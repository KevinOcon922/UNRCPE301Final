PK
     t$v[e�{��~ �~    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2":["pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5":["pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19":["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23":["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28":[],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29":["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"],"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16"],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29":[],"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg":["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg":["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos":["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg":[],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos"],"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos":["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg":["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25"],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-neg":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-pos":[],"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_0":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_1":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_2":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_3":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_4":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_5":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_6":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_7":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8":["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_10":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_11":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_12":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_13":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_14":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_15":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_18":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_19":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_20":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_21":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_22":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_23":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_26":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_27":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_32":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_34":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_35":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_36":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_37":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_40":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_41":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_42":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_43":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_46":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_56":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_57":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_58":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_59":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_60":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_61":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8"],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_68":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_69":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_70":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_71":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_72":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_73":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_74":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_75":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_76":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_77":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_78":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_79":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_80":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_81":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_82":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_83":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84":[],"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_85":[],"pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_0":[],"pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29"],"pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_0":[],"pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19"],"pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_0":[],"pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23"],"pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_0":[],"pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_1":[],"pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_0":[],"pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_1":[],"pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_2":[],"pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_3":[],"pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_0":[],"pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_1":[],"pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_2":[],"pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_3":[],"pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_0":[],"pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_1":[],"pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_0":[],"pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_1":[],"pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_0":[],"pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_1":[],"pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_2":[],"pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_3":[],"pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_0":[],"pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_1":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_0":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_2":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_4":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_6":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_8":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_10":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_12":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_14":[],"pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15":[],"pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2"],"pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5"],"pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_0":[],"pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_1":[],"pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_2":[],"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"],"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"],"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg"],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_0":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_1":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_2":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_3":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_4":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_5":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_6":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_7":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_8":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_9":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_10":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_11":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_12":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_13":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_14":[],"pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_15":[],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6":["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7":["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8":["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9":["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"],"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10":["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"],"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6"],"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7"],"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"],"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9"],"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10"],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg"],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_2":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_3":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_8":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_11":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_12":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_13":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_14":[],"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_15":[],"pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0":[],"pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1":[],"pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2":[],"pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3":[],"pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_4":[],"pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_0":[],"pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_1":[],"pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_0":[],"pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_1":[],"pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_0":[],"pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_1":[],"pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_0":[],"pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_1":[]},"pin_to_color":{"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0":"#bb00ff","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1":"#ff6600","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2":"#ff3232","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2":"#FF0000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3":"#189AB4","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3":"#9caeaa","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5":"#1464c8","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5":"#189AB4","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6":"#90FB92","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7":"#FF0000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8":"#FF0000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9":"#bd684c","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10":"#189AB4","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11":"#999999","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14":"#735348","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19":"#e9e943","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23":"#74b576","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26":"#e94343","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28":"#000000","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29":"#58a5e1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8":"#005F39","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10":"#95003A","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15":"#FF937E","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16":"#001544","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17":"#91D0CB","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18":"#007DB5","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25":"#189AB4","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26":"#FF0000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27":"#e5d545","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28":"#8b7d04","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29":"#000000","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos":"#FF0000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg":"#189AB4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos":"#FF0000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg":"#189AB4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos":"#FF0000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg":"#189AB4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos":"#FF0000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg":"#189AB4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg":"#189AB4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg":"#189AB4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos":"#FF0000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg":"#000000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos":"#FF0000","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos":"#FF0000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg":"#189AB4","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-neg":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-pos":"#000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_0":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_1":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_2":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_3":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_4":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_5":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_6":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_7":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8":"#dddddd","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9":"#bd684c","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_10":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_11":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_12":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_13":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_14":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_15":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16":"#8b7d04","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17":"#e5d545","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_18":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_19":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_20":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_21":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_22":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_23":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_26":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_27":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28":"#5FAD4E","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29":"#ed81ef","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30":"#f90158","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31":"#e2fe0b","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_32":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33":"#bb00ff","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_34":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_35":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_36":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_37":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38":"#FF0000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39":"#189AB4","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_40":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_41":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_42":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_43":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44":"#999999","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45":"#735348","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_46":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47":"#9caeaa","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48":"#90FB92","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49":"#ff6600","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52":"#e9e943","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53":"#74b576","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54":"#e94343","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55":"#58a5e1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_56":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_57":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_58":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_59":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_60":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_61":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62":"#007DB5","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63":"#91D0CB","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64":"#001544","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65":"#FF937E","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66":"#95003A","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67":"#005F39","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_68":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_69":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_70":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_71":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_72":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_73":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_74":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_75":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_76":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_77":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_78":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_79":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_80":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_81":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_82":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_83":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84":"#000000","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_85":"#000000","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_0":"#000000","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1":"#58a5e1","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_0":"#000000","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1":"#e9e943","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_0":"#000000","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1":"#74b576","pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_0":"#000000","pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_1":"#000000","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_0":"#000000","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_1":"#000000","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_2":"#000000","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_3":"#000000","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_0":"#000000","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_1":"#000000","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_2":"#000000","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_3":"#000000","pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_0":"#000000","pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_1":"#000000","pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_0":"#000000","pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_1":"#000000","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_0":"#000000","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_1":"#000000","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_2":"#000000","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_3":"#000000","pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_0":"#000000","pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_1":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_0":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_2":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_4":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_6":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_8":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_10":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_12":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_14":"#000000","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15":"#000000","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0":"#ff3232","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1":"#1464c8","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_0":"#000000","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_1":"#000000","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_2":"#000000","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0":"#dddddd","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1":"#FF0000","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2":"#189AB4","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_0":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_1":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_2":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_3":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_4":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_5":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_6":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_7":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_8":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_9":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_10":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_11":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_12":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_13":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_14":"#000000","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_15":"#000000","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0":"#5FAD4E","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1":"#ed81ef","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2":"#f90158","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3":"#e2fe0b","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4":"#FF0000","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5":"#189AB4","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6":"#1642b2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7":"#ef9cdb","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8":"#eed145","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9":"#f2681c","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10":"#cc1212","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0":"#1642b2","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1":"#ef9cdb","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2":"#eed145","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3":"#f2681c","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4":"#cc1212","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1":"#189AB4","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_2":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_3":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4":"#FF0000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5":"#189AB4","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_8":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_11":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_12":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_13":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_14":"#000000","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_15":"#000000","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0":"#000000","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1":"#000000","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2":"#000000","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3":"#000000","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_4":"#000000","pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_0":"#000000","pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_1":"#000000","pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_0":"#000000","pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_1":"#000000","pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_0":"#000000","pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_1":"#000000","pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_0":"#000000","pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_1":"#000000"},"pin_to_state":{"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29":"neutral","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29":"neutral","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos":"neutral","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-neg":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-pos":"neutral","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_0":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_1":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_2":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_3":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_4":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_5":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_6":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_7":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_10":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_11":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_12":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_13":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_14":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_15":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_18":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_19":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_20":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_21":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_22":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_23":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_26":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_27":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_32":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_34":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_35":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_36":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_37":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_40":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_41":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_42":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_43":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_46":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_56":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_57":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_58":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_59":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_60":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_61":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_68":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_69":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_70":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_71":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_72":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_73":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_74":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_75":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_76":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_77":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_78":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_79":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_80":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_81":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_82":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_83":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84":"neutral","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_85":"neutral","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_0":"neutral","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1":"neutral","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_0":"neutral","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1":"neutral","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_0":"neutral","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1":"neutral","pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_0":"neutral","pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_1":"neutral","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_0":"neutral","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_1":"neutral","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_2":"neutral","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_3":"neutral","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_0":"neutral","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_1":"neutral","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_2":"neutral","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_3":"neutral","pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_0":"neutral","pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_1":"neutral","pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_0":"neutral","pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_1":"neutral","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_0":"neutral","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_1":"neutral","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_2":"neutral","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_3":"neutral","pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_0":"neutral","pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_1":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_0":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_2":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_4":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_6":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_8":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_10":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_12":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_14":"neutral","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15":"neutral","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0":"neutral","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1":"neutral","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_0":"neutral","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_1":"neutral","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_2":"neutral","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0":"neutral","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1":"neutral","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_0":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_1":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_2":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_3":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_4":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_5":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_6":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_7":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_8":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_9":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_10":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_11":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_12":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_13":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_14":"neutral","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_15":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9":"neutral","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10":"neutral","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0":"neutral","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1":"neutral","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2":"neutral","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3":"neutral","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_2":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_3":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_8":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_11":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_12":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_13":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_14":"neutral","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_15":"neutral","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0":"neutral","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1":"neutral","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2":"neutral","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3":"neutral","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_4":"neutral","pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_0":"neutral","pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_1":"neutral","pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_0":"neutral","pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_1":"neutral","pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_0":"neutral","pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_1":"neutral","pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_0":"neutral","pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_1":"neutral"},"next_color_idx":31,"wires_placed_in_order":[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-pos"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_1_polarity-neg"],["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-neg","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-neg"],["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62_polarity-pos","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_62_polarity-pos"],["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62_polarity-neg","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_62_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_4","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_4_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_8","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_8_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_11","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_11_polarity-neg"],["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2"],["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_6"],["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_13"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_6","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_13","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_15","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_19","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_1","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_2","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_5","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_7_polarity-neg"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_27"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_28"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_29"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_30"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_31"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_32"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_33"],["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_34"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_27"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_33","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_33","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_29","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_25","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_25_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_23","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_23_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_24","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"],["pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_31"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_35","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_29","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_41","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_43","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_47_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_42","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_48_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_47","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_43_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_48","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_42_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_49","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_41_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_50","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_51","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_40_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_52","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_57","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_58","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_59","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_60","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_61","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_39_polarity-pos"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_38_polarity-neg"],["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"],["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2_polarity-pos"],["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_3_polarity-neg"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"],["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6"],["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7"],["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7"],["pin-type-fake_2","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-fake_3"],["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_51_polarity-neg","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36"],["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_52_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"],["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1"],["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2"],["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6"],["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11"],["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos"],["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg"],["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos"],["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg"],["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29"],["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23"],["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"],["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50"],["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg"],["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9"],["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"],["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg"],["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1"],["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"],["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"],["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg"],["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"],["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"],["pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24"],["pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1"],["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"],["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-pos"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_1_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-neg","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-neg"]]],[[],[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62_polarity-pos","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_62_polarity-pos"]]],[[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-neg","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-neg"]],[]],[[],[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62_polarity-neg","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_62_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-neg"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-neg"]],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_4","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_4_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_8","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_8_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_11","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_11_polarity-neg"]]],[[],[["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2"]]],[[],[["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_6"]]],[[],[["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_13"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_6","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_13","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_15","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_19","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_1","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-pos"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_1","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-pos"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_2","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-pos"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_5","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_7_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_27"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_28"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_29"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_30"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_31"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_32"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_33"]]],[[],[["pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_34"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_27"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_33","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_33","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_33","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34_polarity-pos"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_29","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_34","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_33","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_32","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_31","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_30","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_29","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_28","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_27","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1"]],[]],[[],[]],[[],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_33","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_29","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34_polarity-pos"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_25","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_25_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_23","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_23_polarity-pos"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_24","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36_polarity-pos"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]]],[[],[["pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_31"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_35","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_29","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_41","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_43","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_47_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_42","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_48_polarity-pos"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_41","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_43","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_47_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_42","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_48_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62_polarity-pos","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_62_polarity-pos"]],[]],[[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62_polarity-neg","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_62_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_47","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_43_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_48","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_42_polarity-pos"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_49","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_41_polarity-pos"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_50","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_51","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_40_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_52","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_57","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_58","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_59","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_60","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_61","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_39_polarity-pos"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_38_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36_polarity-pos"]],[]],[[],[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"]]],[[],[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2_polarity-pos"]]],[[],[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_3_polarity-neg"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4"]]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"]]],[[],[["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6"]]],[[],[["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7"]]],[[],[["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"]],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5"]],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_29","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_30","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_35","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_19","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_15","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_60","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_59","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_58","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_57","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_52","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_50","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_6","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_13","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]],[]],[[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_3_polarity-neg"]],[]],[[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2_polarity-pos"]],[]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_1_polarity-neg"]],[]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-pos"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_24","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_31","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_34","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]],[]],[[],[]],[[],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36"]],[]],[[],[["pin-type-fake_2","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36"]]],[[],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-fake_3"]]],[[],[]],[[],[]],[[],[]],[[["pin-type-fake_2","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36"]],[]],[[],[["pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_51_polarity-neg","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36"]]],[[],[]],[[["pin-type-fake_3","pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32"]],[]],[[],[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_52_polarity-neg"]]],[[],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_36","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_51_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_52_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_62","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_38_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_61","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_39_polarity-pos"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_51","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_40_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_49","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_41_polarity-pos"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_48","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_42_polarity-pos"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_47","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_43_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_2","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_6","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_13","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"]]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_2","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_0_polarity-pos"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_5","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_7_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_0_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_4","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_4_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_8","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_8_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_11","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_11_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_23","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_23_polarity-pos"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_25","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_1_25_polarity-neg"]],[]],[[["pin-type-breadboard_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32","pin-type-power-rail_5689fad3-77a5-4981-a424-b3d9978fd7e9_0_32_polarity-neg"]],[]],[[],[["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1"]],[]],[[],[["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2"]]],[[],[["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6"]]],[[],[["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1"]],[]],[[],[["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg"]],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos"]]],[[],[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos"]],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg"]]],[[],[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg"]],[]],[[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg"]],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg"]]],[[],[]],[[],[]],[[],[["pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29"]]],[[],[["pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23"]]],[[],[["pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"]],[]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"]],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg"]],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]]],[[],[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"]],[]],[[],[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos"]]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos"]],[]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg"]]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"]]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"]],[]],[[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"]],[]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]],[]],[[],[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos"]],[]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg"]],[]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"]]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos"]]],[[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"]]],[[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos"]],[]],[[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg"]],[]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9"]]],[[],[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"]]],[[],[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg"]]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"]],[]],[[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"]],[]],[[],[["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"]]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]],[]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1"]]],[[],[["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9"]],[]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"]]],[[],[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"]]],[[["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2"]],[]],[[],[["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"]],[]],[[],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg"]]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg"]]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]],[]],[[],[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"]]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos"]],[]],[[["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"]]],[[],[["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"]]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg"]],[]],[[["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"]]],[[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"]],[]],[[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"]],[]],[[],[["pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24"]]],[[],[["pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1"]]],[[],[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0"]]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3"]],[]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2"]],[]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1"]],[]],[[["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"]]],[[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"]],[]],[[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg"]],[]],[[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos"]],[]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"]]],[[],[["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0":"0000000000000028","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1":"0000000000000026","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2":"0000000000000023","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2":"0000000000000017","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3":"0000000000000008","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3":"0000000000000055","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5":"0000000000000022","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5":"0000000000000001","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6":"0000000000000027","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7":"0000000000000007","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8":"0000000000000002","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9":"0000000000000041","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10":"0000000000000003","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11":"0000000000000010","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14":"0000000000000009","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19":"0000000000000006","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23":"0000000000000005","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26":"0000000000000011","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28":"_","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29":"0000000000000004","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5":"0000000000000029","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5":"0000000000000029","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6":"0000000000000030","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6":"0000000000000030","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7":"0000000000000031","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7":"0000000000000031","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8":"0000000000000035","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9":"0000000000000032","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9":"0000000000000032","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10":"0000000000000036","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15":"0000000000000037","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16":"0000000000000038","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17":"0000000000000039","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18":"0000000000000040","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19":"0000000000000034","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19":"0000000000000034","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20":"0000000000000033","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20":"0000000000000033","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25":"0000000000000013","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26":"0000000000000014","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27":"0000000000000016","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28":"0000000000000053","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29":"_","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos":"0000000000000047","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg":"0000000000000046","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_0_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos":"0000000000000017","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg":"0000000000000008","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_4_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_4_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_6_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos":"0000000000000007","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg":"0000000000000001","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_8_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos":"0000000000000002","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_9_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_10_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg":"0000000000000003","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_11_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_12_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_12_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_13_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_13_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_14_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_15_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_15_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_16_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_16_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_17_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_17_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_18_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_18_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_19_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_20_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_20_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_21_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_21_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_22_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_22_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_23_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_24_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_24_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_25_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_25_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_26_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg":"0000000000000012","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_27_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_28_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-pos":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg":"0000000000000054","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos":"0000000000000015","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-neg":"_","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos":"0000000000000018","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg":"0000000000000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos":"0000000000000042","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg":"0000000000000021","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_0_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos":"0000000000000019","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg":"0000000000000043","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_1_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_2_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_2_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_3_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_3_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_4_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_4_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg":"0000000000000029","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos":"0000000000000030","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos":"0000000000000031","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_8_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg":"0000000000000032","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_10_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_11_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_11_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_12_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_12_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_13_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_13_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_14_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_14_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_15_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_16_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_17_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos":"0000000000000018","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos":"0000000000000034","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg":"0000000000000000","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg":"0000000000000033","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_21_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_21_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_22_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos":"0000000000000014","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_23_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg":"0000000000000013","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_24_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_24_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_25_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_26_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_27_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_28_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_29_polarity-neg":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-pos":"_","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_29_polarity-neg":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_0":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_1":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_2":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_3":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_4":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_5":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_6":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_7":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8":"0000000000000020","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9":"0000000000000041","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_10":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_11":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_12":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_13":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_14":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_15":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16":"0000000000000053","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17":"0000000000000016","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_18":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_19":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_20":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_21":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_22":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_23":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_24":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_25":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_26":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_27":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28":"0000000000000045","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29":"0000000000000044","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30":"0000000000000025","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31":"0000000000000024","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_32":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33":"0000000000000028","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_34":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_35":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_36":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_37":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38":"0000000000000042","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39":"0000000000000021","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_40":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_41":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_42":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_43":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44":"0000000000000010","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45":"0000000000000009","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_46":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47":"0000000000000055","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48":"0000000000000027","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49":"0000000000000026","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_50":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_51":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52":"0000000000000006","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53":"0000000000000005","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54":"0000000000000011","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55":"0000000000000004","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_56":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_57":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_58":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_59":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_60":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_61":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62":"0000000000000040","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63":"0000000000000039","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64":"0000000000000038","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65":"0000000000000037","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66":"0000000000000036","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67":"0000000000000035","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_68":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_69":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_70":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_71":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_72":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_73":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_74":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_75":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_76":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_77":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_78":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_79":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_80":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_81":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_82":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_83":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_84":"_","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_85":"_","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_0":"_","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1":"0000000000000004","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_0":"_","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1":"0000000000000006","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_0":"_","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1":"0000000000000005","pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_0":"_","pin-type-component_9599c2c6-ff11-4398-b0b0-57d2801063a2_1":"_","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_0":"_","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_1":"_","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_2":"_","pin-type-component_0bb3fad2-c6fc-4e08-b85d-d0ae222291a4_3":"_","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_0":"_","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_1":"_","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_2":"_","pin-type-component_a35b23da-4320-4bb1-9803-5623435010b8_3":"_","pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_0":"_","pin-type-component_35403b54-b36e-41ad-adc9-689326b1737d_1":"_","pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_0":"_","pin-type-component_d8350423-52d2-45ba-9cfc-9ffab1e52410_1":"_","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_0":"_","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_1":"_","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_2":"_","pin-type-component_f4b5bb34-dfd2-4497-8b35-3c669d760eef_3":"_","pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_0":"_","pin-type-component_0f89696f-8c6b-487e-8d1f-581cd6a2b8bb_1":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_0":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_1":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_2":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_3":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_4":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_5":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_6":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_7":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_8":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_9":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_10":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_11":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_12":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_13":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_14":"_","pin-type-component_46ad218f-026e-4be7-9a05-692d65968ceb_15":"_","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0":"0000000000000023","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1":"0000000000000022","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_0":"_","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_1":"_","pin-type-component_25f1d489-7130-4e16-bf56-2cf3a4b82b0f_2":"_","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0":"0000000000000020","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1":"0000000000000019","pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2":"0000000000000043","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_0":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_1":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_2":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_3":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_4":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_5":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_6":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_7":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_8":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_9":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_10":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_11":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_12":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_13":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_14":"_","pin-type-component_03536000-14c0-4aaf-abcc-70e8ef6b2088_15":"_","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0":"0000000000000045","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1":"0000000000000044","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2":"0000000000000025","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3":"0000000000000024","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4":"0000000000000047","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5":"0000000000000046","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6":"0000000000000048","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7":"0000000000000049","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8":"0000000000000050","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9":"0000000000000051","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10":"0000000000000052","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0":"0000000000000048","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1":"0000000000000049","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2":"0000000000000050","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3":"0000000000000051","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4":"0000000000000052","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_0":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1":"0000000000000054","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_2":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_3":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4":"0000000000000015","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5":"0000000000000012","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_6":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_7":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_8":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_9":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_10":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_11":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_12":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_13":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_14":"_","pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_15":"_","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_0":"_","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_1":"_","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_2":"_","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_3":"_","pin-type-component_ed7be971-3bf8-4999-a879-84514691bc16_4":"_","pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_0":"_","pin-type-component_477ab0cf-d7c8-4735-9d85-297b1c25bcdd_1":"_","pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_0":"_","pin-type-component_56960671-d035-4d6b-9122-a3075a17d45a_1":"_","pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_0":"_","pin-type-component_5a09c35a-bb24-444f-b5a5-73cfd27e91a0_1":"_","pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_0":"_","pin-type-component_3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7_1":"_"},"component_id_to_pins":{"e089bc97-3efd-4a29-a939-30b226883bf4":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","42","43","44","45","46","47","48","49","50","51","52","53","54","55","56","57","58","59","60","61","62","63","64","65","66","67","68","69","70","71","72","73","74","75","76","77","78","79","80","81","82","83","84","85"],"a8f06db4-bc8a-4ced-9f16-e6b21dbe1539":["0","1"],"a4427fbb-4a98-452f-b0a1-621dd7a1661f":["0","1"],"5b6e25a5-f561-4e8d-a22d-e361c10aa6f3":["0","1"],"9599c2c6-ff11-4398-b0b0-57d2801063a2":["0","1"],"0bb3fad2-c6fc-4e08-b85d-d0ae222291a4":["0","1","2","3"],"a35b23da-4320-4bb1-9803-5623435010b8":["0","1","2","3"],"35403b54-b36e-41ad-adc9-689326b1737d":["0","1"],"d8350423-52d2-45ba-9cfc-9ffab1e52410":["0","1"],"f4b5bb34-dfd2-4497-8b35-3c669d760eef":["0","1","2","3"],"0f89696f-8c6b-487e-8d1f-581cd6a2b8bb":["0","1"],"46ad218f-026e-4be7-9a05-692d65968ceb":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"047cb0d4-3606-44fe-91b7-6e30f1913e78":["0","1"],"25f1d489-7130-4e16-bf56-2cf3a4b82b0f":["0","1","2"],"f9130057-4ade-4f7f-a4ec-80702a655d28":["0","1","2"],"03536000-14c0-4aaf-abcc-70e8ef6b2088":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"54195fcb-e342-4208-b4ce-f4de03f5d795":["0","1","2","3","4","5","6","7","8","9","10"],"b466983e-1896-401c-90c5-57535cb2e5a6":["0","1","2","3","4"],"1c5b82ec-d40c-4873-a511-0cb71ebcb6c9":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"cf24b1b8-b621-4d44-91d7-a5bfcba42892":[],"a29b71f0-9777-419b-92b7-b0c33062b8d8":[],"aa98d916-656a-4f5c-9420-ef145600d396":[],"6ff94e4c-22b2-46b8-9016-5ceb2c80493e":[],"958e2f7d-be7f-4a65-aac7-b7f6a8f0ab67":[],"d8ce3ba2-5633-461e-bd3b-48cbf14f7e4c":[],"465db3f5-2c24-48c7-9f83-db45be687fdb":[],"7ed77f21-a242-4d15-8707-6b1df9e1155e":[],"e42acb99-bbba-4da4-8d6d-7c9b539be5b4":[],"f2d2aeb9-c40a-44f4-af90-aa33bfe3bc13":[],"adffc0fb-edf6-4614-8d9e-668af8e616c8":[],"ed7be971-3bf8-4999-a879-84514691bc16":["0","1","2","3","4"],"477ab0cf-d7c8-4735-9d85-297b1c25bcdd":["0","1"],"56960671-d035-4d6b-9122-a3075a17d45a":["0","1"],"5a09c35a-bb24-444f-b5a5-73cfd27e91a0":["0","1"],"3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7":["0","1"],"187edb3a-243a-4ca3-8428-c5a109bbe2d4":[]},"uid_to_net":{"_":[],"0000000000000020":["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8"],"0000000000000001":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg"],"0000000000000002":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos"],"0000000000000003":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg"],"0000000000000004":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29","pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55"],"0000000000000005":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23","pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53"],"0000000000000006":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19","pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52"],"0000000000000007":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos"],"0000000000000008":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg"],"0000000000000017":["pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2"],"0000000000000021":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg"],"0000000000000027":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48"],"0000000000000022":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1"],"0000000000000023":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2","pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0"],"0000000000000026":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49"],"0000000000000028":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33"],"0000000000000009":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45"],"0000000000000010":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44"],"0000000000000029":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg"],"0000000000000030":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos"],"0000000000000031":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos"],"0000000000000032":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg"],"0000000000000033":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg"],"0000000000000034":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19","pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos"],"0000000000000035":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67"],"0000000000000036":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66"],"0000000000000037":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65"],"0000000000000038":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64"],"0000000000000039":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63"],"0000000000000040":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62"],"0000000000000043":["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg"],"0000000000000019":["pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos"],"0000000000000042":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos"],"0000000000000015":["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos"],"0000000000000024":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31"],"0000000000000025":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30"],"0000000000000044":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29"],"0000000000000045":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28"],"0000000000000046":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg"],"0000000000000047":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos"],"0000000000000048":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0"],"0000000000000049":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1"],"0000000000000051":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3"],"0000000000000052":["pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10","pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4"],"0000000000000050":["pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2","pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8"],"0000000000000041":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9"],"0000000000000011":["pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54"],"0000000000000054":["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg"],"0000000000000055":["pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47","pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3"],"0000000000000000":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg"],"0000000000000018":["pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos"],"0000000000000012":["pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5","pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg"],"0000000000000013":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg"],"0000000000000014":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26","pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos"],"0000000000000016":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17"],"0000000000000053":["pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28","pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16"]},"uid_to_text_label":{"0000000000000020":"Net 20","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000017":"Net 17","0000000000000021":"Net 21","0000000000000027":"Net 27","0000000000000022":"Net 22","0000000000000023":"Net 23","0000000000000026":"Net 26","0000000000000028":"Net 28","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000029":"Net 29","0000000000000030":"Net 30","0000000000000031":"Net 31","0000000000000032":"Net 32","0000000000000033":"Net 33","0000000000000034":"Net 34","0000000000000035":"Net 35","0000000000000036":"Net 36","0000000000000037":"Net 37","0000000000000038":"Net 38","0000000000000039":"Net 39","0000000000000040":"Net 40","0000000000000043":"Net 43","0000000000000019":"Net 19","0000000000000042":"Net 42","0000000000000015":"Net 15","0000000000000024":"Net 24","0000000000000025":"Net 25","0000000000000044":"Net 44","0000000000000045":"Net 45","0000000000000046":"Net 46","0000000000000047":"Net 47","0000000000000048":"Net 48","0000000000000049":"Net 49","0000000000000051":"Net 51","0000000000000052":"Net 52","0000000000000050":"Net 50","0000000000000041":"Net 41","0000000000000011":"Net 11","0000000000000054":"Net 54","0000000000000055":"Net 55","0000000000000000":"Net 0","0000000000000018":"Net 18","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000016":"Net 16","0000000000000053":"Net 53"},"all_breadboard_info_list":["5689fad3-77a5-4981-a424-b3d9978fd7e9_63_2_True_1127_-447.0000000000006_left","baacc681-4994-4064-8b3a-269f4fbd62a9_30_2_True_879.5000000000001_-229.49999999999997_left","d3e67062-b31b-41bc-8e97-0bb2a0d8f023_30_2_True_1269.5_145.50000000000003_left"],"breadboard_info_list":["baacc681-4994-4064-8b3a-269f4fbd62a9_30_2_True_879.5000000000001_-229.49999999999997_left","d3e67062-b31b-41bc-8e97-0bb2a0d8f023_30_2_True_1269.5_145.50000000000003_left"],"componentsData":[{"compProperties":{},"position":[718.7803885000003,372.5000179999996],"typeId":"972688b5-e2a3-1d53-e820-bc24d2f5082a","componentVersion":15,"instanceId":"e089bc97-3efd-4a29-a939-30b226883bf4","orientation":"up","circleData":[[872.5,515],[887.4999819999998,515],[902.4978804999998,515],[917.5020294999999,515],[932.5020115,515],[947.4999114999998,515],[962.4998934999999,515],[977.4977919999999,515],[737.5001575000005,515],[752.4980575000004,515],[767.5022065000003,515],[782.5021885000003,515],[797.5000870000001,515],[812.5000705000002,515],[827.4979690000002,515],[842.5021180000001,515],[947.4999114999998,229.99999999999977],[932.5020115,229.99999999999977],[917.5020294999999,229.99999999999977],[902.4978804999998,229.99999999999977],[887.4999819999998,229.99999999999977],[872.5,229.99999999999977],[857.5021000000002,229.99999999999977],[842.5021180000001,229.99999999999977],[548.4982975000004,229.99999999999977],[563.5003630000004,229.99999999999977],[578.5003450000004,229.99999999999977],[593.5003270000004,229.99999999999977],[608.5003105000004,229.99999999999977],[623.5002925000005,229.99999999999977],[638.5002745000004,229.99999999999977],[653.5002565000004,229.99999999999977],[668.5002400000004,229.99999999999977],[683.5002220000005,229.99999999999977],[602.5003165000004,515],[617.5003000000004,515],[632.5023655000005,515],[647.5002640000004,515],[662.5002460000004,515],[677.5002280000004,515],[692.5002115000003,515],[707.5022770000004,515],[812.5000705000002,229.99999999999977],[797.5000870000001,229.99999999999977],[782.5021885000003,229.99999999999977],[767.5022065000003,229.99999999999977],[752.4980575000004,229.99999999999977],[737.5001575000005,229.99999999999977],[722.5001755000004,229.99999999999977],[707.5022770000004,229.99999999999977],[992.5019409999998,229.99999999999977],[1007.5019245,229.99999999999977],[992.5019409999998,244.99999999999977],[1007.5019245,244.99999999999977],[992.5019409999998,259.9999999999998],[1007.5019245,259.9999999999998],[992.5019409999998,274.9999999999998],[1007.5019245,274.9999999999998],[992.5019409999998,289.9999999999998],[1007.5019245,289.9999999999998],[992.5019409999998,304.9999999999998],[1007.5019245,304.9999999999998],[992.5019409999998,319.9999999999998],[1007.5019245,319.9999999999998],[992.5019409999998,334.9999999999998],[1007.5019245,334.9999999999998],[992.5019409999998,349.9999999999998],[1007.5019245,349.9999999999998],[992.5019409999998,364.9999999999998],[1007.5019245,364.9999999999998],[992.5019409999998,379.99999999999983],[1007.5019245,379.99999999999983],[992.5019409999998,394.99999999999983],[1007.5019245,394.99999999999983],[992.5019409999998,409.99999999999983],[1007.5019245,409.99999999999983],[992.5019409999998,424.99999999999983],[1007.5019245,424.99999999999983],[992.5019409999998,439.99999999999983],[1007.5019245,439.99999999999983],[992.5019409999998,454.99999999999983],[1007.5019245,454.99999999999983],[992.5019409999998,469.99999999999983],[1007.5019245,469.99999999999983],[992.5019409999998,484.99999999999983],[1007.5019245,484.99999999999983]],"code":"512,folder,{\"name\":\"sketch\",\"id\":\"8da69639-5087-4181-b1f0-3488098e23de\",\"explorerHtmlId\":\"b3a92ac7-826f-4994-b25c-b42d39484557\",\"nameHtmlId\":\"8b794d20-4c52-45c3-9f37-6a22aac27f55\",\"nameInputHtmlId\":\"9550f4a1-68f4-4ed9-a134-ca05b4b8faf9\",\"explorerChildHtmlId\":\"eca1c1cf-43f2-4319-a243-21b7b57d9779\",\"explorerCarrotOpenHtmlId\":\"461264a7-7407-4d1d-a6f7-935240040acb\",\"explorerCarrotClosedHtmlId\":\"c592a505-6ddc-434d-aa6b-8e1796d56299\",\"arduinoBoardFqbn\":\"arduino:avr:mega\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"c2d8af3e-8b3b-4811-9f34-f07b1f0ff89e\",\"explorerHtmlId\":\"c98f0a15-2576-4cbb-a5e0-3eff17e142c7\",\"nameHtmlId\":\"a2e90789-2d60-4844-83ca-24ce9c86fa45\",\"nameInputHtmlId\":\"3a693928-cb0f-4856-a531-1df5db87ed36\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"5aff0c0c-2775-4600-9134-54add2e1cee8\",\"explorerHtmlId\":\"954a1429-055a-4071-bded-f45996928055\",\"nameHtmlId\":\"5b3a3f40-9662-40d1-8521-20614dcb481f\",\"nameInputHtmlId\":\"d20aae69-4572-457d-b32e-1a272264e9d9\",\"code\":\"\"},0,","codeLabelPosition":[718.7803885000004,215.01411799999966],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[174.58349499999647,577.2166699999998],"typeId":"97784b10-4dcd-a3be-9167-75f1272c8490","componentVersion":1,"instanceId":"f9130057-4ade-4f7f-a4ec-80702a655d28","orientation":"right","circleData":[[347.5,560],[347.5,575],[347.5,590]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1258.0816210000003,-2.11849149999901],"typeId":"307d45d2-aa1f-05de-326e-55c453eb206e","componentVersion":4,"instanceId":"1c5b82ec-d40c-4873-a511-0cb71ebcb6c9","orientation":"up","circleData":[[1187.5,-145.00000000000006],[1187.5,-130.0000000000001],[1247.5,-145.00000000000006],[1247.5,-130.00000000000034],[1187.6500000000005,123.80000000000177],[1187.6500000000005,139.1000000000011],[1247.3805730000004,123.81528650000178],[1247.3652865000004,138.98057300000102],[1203.1000000000004,-55.29999999999973],[1218.1000000000004,-55.29999999999973],[1233.1000000000004,-55.29999999999973],[1248.1000000000004,-55.29999999999973],[1203.1000000000004,-40.2999999999996],[1218.1000000000004,-40.2999999999996],[1233.1000000000004,-40.2999999999996],[1248.1000000000004,-40.2999999999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[508.7155825000001,88.8005584999998],"typeId":"ecbd5bee-2226-4f1c-8fdb-aaff666e8628","componentVersion":1,"instanceId":"54195fcb-e342-4208-b4ce-f4de03f5d795","orientation":"right","circleData":[[557.5,140],[557.5,125.50958600000004],[558.949036,112.46820799999992],[558.949036,99.42688850000005],[529.1097235,34.42580600000022],[543.505591,33.526101500000124],[480.52372000000014,151.39208599999984],[481.4234845000001,138.79574749999995],[481.4234845000001,127.09911349999999],[481.4234845000001,115.40247949999994],[482.32318900000007,101.90637800000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[418.9273495000007,-104.31239349999959],"typeId":"7115dd0c-9076-1603-96e1-f4f66aa483df","componentVersion":7,"instanceId":"047cb0d4-3606-44fe-91b7-6e30f1913e78","orientation":"down","circleData":[[602.5,-55.00000000000003],[602.5,-153.8379999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"181","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1361.4770754999997,546.5344084999999],"typeId":"23598c1c-7607-4538-b177-9ab948fb1937","componentVersion":3,"instanceId":"03536000-14c0-4aaf-abcc-70e8ef6b2088","orientation":"up","circleData":[[1172.5,455],[1187.5020834999998,455],[1202.4999999999998,455],[1217.4999999999998,455],[1232.5020834999998,455],[1247.4999999999998,455],[1262.5020834999998,455],[1277.4999999999998,455],[1292.4999999999998,455],[1307.4999999999998,455],[1322.4999999999998,455],[1337.5020834999998,455],[1352.4999999999998,455],[1367.4999999999986,455],[1382.5020834999991,455],[1397.4999999999968,455]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"28BYJ-48 Stepper Motor","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#ffffff","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[289.6900363232473,64.69742282664527],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"cf24b1b8-b621-4d44-91d7-a5bfcba42892","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"DC Gear Motor (3-6V)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[536.4393288796678,-187.43397919321],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"a29b71f0-9777-419b-92b7-b0c33062b8d8","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"DHT11","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[831.273340801352,-186.299531050575],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"aa98d916-656a-4f5c-9420-ef145600d396","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Water Level Sensor","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[181.05295828959504,494.6940297400324],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"6ff94e4c-22b2-46b8-9016-5ceb2c80493e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Arduino Mega 2560","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[351.7895325351838,374.3098845483647],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"958e2f7d-be7f-4a65-aac7-b7f6a8f0ab67","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LCD Display","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1067.7203638622111,617.000898110022],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"d8ce3ba2-5633-461e-bd3b-48cbf14f7e4c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Power Supply Module","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1270.0456979671255,-189.1692806246767],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"465db3f5-2c24-48c7-9f83-db45be687fdb","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Potentiometer","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[838.5892144950641,-43.270675242585234],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"7ed77f21-a242-4d15-8707-6b1df9e1155e","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Push Buttons","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[909.5264903944395,41.28726466905661],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"e42acb99-bbba-4da4-8d6d-7c9b539be5b4","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LEDs","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1067.7282863150049,-60.362173735363854],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"f2d2aeb9-c40a-44f4-af90-aa33bfe3bc13","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"28BYJ-48 Motor Driver","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#ffffff","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[509.8240899189391,-5.546514544180802],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"adffc0fb-edf6-4614-8d9e-668af8e616c8","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[159.063541,124.99791650000023],"typeId":"de09217e-3b73-b82d-0145-70b2df9a4b72","componentVersion":1,"instanceId":"b466983e-1896-401c-90c5-57535cb2e5a6","orientation":"left","circleData":[[407.5,155],[407.5,140.00208350000014],[407.5,124.99791650000009],[407.5,110.00104099999992],[407.5,95.00104100000016]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"initTime":{"version":2,"id":"initTime","label":"Initial Time","description":"Initial time of the RTC: \"0\", \"now\", or a valid ISO 8601 date string","units":"","type":"string","value":"now","displayFormat":"input","showOnComp":false}},"position":[1513.896763,229.63745299999977],"typeId":"9f0127e3-b141-4b6c-b341-c271412e4837","componentVersion":2,"instanceId":"ed7be971-3bf8-4999-a879-84514691bc16","orientation":"left","circleData":[[1472.5,290],[1487.5,290],[1502.5,290],[1517.5,290],[1532.4999999999998,290]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1137.5000244999992,7.500006500000104],"typeId":"117aab52-1b06-40f5-98b6-df63a601b0e6","componentVersion":3,"instanceId":"a8f06db4-bc8a-4ced-9f16-e6b21dbe1539","orientation":"up","circleData":[[1127.499999999999,50.00000000000012],[1150.761384999999,49.87209200000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1090.0478664999987,22.2029990000001],"typeId":"5f0a7f7f-5908-4e39-94d8-2714a0462581","componentVersion":2,"instanceId":"9599c2c6-ff11-4398-b0b0-57d2801063a2","orientation":"up","circleData":[[1082.4999999999986,50.00000000000012],[1097.4999999999986,50.00000000000012]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[742.1402533379207,-45.68155936351795],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"0f89696f-8c6b-487e-8d1f-581cd6a2b8bb","orientation":"up","circleData":[[737.5000000000001,-54.9999999999996],[752.5000000000001,-54.9999999999996]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[759.9999984999996,-144.99991599999956],"typeId":"a76bb123-3d3c-417d-b1f3-c8417efb7bc7","componentVersion":1,"instanceId":"f4b5bb34-dfd2-4497-8b35-3c669d760eef","orientation":"up","circleData":[[737.4999999999997,-84.9999999999998],[752.4999999999997,-84.9999999999998],[767.4999999999995,-84.9999999999998],[782.4999999999995,-84.9999999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1047.5000244999983,7.500024500000144],"typeId":"a70bb5a8-99ed-4f1b-882e-eac0873b75ef","componentVersion":5,"instanceId":"5b6e25a5-f561-4e8d-a22d-e361c10aa6f3","orientation":"up","circleData":[[1037.4999999999982,50.00000000000012],[1060.7613849999984,49.872090500000134]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"PTS645SL50-2 LFS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"C&K Components","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[932.2705000000001,-2.498499999999126],"typeId":"232ac546-6e45-4194-9a27-0fa614949a21","componentVersion":3,"instanceId":"a35b23da-4320-4bb1-9803-5623435010b8","orientation":"down","circleData":[[917.5000000000001,20.0000000000005],[917.5000000000001,-24.99999999999941],[947.4999999999995,20.0000000000005],[947.5000000000002,-24.99999999999941]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"","type":"string","value":"10000","displayFormat":"dropdown","options":[{"label":"100","value":"100"},{"label":"1000","value":"1000"},{"label":"10000","value":"10000"},{"label":"100000","value":"100000"},{"label":"1000000","value":"1000000"}],"showOnComp":false,"isVisibleToUser":true,"name":"Resistance","required":true}},"position":[842.5,-3.2499999999997726],"typeId":"cc03c8ee-909a-4085-863c-ededb100351c","componentVersion":3,"instanceId":"25f1d489-7130-4e16-bf56-2cf3a4b82b0f","orientation":"down","circleData":[[857.5,-24.999999999999694],[842.5000000000002,18.500000000000213],[827.5000000000002,-24.999999999999694]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"PTS645SL50-2 LFS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"C&K Components","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[887.2705000000005,-2.498499999999126],"typeId":"232ac546-6e45-4194-9a27-0fa614949a21","componentVersion":3,"instanceId":"0bb3fad2-c6fc-4e08-b85d-d0ae222291a4","orientation":"down","circleData":[[872.4999999999999,20.000000000000497],[872.5,-24.999999999999467],[902.5,20.000000000000497],[902.5,-24.999999999999467]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[987.5000245000003,7.499988500000207],"typeId":"1310de1e-180e-4aed-a1c6-f80032a2bfde","componentVersion":4,"instanceId":"a4427fbb-4a98-452f-b0a1-621dd7a1661f","orientation":"up","circleData":[[977.5000000000001,50.00000000000012],[1000.7613850000009,49.87209200000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4700","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[902.5000000000002,-92.5],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"35403b54-b36e-41ad-adc9-689326b1737d","orientation":"left","circleData":[[902.5000000000002,-54.9999999999996],[902.5000000000002,-130.00000000000014]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[760.0000000000001,-1.4950014999993968],"typeId":"155f7657-2d2d-eaf2-280f-5c76a41d0679","componentVersion":1,"instanceId":"46ad218f-026e-4be7-9a05-692d65968ceb","orientation":"up","circleData":[[707.5000000000001,20.0000000000005],[707.5000000000001,-22.99000299999944],[812.5000015000003,20.0000000000005],[812.5000015000003,-22.99000299999944],[722.5000000000001,20.0000000000005],[722.5000000000001,-22.99000299999944],[737.5000000000001,20.0000000000005],[737.5000000000001,-22.99000299999944],[752.5000000000001,20.0000000000005],[752.5000000000001,-22.99000299999944],[767.5000015000002,20.0000000000005],[767.5000015000002,-22.99000299999944],[782.5000015000002,20.0000000000005],[782.5000015000002,-22.99000299999944],[797.5000015000003,20.0000000000005],[797.5000015000003,-22.99000299999944]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4700","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[947.4999999999995,-92.5],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"d8350423-52d2-45ba-9cfc-9ffab1e52410","orientation":"left","circleData":[[947.5000000000001,-54.9999999999996],[947.5000000000001,-129.9999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[977.5,102.5],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"477ab0cf-d7c8-4735-9d85-297b1c25bcdd","orientation":"left","circleData":[[977.5000000000001,125],[977.5000000000001,80]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[1037.5,102.50000000000003],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"56960671-d035-4d6b-9122-a3075a17d45a","orientation":"left","circleData":[[1037.5,125],[1037.5,79.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[1082.5,102.49999999999997],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"5a09c35a-bb24-444f-b5a5-73cfd27e91a0","orientation":"left","circleData":[[1082.5,125],[1082.5,79.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[1127.5,102.5],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"3a30102b-0e2b-4ec7-854f-76a7ba9ccbb7","orientation":"left","circleData":[[1127.5,125],[1127.5,80.00000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"RTC DS1307","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"12","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1514.426481794541,133.33159025673595],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":3,"instanceId":"187edb3a-243a-4ca3-8428-c5a109bbe2d4","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-219.99992","left":"-108.74896","width":"1707.04686","height":"873.43325","x":"-108.74896","y":"-219.99992"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#dddddd\",\"startPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8\",\"endPinId\":\"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0\",\"rawStartPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_8\",\"rawEndPinId\":\"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"737.5001575000_515.0000000000\\\",\\\"737.5001575000_560.0000000000\\\",\\\"347.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_1_5_3\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_7_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_-70.0000000000\\\",\\\"812.5000000000_-70.0000000000\\\",\\\"812.5000000000_-145.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_3\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_8_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_-70.0000000000\\\",\\\"827.5000000000_-130.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_3\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_10_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_-70.0000000000\\\",\\\"857.5000000000_-145.0000000000\\\"]}\"}","{\"color\":\"#58a5e1\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29\",\"endPinId\":\"pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_2\",\"rawEndPinId\":\"pin-type-component_a8f06db4-bc8a-4ced-9f16-e6b21dbe1539_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_50.0000000000\\\",\\\"1150.7613850000_50.0000000000\\\",\\\"1150.7613850000_49.8720920000\\\"]}\"}","{\"color\":\"#58a5e1\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_0\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_55\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_80.0000000000\\\",\\\"1142.5000000000_95.0000000000\\\",\\\"1037.5000000000_95.0000000000\\\",\\\"1037.5000000000_260.0000000000\\\",\\\"1007.5019245000_260.0000000000\\\"]}\"}","{\"color\":\"#74b576\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23\",\"endPinId\":\"pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_2\",\"rawEndPinId\":\"pin-type-component_5b6e25a5-f561-4e8d-a22d-e361c10aa6f3_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_50.0000000000\\\",\\\"1060.7613850000_50.0000000000\\\",\\\"1060.7613850000_49.8720905000\\\"]}\"}","{\"color\":\"#74b576\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_23_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_53\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_65.0000000000\\\",\\\"1007.5000000000_65.0000000000\\\",\\\"1007.5000000000_200.0000000000\\\",\\\"1007.5019245000_200.0000000000\\\",\\\"1007.5019245000_245.0000000000\\\"]}\"}","{\"color\":\"#e9e943\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19\",\"endPinId\":\"pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_2\",\"rawEndPinId\":\"pin-type-component_a4427fbb-4a98-452f-b0a1-621dd7a1661f_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_50.0000000000\\\",\\\"1000.7613850000_50.0000000000\\\",\\\"1000.7613850000_49.8720920000\\\"]}\"}","{\"color\":\"#e9e943\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_19_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_52\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_65.0000000000\\\",\\\"992.5000000000_200.0000000000\\\",\\\"992.5019410000_200.0000000000\\\",\\\"992.5019410000_245.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_0\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_7_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_80.0000000000\\\",\\\"812.5000000000_140.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_0\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_3_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"752.5000000000_80.0000000000\\\",\\\"752.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_1_2_3\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_1_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"737.5000000000_-70.0000000000\\\",\\\"722.5000000000_-70.0000000000\\\",\\\"722.5000000000_-130.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg\",\"rawStartPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_39\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5002280000_515.0000000000\\\",\\\"677.5002280000_537.5000000000\\\",\\\"1090.0000000000_537.5000000000\\\",\\\"1090.0000000000_500.0000000000\\\",\\\"1097.5000000000_500.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_6_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_48\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_65.0000000000\\\",\\\"797.5000000000_185.0000000000\\\",\\\"722.5001755000_185.0000000000\\\",\\\"722.5001755000_230.0000000000\\\"]}\"}","{\"color\":\"#1464c8\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5\",\"endPinId\":\"pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_5_3\",\"rawEndPinId\":\"pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_35.0000000000\\\",\\\"647.5000000000_35.0000000000\\\",\\\"647.5000000000_-153.8380000000\\\",\\\"602.5000000000_-153.8380000000\\\"]}\"}","{\"color\":\"#ff3232\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2\",\"endPinId\":\"pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_2_2\",\"rawEndPinId\":\"pin-type-component_047cb0d4-3606-44fe-91b7-6e30f1913e78_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"737.5000000000_50.0000000000\\\",\\\"632.5000000000_50.0000000000\\\",\\\"632.5000000000_-55.0000000000\\\",\\\"602.5000000000_-55.0000000000\\\"]}\"}","{\"color\":\"#ff6600\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_1_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_49\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.5000000000_65.0000000000\\\",\\\"730.0000000000_65.0000000000\\\",\\\"730.0000000000_177.5000000000\\\",\\\"707.5022770000_177.5000000000\\\",\\\"707.5022770000_230.0000000000\\\"]}\"}","{\"color\":\"#bb00ff\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_0\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_33\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.5000000000_80.0000000000\\\",\\\"715.0000000000_80.0000000000\\\",\\\"715.0000000000_170.0000000000\\\",\\\"683.5002220000_170.0000000000\\\",\\\"683.5002220000_230.0000000000\\\"]}\"}","{\"color\":\"#735348\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_14_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_45\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"917.5000000000_65.0000000000\\\",\\\"857.5000000000_65.0000000000\\\",\\\"857.5000000000_200.0000000000\\\",\\\"767.5022065000_200.0000000000\\\",\\\"767.5022065000_230.0000000000\\\"]}\"}","{\"color\":\"#999999\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_11_0\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_44\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_80.0000000000\\\",\\\"872.5000000000_207.5000000000\\\",\\\"782.5021885000_207.5000000000\\\",\\\"782.5021885000_230.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5\",\"endPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_5_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1172.5000000000_395.0000000000\\\",\\\"1172.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_5_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1172.5000000000_305.0000000000\\\",\\\"1172.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6\",\"endPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_6_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.5000000000_395.0000000000\\\",\\\"1187.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_6_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.5000000000_305.0000000000\\\",\\\"1187.5000000000_245.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7\",\"endPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_7_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1202.5000000000_395.0000000000\\\",\\\"1202.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_7_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1202.5000000000_305.0000000000\\\",\\\"1202.5000000000_245.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9\",\"endPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_9_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1232.5000000000_395.0000000000\\\",\\\"1232.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_9_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1232.5000000000_305.0000000000\\\",\\\"1232.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20\",\"endPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_20_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1397.5000000000_395.0000000000\\\",\\\"1397.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_20_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1397.5000000000_305.0000000000\\\",\\\"1397.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19\",\"endPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_19_4\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1382.5000000000_395.0000000000\\\",\\\"1382.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1382.5000000000_305.0000000000\\\",\\\"1382.5000000000_245.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_8_2\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_67\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1217.5000000000_425.0000000000\\\",\\\"1045.0000000000_425.0000000000\\\",\\\"1045.0000000000_357.5000000000\\\",\\\"1007.5019245000_357.5000000000\\\",\\\"1007.5019245000_350.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_10_3\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_66\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1247.5000000000_410.0000000000\\\",\\\"1052.5000000000_410.0000000000\\\",\\\"1052.5000000000_342.5000000000\\\",\\\"992.5019410000_342.5000000000\\\",\\\"992.5019410000_350.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_15_2\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_65\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1322.5000000000_425.0000000000\\\",\\\"1322.5000000000_335.0000000000\\\",\\\"1007.5019245000_335.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_16_3\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_64\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1337.5000000000_410.0000000000\\\",\\\"1337.5000000000_327.5000000000\\\",\\\"992.5019410000_327.5000000000\\\",\\\"992.5019410000_335.0000000000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_17_4\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_63\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1352.5000000000_395.0000000000\\\",\\\"1352.5000000000_320.0000000000\\\",\\\"1007.5019245000_320.0000000000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_18_2\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_62\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1367.5000000000_425.0000000000\\\",\\\"1367.5000000000_312.5000000000\\\",\\\"992.5019410000_312.5000000000\\\",\\\"992.5019410000_320.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg\",\"rawStartPinId\":\"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_2\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"347.5000000000_590.0000000000\\\",\\\"1120.0000000000_590.0000000000\\\",\\\"1120.0000000000_500.0000000000\\\",\\\"1112.5000000000_500.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos\",\"rawStartPinId\":\"pin-type-component_f9130057-4ade-4f7f-a4ec-80702a655d28_1\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_1_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"347.5000000000_575.0000000000\\\",\\\"1112.5000000000_575.0000000000\\\",\\\"1112.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos\",\"rawStartPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_38\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_0_0_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5002460000_515.0000000000\\\",\\\"662.5002460000_545.0000000000\\\",\\\"1097.5000000000_545.0000000000\\\",\\\"1097.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos\",\"rawStartPinId\":\"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_4\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_29_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.6500000000_123.8000000000\\\",\\\"1157.5000000000_123.8000000000\\\",\\\"1157.5000000000_140.0000000000\\\",\\\"1142.5000000000_140.0000000000\\\"]}\"}","{\"color\":\"#e2fe0b\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_3\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_31\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"558.9490360000_99.4268885000\\\",\\\"655.0000000000_99.4268885000\\\",\\\"655.0000000000_230.0000000000\\\",\\\"653.5002565000_230.0000000000\\\"]}\"}","{\"color\":\"#f90158\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_2\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_30\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"558.9490360000_112.4682080000\\\",\\\"640.0000000000_112.4682080000\\\",\\\"640.0000000000_230.0000000000\\\",\\\"638.5002745000_230.0000000000\\\"]}\"}","{\"color\":\"#ed81ef\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_29\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5000000000_125.5095860000\\\",\\\"625.0000000000_125.5095860000\\\",\\\"625.0000000000_230.0000000000\\\",\\\"623.5002925000_230.0000000000\\\"]}\"}","{\"color\":\"#5FAD4E\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_0\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5000000000_140.0000000000\\\",\\\"610.0000000000_140.0000000000\\\",\\\"610.0000000000_230.0000000000\\\",\\\"608.5003105000_230.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_5\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"543.5055910000_33.5261015000\\\",\\\"543.5055910000_27.5000000000\\\",\\\"617.5000000000_27.5000000000\\\",\\\"617.5000000000_72.5000000000\\\",\\\"685.0000000000_72.5000000000\\\",\\\"685.0000000000_125.0000000000\\\",\\\"707.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_4\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_0_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"529.1097235000_34.4258060000\\\",\\\"529.1097235000_42.5000000000\\\",\\\"602.5000000000_42.5000000000\\\",\\\"602.5000000000_87.5000000000\\\",\\\"670.0000000000_87.5000000000\\\",\\\"670.0000000000_140.0000000000\\\",\\\"707.5000000000_140.0000000000\\\"]}\"}","{\"color\":\"#1642b2\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6\",\"endPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_6\",\"rawEndPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"480.5237200000_151.3920860000\\\",\\\"480.5237200000_155.0000000000\\\",\\\"407.5000000000_155.0000000000\\\"]}\"}","{\"color\":\"#ef9cdb\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7\",\"endPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_7\",\"rawEndPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"481.4234845000_138.7957475000\\\",\\\"481.4234845000_140.0020835000\\\",\\\"407.5000000000_140.0020835000\\\"]}\"}","{\"color\":\"#f2681c\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9\",\"endPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_9\",\"rawEndPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"481.4234845000_115.4024795000\\\",\\\"481.4234845000_110.0000000000\\\",\\\"407.5000000000_110.0000000000\\\",\\\"407.5000000000_110.0010410000\\\"]}\"}","{\"color\":\"#cc1212\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10\",\"endPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_10\",\"rawEndPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"482.3231890000_101.9063780000\\\",\\\"482.3231890000_95.0000000000\\\",\\\"452.4115945000_95.0000000000\\\",\\\"452.4115945000_95.0010410000\\\",\\\"407.5000000000_95.0010410000\\\"]}\"}","{\"color\":\"#eed145\",\"startPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8\",\"endPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2\",\"rawStartPinId\":\"pin-type-component_54195fcb-e342-4208-b4ce-f4de03f5d795_8\",\"rawEndPinId\":\"pin-type-component_b466983e-1896-401c-90c5-57535cb2e5a6_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"481.4234845000_127.0991135000\\\",\\\"481.4234845000_125.0000000000\\\",\\\"407.5000000000_125.0000000000\\\",\\\"407.5000000000_124.9979165000\\\"]}\"}","{\"color\":\"#bd684c\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_9_2\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_50.0000000000\\\",\\\"932.5000000000_50.0000000000\\\",\\\"932.5000000000_170.0000000000\\\",\\\"1060.0000000000_170.0000000000\\\",\\\"1060.0000000000_560.0000000000\\\",\\\"752.4980575000_560.0000000000\\\",\\\"752.4980575000_515.0000000000\\\"]}\"}","{\"color\":\"#e94343\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_0_26_0\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_54\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1097.5000000000_80.0000000000\\\",\\\"1022.5000000000_80.0000000000\\\",\\\"1022.5000000000_252.5000000000\\\",\\\"992.5019410000_252.5000000000\\\",\\\"992.5019410000_260.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg\",\"rawStartPinId\":\"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_1\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_28_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.5000000000_-130.0000000000\\\",\\\"1187.5000000000_-115.0000000000\\\",\\\"1127.5000000000_-115.0000000000\\\",\\\"1127.5000000000_-145.0000000000\\\"]}\"}","{\"color\":\"#9caeaa\",\"startPinId\":\"pin-type-breadboard_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_baacc681-4994-4064-8b3a-269f4fbd62a9_1_3_3\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_47\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"752.5000000000_-70.0000000000\\\",\\\"752.5000000000_-62.5000000000\\\",\\\"820.0000000000_-62.5000000000\\\",\\\"820.0000000000_192.5000000000\\\",\\\"737.5001575000_192.5000000000\\\",\\\"737.5001575000_230.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_19_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_-145.0000000000\\\",\\\"1142.5000000000_-167.5000000000\\\",\\\"1382.5000000000_-167.5000000000\\\",\\\"1382.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos\",\"rawStartPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_1_29_polarity-pos\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_18_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1142.5000000000_-130.0000000000\\\",\\\"1157.5000000000_-130.0000000000\\\",\\\"1157.5000000000_-160.0000000000\\\",\\\"1367.5000000000_-160.0000000000\\\",\\\"1367.5000000000_245.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5\",\"endPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg\",\"rawStartPinId\":\"pin-type-component_1c5b82ec-d40c-4873-a511-0cb71ebcb6c9_5\",\"rawEndPinId\":\"pin-type-power-rail_baacc681-4994-4064-8b3a-269f4fbd62a9_0_27_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.6500000000_139.1000000000\\\",\\\"1187.6500000000_155.0000000000\\\",\\\"1112.5000000000_155.0000000000\\\",\\\"1112.5000000000_125.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_25_3\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_23_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1472.5000000000_305.0000000000\\\",\\\"1442.5000000000_305.0000000000\\\",\\\"1442.5000000000_230.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26\",\"endPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_26_2\",\"rawEndPinId\":\"pin-type-power-rail_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_22_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1487.5000000000_320.0000000000\\\",\\\"1427.5000000000_320.0000000000\\\",\\\"1427.5000000000_245.0000000000\\\"]}\"}","{\"color\":\"#e5d545\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_27_1\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_17\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1502.5000000000_335.0000000000\\\",\\\"1420.0000000000_335.0000000000\\\",\\\"1420.0000000000_192.5000000000\\\",\\\"932.5020115000_192.5000000000\\\",\\\"932.5020115000_230.0000000000\\\"]}\"}","{\"color\":\"#8b7d04\",\"startPinId\":\"pin-type-breadboard_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28\",\"endPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_d3e67062-b31b-41bc-8e97-0bb2a0d8f023_1_28_0\",\"rawEndPinId\":\"pin-type-component_e089bc97-3efd-4a29-a939-30b226883bf4_16\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1517.5000000000_350.0000000000\\\",\\\"1412.5000000000_350.0000000000\\\",\\\"1412.5000000000_200.0000000000\\\",\\\"947.4999115000_200.0000000000\\\",\\\"947.4999115000_230.0000000000\\\"]}\"}"],"projectDescription":""}PK
     t$v[               jsons/PK
     t$v[��2��  ��     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino Mega 2560","category":["User Defined"],"userDefined":true,"id":"972688b5-e2a3-1d53-e820-bc24d2f5082a","subtypeDescription":"","subtypePic":"b949fd05-6e10-4256-9d1b-e11f1f9900de.png","fqbn":"arduino:avr:mega","iconPic":"01119c27-1bad-421a-afe4-dfb48490a906.png","imageLocation":"local_cache","componentVersion":15,"pinInfo":{"numDisplayCols":"42.49620","numDisplayRows":"20.99812","pins":[{"uniquePinIdString":"0","positionMil":"3149.60741,99.90612","isAnchorPin":true,"label":"A8"},{"uniquePinIdString":"1","positionMil":"3249.60729,99.90612","isAnchorPin":false,"label":"A9"},{"uniquePinIdString":"2","positionMil":"3349.59328,99.90612","isAnchorPin":false,"label":"A10"},{"uniquePinIdString":"3","positionMil":"3449.62094,99.90612","isAnchorPin":false,"label":"A11"},{"uniquePinIdString":"4","positionMil":"3549.62082,99.90612","isAnchorPin":false,"label":"A12"},{"uniquePinIdString":"5","positionMil":"3649.60682,99.90612","isAnchorPin":false,"label":"A13"},{"uniquePinIdString":"6","positionMil":"3749.60670,99.90612","isAnchorPin":false,"label":"A14"},{"uniquePinIdString":"7","positionMil":"3849.59269,99.90612","isAnchorPin":false,"label":"A15"},{"uniquePinIdString":"8","positionMil":"2249.60846,99.90612","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2349.59446,99.90612","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2449.62212,99.90612","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2549.62200,99.90612","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2649.60799,99.90612","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2749.60788,99.90612","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"2849.59387,99.90612","isAnchorPin":false,"label":"A6"},{"uniquePinIdString":"15","positionMil":"2949.62153,99.90612","isAnchorPin":false,"label":"A7"},{"uniquePinIdString":"16","positionMil":"3649.60682,1999.90612","isAnchorPin":false,"label":"D21"},{"uniquePinIdString":"17","positionMil":"3549.62082,1999.90612","isAnchorPin":false,"label":"D20"},{"uniquePinIdString":"18","positionMil":"3449.62094,1999.90612","isAnchorPin":false,"label":"D19"},{"uniquePinIdString":"19","positionMil":"3349.59328,1999.90612","isAnchorPin":false,"label":"D18"},{"uniquePinIdString":"20","positionMil":"3249.60729,1999.90612","isAnchorPin":false,"label":"D17"},{"uniquePinIdString":"21","positionMil":"3149.60741,1999.90612","isAnchorPin":false,"label":"D16"},{"uniquePinIdString":"22","positionMil":"3049.62141,1999.90612","isAnchorPin":false,"label":"D15"},{"uniquePinIdString":"23","positionMil":"2949.62153,1999.90612","isAnchorPin":false,"label":"D14"},{"uniquePinIdString":"24","positionMil":"989.59606,1999.90612","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"25","positionMil":"1089.60983,1999.90612","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"26","positionMil":"1189.60971,1999.90612","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"27","positionMil":"1289.60959,1999.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"28","positionMil":"1389.60948,1999.90612","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"29","positionMil":"1489.60936,1999.90612","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"30","positionMil":"1589.60924,1999.90612","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"31","positionMil":"1689.60912,1999.90612","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"32","positionMil":"1789.60901,1999.90612","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"33","positionMil":"1889.60889,1999.90612","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"34","positionMil":"1349.60952,99.90612","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"35","positionMil":"1449.60941,99.90612","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"36","positionMil":"1549.62318,99.90612","isAnchorPin":false,"label":"RESET"},{"uniquePinIdString":"37","positionMil":"1649.60917,99.90612","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"38","positionMil":"1749.60905,99.90612","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"39","positionMil":"1849.60893,99.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"40","positionMil":"1949.60882,99.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"41","positionMil":"2049.62259,99.90612","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"42","positionMil":"2749.60788,1999.90612","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"43","positionMil":"2649.60799,1999.90612","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"44","positionMil":"2549.62200,1999.90612","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"45","positionMil":"2449.62212,1999.90612","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"46","positionMil":"2349.59446,1999.90612","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"47","positionMil":"2249.60846,1999.90612","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"48","positionMil":"2149.60858,1999.90612","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"49","positionMil":"2049.62259,1999.90612","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"50","positionMil":"3949.62035,1999.90612","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"51","positionMil":"4049.62024,1999.90612","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"52","positionMil":"3949.62035,1899.90612","isAnchorPin":false,"label":"D22"},{"uniquePinIdString":"53","positionMil":"4049.62024,1899.90612","isAnchorPin":false,"label":"D23"},{"uniquePinIdString":"54","positionMil":"3949.62035,1799.90612","isAnchorPin":false,"label":"D24"},{"uniquePinIdString":"55","positionMil":"4049.62024,1799.90612","isAnchorPin":false,"label":"D25"},{"uniquePinIdString":"56","positionMil":"3949.62035,1699.90612","isAnchorPin":false,"label":"D26"},{"uniquePinIdString":"57","positionMil":"4049.62024,1699.90612","isAnchorPin":false,"label":"D27"},{"uniquePinIdString":"58","positionMil":"3949.62035,1599.90612","isAnchorPin":false,"label":"D28"},{"uniquePinIdString":"59","positionMil":"4049.62024,1599.90612","isAnchorPin":false,"label":"D29"},{"uniquePinIdString":"60","positionMil":"3949.62035,1499.90612","isAnchorPin":false,"label":"D30"},{"uniquePinIdString":"61","positionMil":"4049.62024,1499.90612","isAnchorPin":false,"label":"D31"},{"uniquePinIdString":"62","positionMil":"3949.62035,1399.90612","isAnchorPin":false,"label":"D32"},{"uniquePinIdString":"63","positionMil":"4049.62024,1399.90612","isAnchorPin":false,"label":"D33"},{"uniquePinIdString":"64","positionMil":"3949.62035,1299.90612","isAnchorPin":false,"label":"D34"},{"uniquePinIdString":"65","positionMil":"4049.62024,1299.90612","isAnchorPin":false,"label":"D35"},{"uniquePinIdString":"66","positionMil":"3949.62035,1199.90612","isAnchorPin":false,"label":"D36"},{"uniquePinIdString":"67","positionMil":"4049.62024,1199.90612","isAnchorPin":false,"label":"D37"},{"uniquePinIdString":"68","positionMil":"3949.62035,1099.90612","isAnchorPin":false,"label":"D38"},{"uniquePinIdString":"69","positionMil":"4049.62024,1099.90612","isAnchorPin":false,"label":"D39"},{"uniquePinIdString":"70","positionMil":"3949.62035,999.90612","isAnchorPin":false,"label":"D40"},{"uniquePinIdString":"71","positionMil":"4049.62024,999.90612","isAnchorPin":false,"label":"D41"},{"uniquePinIdString":"72","positionMil":"3949.62035,899.90612","isAnchorPin":false,"label":"D42"},{"uniquePinIdString":"73","positionMil":"4049.62024,899.90612","isAnchorPin":false,"label":"D43"},{"uniquePinIdString":"74","positionMil":"3949.62035,799.90612","isAnchorPin":false,"label":"D44"},{"uniquePinIdString":"75","positionMil":"4049.62024,799.90612","isAnchorPin":false,"label":"D45"},{"uniquePinIdString":"76","positionMil":"3949.62035,699.90612","isAnchorPin":false,"label":"D46"},{"uniquePinIdString":"77","positionMil":"4049.62024,699.90612","isAnchorPin":false,"label":"D47"},{"uniquePinIdString":"78","positionMil":"3949.62035,599.90612","isAnchorPin":false,"label":"D48"},{"uniquePinIdString":"79","positionMil":"4049.62024,599.90612","isAnchorPin":false,"label":"D49"},{"uniquePinIdString":"80","positionMil":"3949.62035,499.90612","isAnchorPin":false,"label":"D50"},{"uniquePinIdString":"81","positionMil":"4049.62024,499.90612","isAnchorPin":false,"label":"D51"},{"uniquePinIdString":"82","positionMil":"3949.62035,399.90612","isAnchorPin":false,"label":"D52"},{"uniquePinIdString":"83","positionMil":"4049.62024,399.90612","isAnchorPin":false,"label":"D53"},{"uniquePinIdString":"84","positionMil":"3949.62035,299.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"85","positionMil":"4049.62024,299.90612","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/05e0cc9a-68eb-4905-ae12-aaf8623b6ed7.svg","propertiesV2":[]},{"subtypeName":"Water Level Sensor","category":["Input"],"userDefined":false,"id":"97784b10-4dcd-a3be-9167-75f1272c8490","subtypeDescription":"","subtypePic":"0657d52a-d145-430e-bb7e-5d1be0618b5b.png","pinInfo":{"numDisplayCols":"7.873610000","numDisplayRows":"24.409700000","pins":[{"uniquePinIdString":"0","positionMil":"278.9027,2373.2617","isAnchorPin":true,"label":"SIG"},{"uniquePinIdString":"1","positionMil":"378.9027,2373.2617","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"478.9027,2373.2617","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"iconPic":"8ade0660-1c92-4b58-a3e7-adda420d3982.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"MB102 Breadboard Power Supply Module 3.3V/5V","category":["User Defined"],"userDefined":true,"id":"307d45d2-aa1f-05de-326e-55c453eb206e","subtypeDescription":"","subtypePic":"fd3ac6b5-800b-45c8-a4ce-2476671127d4.png","iconPic":"915d9337-ea3e-4fec-8caa-7acd53f715e1.png","imageLocation":"local_cache","componentVersion":4,"pinInfo":{"numDisplayCols":"12.59843","numDisplayRows":"20.86614","pins":[{"uniquePinIdString":"0","positionMil":"159.37736,1995.85039","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"159.37736,1895.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"559.37736,1995.85039","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"3","positionMil":"559.37736,1895.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"160.37736,203.85039","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"5","positionMil":"160.37736,101.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"558.58118,203.74848","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"7","positionMil":"558.47927,102.64657","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"8","positionMil":"263.37736,1397.85039","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"9","positionMil":"363.37736,1397.85039","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"10","positionMil":"463.37736,1397.85039","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"11","positionMil":"563.37736,1397.85039","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"12","positionMil":"263.37736,1297.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"13","positionMil":"363.37736,1297.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"463.37736,1297.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"15","positionMil":"563.37736,1297.85039","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"28BYJ-48 Motor Driver","category":["User Defined"],"id":"ecbd5bee-2226-4f1c-8fdb-aaff666e8628","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"00941d67-c746-454a-b945-4fddefc776b2.png","iconPic":"ef87c5cc-d843-475d-a868-97060fb00c54.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"10.89860","pins":[{"uniquePinIdString":"0","positionMil":"841.32961,870.15945","isAnchorPin":true,"label":"IN1"},{"uniquePinIdString":"1","positionMil":"744.72685,870.15945","isAnchorPin":false,"label":"IN2"},{"uniquePinIdString":"2","positionMil":"657.78433,879.81969","isAnchorPin":false,"label":"IN3"},{"uniquePinIdString":"3","positionMil":"570.84220,879.81969","isAnchorPin":false,"label":"IN4"},{"uniquePinIdString":"4","positionMil":"137.50165,680.89094","isAnchorPin":false,"label":"Vcc"},{"uniquePinIdString":"5","positionMil":"131.50362,776.86339","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"917.27685,356.98425","isAnchorPin":false,"label":"blue"},{"uniquePinIdString":"7","positionMil":"833.30126,362.98268","isAnchorPin":false,"label":"pink"},{"uniquePinIdString":"8","positionMil":"755.32370,362.98268","isAnchorPin":false,"label":"yellow"},{"uniquePinIdString":"9","positionMil":"677.34614,362.98268","isAnchorPin":false,"label":"orange"},{"uniquePinIdString":"10","positionMil":"587.37213,368.98071","isAnchorPin":false,"label":"red"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"DC Gear Motor (3-6V)","category":["User Defined"],"userDefined":true,"id":"7115dd0c-9076-1603-96e1-f4f66aa483df","subtypeDescription":"","subtypePic":"e2e2c934-b375-45fc-834c-534243cbf361.png","iconPic":"6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png","imageLocation":"local_cache","componentVersion":7,"pinInfo":{"numDisplayCols":"26.87010","numDisplayRows":"12.94650","pins":[{"uniquePinIdString":"0","positionMil":"119.68733,976.07429","isAnchorPin":true,"label":"V+"},{"uniquePinIdString":"1","positionMil":"119.68733,317.15429","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/7f9ce5f4-cc5c-40e6-be98-a947128d0a84.svg","propertiesV2":[]},{"subtypeName":"LCD Display (16 pin)","category":["User Defined"],"userDefined":true,"id":"23598c1c-7607-4538-b177-9ab948fb1937","subtypeDescription":"","subtypePic":"31959ea2-aec5-42cb-a646-ec7cb3b6e41e.png","pinInfo":{"numDisplayCols":"31.57611","numDisplayRows":"14.25319","pins":[{"uniquePinIdString":"0","positionMil":"318.95833,1322.88889","isAnchorPin":true,"label":"VSS"},{"uniquePinIdString":"1","positionMil":"418.97222,1322.88889","isAnchorPin":false,"label":"VDD"},{"uniquePinIdString":"2","positionMil":"518.95833,1322.88889","isAnchorPin":false,"label":"VO"},{"uniquePinIdString":"3","positionMil":"618.95833,1322.88889","isAnchorPin":false,"label":"RS"},{"uniquePinIdString":"4","positionMil":"718.97222,1322.88889","isAnchorPin":false,"label":"R_W"},{"uniquePinIdString":"5","positionMil":"818.95833,1322.88889","isAnchorPin":false,"label":"E"},{"uniquePinIdString":"6","positionMil":"918.97222,1322.88889","isAnchorPin":false,"label":"DB0"},{"uniquePinIdString":"7","positionMil":"1018.95833,1322.88889","isAnchorPin":false,"label":"DB1"},{"uniquePinIdString":"8","positionMil":"1118.95833,1322.88889","isAnchorPin":false,"label":"DB2"},{"uniquePinIdString":"9","positionMil":"1218.95833,1322.88889","isAnchorPin":false,"label":"DB3"},{"uniquePinIdString":"10","positionMil":"1318.95833,1322.88889","isAnchorPin":false,"label":"DB4"},{"uniquePinIdString":"11","positionMil":"1418.97222,1322.88889","isAnchorPin":false,"label":"DB5"},{"uniquePinIdString":"12","positionMil":"1518.95833,1322.88889","isAnchorPin":false,"label":"DB6"},{"uniquePinIdString":"13","positionMil":"1618.95833,1322.88889","isAnchorPin":false,"label":"DB7"},{"uniquePinIdString":"14","positionMil":"1718.97222,1322.88889","isAnchorPin":false,"label":"A"},{"uniquePinIdString":"15","positionMil":"1818.95833,1322.88889","isAnchorPin":false,"label":"K"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"181","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"ce527fa2-4558-4370-a5e7-21077342728a.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"28BYJ-48 Stepper Motor","category":["Output"],"userDefined":true,"id":"de09217e-3b73-b82d-0145-70b2df9a4b72","subtypeDescription":"","subtypePic":"27b84e47-6648-4cee-a869-6ff1a6fc12fe.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"21.25000","numDisplayRows":"34.37500","pins":[{"uniquePinIdString":"0","positionMil":"862.48611,62.50694","isAnchorPin":true,"label":"BLUE"},{"uniquePinIdString":"1","positionMil":"962.47222,62.50694","isAnchorPin":false,"label":"PINK"},{"uniquePinIdString":"2","positionMil":"1062.50000,62.50694","isAnchorPin":false,"label":"YELLOW"},{"uniquePinIdString":"3","positionMil":"1162.47917,62.50694","isAnchorPin":false,"label":"ORANGE"},{"uniquePinIdString":"4","positionMil":"1262.47917,62.50694","isAnchorPin":false,"label":"RED"}],"pinType":"wired"},"properties":[],"iconPic":"50196d33-890c-4789-8115-a73c306e50dc.png","componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"DS1307 RTC","category":["User Defined"],"id":"9f0127e3-b141-4b6c-b341-c271412e4837","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"f158dbb6-f78a-4fb5-8a82-0ff8626242d4.png","iconPic":"0956fa89-558f-410d-92be-91de6d3dc59e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.07858","numDisplayRows":"8.68668","pins":[{"uniquePinIdString":"0","positionMil":"101.51202,710.31242","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"101.51202,610.31242","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"2","positionMil":"101.51202,510.31242","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"3","positionMil":"101.51202,410.31242","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"4","positionMil":"101.51202,310.31242","isAnchorPin":false,"label":"SQW"}],"pinType":"wired"},"properties":[],"propertiesV2":[{"version":2,"id":"initTime","label":"Initial Time","description":"Initial time of the RTC: \"0\", \"now\", or a valid ISO 8601 date string","units":"","type":"string","value":"now","displayFormat":"input","showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED Two Pin (Blue) ","category":["User Defined"],"id":"117aab52-1b06-40f5-98b6-df63a601b0e6","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"2c98734f-75db-43ce-800c-ea69461525e8.png","iconPic":"d4c851cf-9fb5-43cd-809f-e1699313b4d2.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/1f9f88e9-950f-4940-ab85-21b1c84421ad.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33334","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33371","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18643","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"LED Two Pin (Red)","category":["User Defined"],"id":"5f0a7f7f-5908-4e39-94d8-2714a0462581","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"3d0a314b-f708-4b2c-819f-35c414b123ec.png","iconPic":"6608fa58-7afa-4488-b64c-2b761d69d6bd.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/a9e23d57-c0ac-465e-ae7a-a15cecbcb7b3.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"4.24452","numDisplayRows":"5.30565","pins":[{"uniquePinIdString":"0","positionMil":"161.90689,79.96916","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"261.90689,79.96916","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"DHT11 Humitidy and Temperature Sensor","category":["User Defined"],"userDefined":true,"id":"a76bb123-3d3c-417d-b1f3-c8417efb7bc7","subtypeDescription":"","subtypePic":"779eddd4-9cc6-4216-b155-89a4f50be07b.png","iconPic":"44e1934a-57d6-434e-9b76-9cc9cf9f98cc.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"7.00000","numDisplayRows":"10.00000","pins":[{"uniquePinIdString":"0","positionMil":"200.00001,100.00056","isAnchorPin":true,"label":"VDD"},{"uniquePinIdString":"1","positionMil":"300.00001,100.00056","isAnchorPin":false,"label":"DATA"},{"uniquePinIdString":"2","positionMil":"400.00001,100.00056","isAnchorPin":false,"label":"NULL"},{"uniquePinIdString":"3","positionMil":"500.00001,100.00056","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"componentVersion":1,"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED Two Pin (Green)","category":["User Defined"],"id":"a70bb5a8-99ed-4f1b-882e-eac0873b75ef","componentVersion":5,"userDefined":true,"subtypeDescription":"","subtypePic":"f9728bc6-2422-4ead-9082-90351081a874.png","iconPic":"9ba3df0f-d630-43f7-8169-617793654d93.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/3749fe76-cef7-4b42-9f27-525b8a44301e.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33333","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33333","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18606","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Pushbutton","category":["User Defined"],"userDefined":true,"id":"232ac546-6e45-4194-9a27-0fa614949a21","subtypeDescription":"","subtypePic":"e2a053a3-24a6-43e1-ac97-395cbc045e87.png","pinInfo":{"numDisplayCols":"2.45180","numDisplayRows":"3.30020","pins":[{"uniquePinIdString":"0","positionMil":"221.06000,315.00000","isAnchorPin":true,"label":"Pin 3 (out)"},{"uniquePinIdString":"1","positionMil":"221.06000,15.00000","isAnchorPin":false,"label":"Pin 4 (out)"},{"uniquePinIdString":"2","positionMil":"21.06000,315.00000","isAnchorPin":false,"label":"Pin 1 (in)"},{"uniquePinIdString":"3","positionMil":"21.06000,15.00000","isAnchorPin":false,"label":"Pin 2 (in)"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"PTS645SL50-2 LFS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"C&K Components","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"6b551873-9f16-48c5-b1b9-2fc6ab10f815.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Trimmer Potentiometer","category":["User Defined"],"userDefined":true,"id":"cc03c8ee-909a-4085-863c-ededb100351c","subtypeDescription":"","subtypePic":"b9037746-96b4-41bf-a651-5749520ed4a9.png","pinInfo":{"pins":[{"uniquePinIdString":"0","positionMil":"23.60000,20.00000","isAnchorPin":true,"label":"leg1"},{"uniquePinIdString":"1","positionMil":"123.60000,310.00000","isAnchorPin":false,"label":"wiper"},{"uniquePinIdString":"2","positionMil":"223.60000,20.00000","isAnchorPin":false,"label":"leg2"}],"numDisplayCols":"2.47200","numDisplayRows":"3.30000","pinType":"wired"},"properties":[{"type":"dropdown","name":"Resistance","value":"10000","options":["100","1000","10000","100000","1000000"],"showOnComp":false,"required":true}],"iconPic":"ded7c6f2-b589-43f4-a4a7-c3e3242414e5.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Pushbutton","category":["User Defined"],"userDefined":true,"id":"232ac546-6e45-4194-9a27-0fa614949a21","subtypeDescription":"","subtypePic":"e2a053a3-24a6-43e1-ac97-395cbc045e87.png","pinInfo":{"numDisplayCols":"2.45180","numDisplayRows":"3.30020","pins":[{"uniquePinIdString":"0","positionMil":"221.06000,315.00000","isAnchorPin":true,"label":"Pin 3 (out)"},{"uniquePinIdString":"1","positionMil":"221.06000,15.00000","isAnchorPin":false,"label":"Pin 4 (out)"},{"uniquePinIdString":"2","positionMil":"21.06000,315.00000","isAnchorPin":false,"label":"Pin 1 (in)"},{"uniquePinIdString":"3","positionMil":"21.06000,15.00000","isAnchorPin":false,"label":"Pin 2 (in)"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"PTS645SL50-2 LFS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"C&K Components","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"6b551873-9f16-48c5-b1b9-2fc6ab10f815.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LED Two Pin (Yellow) ","category":["User Defined"],"id":"1310de1e-180e-4aed-a1c6-f80032a2bfde","componentVersion":4,"userDefined":true,"subtypeDescription":"","subtypePic":"42e39361-2f02-4030-a678-a3271aadd3f6.png","iconPic":"a4af1710-95e2-4b5e-9600-8e4d90487313.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/e51a5bd5-4abe-4a22-abdb-307c464150b2.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33334","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33359","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18631","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"L293D H-Bridge","category":["User Defined"],"userDefined":true,"id":"155f7657-2d2d-eaf2-280f-5c76a41d0679","subtypeDescription":"","subtypePic":"022fab5a-d187-48c2-96d7-20ad2a5d1671.png","iconPic":"39d025b2-988a-45cd-b457-87e73cc458ec.png","imageLocation":"local_cache","componentVersion":1,"pinInfo":{"numDisplayCols":"8.00000","numDisplayRows":"3.30000","pins":[{"uniquePinIdString":"0","positionMil":"50.00000,21.69999","isAnchorPin":true,"label":"Enable 1"},{"uniquePinIdString":"1","positionMil":"50.00000,308.30001","isAnchorPin":false,"label":"+V"},{"uniquePinIdString":"2","positionMil":"750.00001,21.69999","isAnchorPin":false,"label":"+Vmotor"},{"uniquePinIdString":"3","positionMil":"750.00001,308.30001","isAnchorPin":false,"label":"Enable 2"},{"uniquePinIdString":"4","positionMil":"150.00000,21.69999","isAnchorPin":false,"label":"In 1"},{"uniquePinIdString":"5","positionMil":"150.00000,308.30001","isAnchorPin":false,"label":"In 4"},{"uniquePinIdString":"6","positionMil":"250.00000,21.69999","isAnchorPin":false,"label":"Out 1 ( Controlled by Enable 1 )"},{"uniquePinIdString":"7","positionMil":"250.00000,308.30001","isAnchorPin":false,"label":"Out 4 ( Controlled by Enable 2 )"},{"uniquePinIdString":"8","positionMil":"350.00000,21.69999","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"9","positionMil":"350.00000,308.30001","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"10","positionMil":"450.00001,21.69999","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"11","positionMil":"450.00001,308.30001","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"12","positionMil":"550.00001,21.69999","isAnchorPin":false,"label":"Out 2 ( Controlled by Enable 1 )"},{"uniquePinIdString":"13","positionMil":"550.00001,308.30001","isAnchorPin":false,"label":"Out 3 ( Controlled by Enable 2 )"},{"uniquePinIdString":"14","positionMil":"650.00001,21.69999","isAnchorPin":false,"label":"In 2"},{"uniquePinIdString":"15","positionMil":"650.00001,308.30001","isAnchorPin":false,"label":"In 3"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     t$v[               images/PK
     t$v[z|S�wq wq /   images/b949fd05-6e10-4256-9d1b-e11f1f9900de.png�PNG

   IHDR  	�  �   �]A�   	pHYs  \F  \F�CA  ��IDATx���`[�������cK��{oH�0�����y��$6��6��EK���i���Reo({�Bd�v����{�Md��I�XwH�~@�$�W��{u|��O�$	�E�?�t�:R��t��p��bHCI�             a�!r[��sq�`<%+w���D�])�Z���y���MUw            H`J)1����}�`<!0%�<��ϕ�)            ���3�}pUp��^���1��/             ��xE��ɞ2�����U"-            �1 ����y�ܟȪx�u�             ͳ?ܗ�oϜ�A�#�Gu�zFyi�fc�Ի            @�(���@N��}���[�O./�x�lC&            �(#�/��1��ʇ�ƃP            `�}�`a6?1�\+            p��#��Cz5����k
u�����l�����7�0��~u�X��* �G�ϖU��B�/���ZN�98,�t��            �k`��r��Mz����+!�6�WZUS���}�R��ܤ�t
f���F�ߧ䃵�	�9�p_,#��*�ϟ�D�	            <�&���Zw�Ǆ�o��+���{�лf��&��c��h�.X.���s����{�2��fO��)��x�%;K:[X!�>\"O/Z}�G�U�`�@����F�           ��T��ʍ��zT?���T�^�Q��].�G�|�=)��>��]q� �kIe�<�t�D��'����[�@�}�:��D2�GG�tX_����(�}��`ld(��{��            ~��t�/#%Y.�[�-Xq�ǟԳ��m�Һ����RQS���������EC{�i}��{k6�Q��b�>�&+w�yJ�P           @�x�����B�d���'<b���Q�Gs�	�z	���ġG�i��b	�>��g�o4�           @����E��㎓���H��A�zwQ��MKN�K�����ٹWl(��z$�}�}2R�#�+���&�Bb\,            �$���ʳdP�6�2#U��Wʊ����W���_K�0���^��
��1��<~������>�a}$��b]��eQ]����!�B �nW�Q<�p_, �[�$���J            xRj�_�5��v��Aٵ�uߢM;�G^��{��ٯ��św�q]���O(x�Si,����j�a��Q]���2ک�@doy�Q��>�#�[(%g            <���V���kY�}�lܻ/�7�s;�|D?i�"]Ftm'����rf�d{Iy��xt�r+�׽U@N��E>X������̒q}�X��X��!�c�E�w��O��]:ggEq�����`�2B            �9�~�\f��@ʪj�?o�
��k�߯�`�Ⱥdg��.9U��߯5��'�X%��h��%�����]u� ��zM����W���?��ē'pI��}�>�"�[(Q            ��nW�!�W\Y-���%y��+dh��r��r���ˎFF�+�����Z'�=��\<�����uaA�����ix�Ͼ���W��"�}��[�O���}            �-U�!�������Z#�س���tm��գ��`_��d�dXk�?����W�l��_���PX�e����`�.�*�)5�T ����l�W�a�2��R��U|�R��C�r#�g~Q�J��qYKeH7�g��?�߼o�y_k         ptc��Zm(c�2��E��D���b#$�a�$��h��F�|\�y�g����?�O)�!��`w��Y-��w�l�-�%��ל0�.�w���u������uJ~��ɯ*�9�!���!�|��a�,  ����<���;�zgϬ�-�Y^��3�|����3Dg�'         Аa�6D�Qo�E�S:s��c^�ԩIYe٣T�7^����8�\n���Eʷُ���C>.l��r�٣��^��G�l/.�K�������YY/$�S�C����}�"؇�3T�O$$  {�'J�%��HѦN�ȓWD��ݛ�����/sd�?ҲK��6��:�Y/5��Hm         �U"�1�e�}^�M���b�M�-�X�]~������K��%g�Q�����Rw}����>v��+�γF[kz�����E���b}���1F���x0���ʴ��!� @�0D6��gH�߷ϸ���'�vSe�ȋ�[M�ѹ���C�j��          q�2�#���Y�{�~�������/}�ʙ�OI�.��P�"钝%?>u�u���F>�f�a���"�p�f9�w��	e�}A@=��ӋVb��`  g����ř{џ�)qa�O񛛙3��~I�lj2?         Ĺ�"�Ҥ��3x�%3'�T�Z�L���;�@���5���?�����/eٶ]}��~�$�{�eF�u���K�a����g˭`_�V뢽�t�WFg`C��iy]E�  �2j̃���V&�|���J�Jgޡ���i}眹��н���         �!a�G�)�)%�N�]$��;�M�۳�̛��9��s�uY)~���IC�KAq���Uh��R��ҿ}+�̬{��u��o|֤�>�t��w��uS�jL�"����Ϙ�W�c� �A�y�l����7e�x���&n5�\��;�?��U)�E         �g��n.�/���&�1���#�je�|�z��]ƶ�Rk�����!�ºhWi�<���{{�T�BMZ��v��%��1C�����6�Rʐ?s���9�  ��T��9ť�w��ֈǕ̸�嬟�9NՄ�e�<_b����Y��s=������7%Z�g���q��g�zW�}�d�Ϛ���d�:�z�C��K���k�����/�%Z�g�Ȩ��?'Z�N��=E{��I{e��h�7��+�<���Τ���굅a<0B�n�/�B<�x��y�����֘��w4?�h�9��K�V�߮�����ooy�|�u����RU۴@_}?a��z{�u���Z�~"^0r��� ���۫�gN~Cb�~�<��0�;�.��o�#:���ߢt��]�^���׼�W��O��w%Z���\��-��M���d��"l_�Q�}��y��^�g����O���jd�◚�'�Y�e���z����Y{$���D����5/�K�߰R�d䥒(|�_�B���h��D����>^8�H�z���h��R{e���x����a)C��h�䧽0�nS����2u��`i�_�U�T��v4?�qO�u��Ҫj�*-�A_�!A�v'��}�_�Y>_�߫�5��Ba�[ur���T�<P��J���JF�s�>  <�<Y�`��s�:��)�h��!����aCS����yf�?;bi]��z���7�o�ߚ_/�     	�0
�ϘP4}�b�EӦ��ܝ����'��ET�۫����ky���Z9�4h>��?��P��B��{���@�  �"˒��y{�8y�ĸ�铞Ϟ�?!���RA         <�0�����7�H�+�1鑬���J��(��p�dx����17��'���C�  �,U)ɧ���{%NΚ�^`�_�m�h.K          �1dM�/����n+�8Q2s�K�S��7�xM�J�VJ)C��ͫ*�1���#� �{�׆C��;)nB}�y?NɿD��y@�*         �G��U)߹���'�����Ϳ�0�Q�`3e����@n^*#�E/`  �`;#tny^�6�SE�&�șu�5o�         �*C���	��o�Z�T�I/s�dV��UM [1r�]� �4C���]S<}�Z�s�3���<�j��\          W�O��O^*q�h���y�̫�#�ق`  3�L+�~��� �2��2P��$��x         \bjfьI�K�(*I�fU�Q'
`;��s�yB�/:� � C���=��D2mZ8iʌ�Cʿ�<�k+         �����4�nI$�Zcܑ����J�� �cZ�h"� �C�

ݢ�n�`���ݒ=e��O=��:�!�pH����[�a����m���m���?~�_�,���A��R[[�ט���)��<��-�n�����S��y��[��y��[�]oTR�3|7렛$����r��1���0���Q9W`Zި!� �c���r�K�*�5��@���c���x�p8,���RQQ!^ԡCGk�e_�f���E�T�>j׮�u2-��?�7�t�^ܾ>�Oڶm��m�0�g�^5_��W^�����L���/*((�ޛ�B�^��&���;�mѢ�u�"�m�`�U�Q���Kh��G�?{
�6����h�=ƌ��&~)	�8s��`i���=h�xHJJ��~Zuu�x�ޗ�ٶx�^���-2��4���}H8�I~�0�W��{m�z��=�O�h�㺴;��=e����r��ee�ɽ:7�o閝�~W�1/sd��ҭUఏ������j)�����*�ZX*�Q�dŠ���_�VQY���r�p������$����{k6����C>~L���1��������$|��f��w�N��.k��ٴ�D����r�$4e�U�İ��r�$))Y���S�}H۾}sݒ�z��!����υ:v�d�[UUUԖ��z��ա����o��ٟ�r��}u��޾Z"m_͋�j���(�3�U����`��TV�;w�Zg����!״���.7����:�ؾёh�F·eN�z��J4��Ϟ@{��Ϟ@��QI{�	^=�0D6�V&�Fٴiac�(_�����yF�.]d��͞{�Jӗ��D�]���y�^�+++�b�O#��\��p��R��Mh�{7?�_yrѪcZ�/'�$�9��A�/�P g�yB�խ���3G5�k���r�˼y�0��	��gjBaYQ�[�l�!7n�ז-�e���W� ��8^�A��.Y��D�_��d����>k����C����F�EC{t�{]_���ǧ'����2C�|� ��'SeΤ襘b����
��?�Dnrk�.�t�'''�6zξpA�gꍄd��0E�^��o"���ؾ��g�ot$y,���o����st%%X{�5^�̉tj�%���Z��7���b�.�u���&�J�7\��7�*ٟ]E��UI{�*/o(C~�s�m�����&~��ڼz�x���nz���2�v�ջ/�g�}�A���у�)ؗ��*��-���)��� �y�{J��t�U�\�X��'�:��.׍l�D������¨��/~v�yf񚨍t�f늳�>%��'�5'כq~�V�����y�^;C}^S8[or����ؾv�T#�h����3�=�����t�8թ�h���+�g$���B����Q������^%�Dk��xCc�:�z�A{��+�У�g������귆/�=�Αx�W�nv��"�S�����}�*�����>]�kˬ����{#�KZR��)��u;h�W-���������->��=g`�G���;�����7�DO�|É��o.$:�;�6�V`)�>i]07_�ts=���+��N�
"�S�S�{a
����޾N�dh���h�l��uN"��"���q�S�z��t�nw�Q����Y�W�&�gg�^٫��IG�?ۋ��,�o�iӼ1,�κ}I0'�Qr�x��a7�B}���D�/�p߱H�ww��*kCRm^i)VXMOQ��7>;�e\3jP��%��.+:�׎\w=6�Q���y��7(j����˹��O�?#%Y����'t�`^�˙��KZræ��a}d���K�V��,<��f�j�y��cZ�ڰ��������R^]#HT�΢��|
� �3�(W�}���n�
"�S(�3�m�R�l_��[���L;9�ف؟�G{��+���^y�[�9nuj�5���j��}�ꬣ^gP�3h�`�gg�^9��Ig�?;����o"�-2�*4����?��in�ݜ�E�[�S����!�̮,�y�?G�;�Hx�P�
��x�붞���7?3O\���:��]���~�U��F4{�Ze��y�z��~w�F�����{Y�wlc=�M;��\:�XXQu�����E��p}�vs�z�`��rƟ Yi)u�풝%/��;rz��V��hT��cUEM���?��ʐ�;Nf��@��y�O�x�����e�l��^'�n�
"�S���`��G�?;���>l_��^�����8�9�v��ӝ9n��������733S�P��uT항

�9���^�W��J��Ys*�U��u핽
b�xC�<�mڭ�^I͘�^ '�k�TO�(��nn��"�^%>s
L��Z<����E�0�[��.ا�O۫��_��I?{m������˛�6D%�w����Zoz�'�Xe��	�iz��h��ƞ�J������ҵ���dh��u��̔�W�-�{�yId�_"Oi� ��n^��GK�*����Կ�3�y����N�)�*�p"\�P�7���k؟����ګ�S��ɩ��tjP�=���S�����p_���k��B}n�b���#��u*�W��u�ڣ F�7|���P*o�y���aN����P_�S��b�G)��%0e��;<�}���d�νҷmK����6)ا�Ž|䀺�O~�Rj�F0�O�[VU#/~�NjCa+X�G�Ӿ7�����ֈ{N[��P.��3���WJ���u��5��5��k˿�D��`�5r����7�tƓ�8^��� �(�1i��Q>���!���n�:L�Gq���'�ۥKWOu��pA(Tf[��;w�X��n_�՛h���z��tr�ϴW��δW�Gwn�6�HJJ��ƨW�]��׌�Nw� ]�޽{m�X�b�EEEV��^�Wwjlٲ%��gګ�I�����n�y���z��k������,����^EO2�'����ޙ�>�,8X�g<�+O�4�~��իm��ljjJ] �:w�,k׮��|A��v�7y����wn0gv���>`����_��u��a}���ޓ���'���S�f���~�\F�z������dH�6u�_�j�5Z�����r��a����T�phoyʼ�z����|�{�r��#�%r�O����w��W�{������K����9��&��5�!θmC 7���صk��޽ۖe�`���ٳGv��i˲;u�,^�����v`����z��}i��ǋ��^E���+V��e��`0(^�ے�˗۲l�֛H�W��vm����Kvv�x����l�2[�=p�@	�%�W�3��
��׮�j�G������l_��L����*:���"%�U=2��Q%�MY��_o^�%W\\,k֬�e������z3)�M�@���:�g�������z�iy�����B��q���[�R~~�I��)�HI�K���G>;���u����WO���`�������k�-W���n�/\Q���t�n���;�Z��]=j`�}'��,�[dÞbIT��.��?�J~p�m���$w�5Zr�yG�81���~G�3�>         �%t����T�<�C�#�wX������{k7��~ݬ�׌t�`_��k�و�>��'<Ғ����n���7�+b���j��߾�u���]�k�,ٴ�D��7�ig�!~�T��7X�K�Ӯ3X������"A0�6�F�/8<}Re�D         ���pHj�޾~��6�}�D��GO�	��أ��k����1W?@�|��Y������5�!��eFZ����P����/\)S�O�SJ�>a�����-_m�)�J+LC||����G��t(�,�)�O�n�iy�>�D�e���|�~�gΤ����BUj�?E         �(1V�μc������*Y O ��(�}@=/~�N�+�%��/e��ʴWO�]=���r_[���.���:\s�4��z��ݳ��Ⱥ�����6N\��w��m2a���i�R ���B�餡���j�֣1���m�82�)eDg�8W:g��`N�n��Z         �f2DV
�h���́��R%*S / �w�}@=�5�����r�C��:����>>hļ�u������Ei�N�L9�O׺�+v˗[w�8=m�������vo�Szw��n�8�l�i�TW��g}9}�7�Y�P�
+�d�;��FX�ń�䪇^�7ÐU�&Rz�ӓ         h&%��5�2��_m��F
���}ٹyF��K�#���W��:ZXS�rC��\So��%��֪��?V׍T7
��.�A���`_d���� [}�2��ws?X,7�&��>�pޠ�2�wg�p�AS�04�!�Z�        @(��L)��])�}�%>�Pe��I�������m�f�^�*�kGn�KKN��׷��_���P���k\X#F�C�����/~�NJ*�%k�����#w=��5�����S��ܚ�K�H�3��\�����~~�r�ܧ��'�VA�(16Y��         ���&A��6�KO"�g!�4�+�Nգ������WZ�/��
�E<� :�����Ez��ݞ�n�l-*=��+jj���k����FLON���'���+qCJ������P�C}+
v�W|sL�[n�b�ß,���:�n�ܫ��=��A�A"~��D�T��         ���{j*C��E��`�=���;ɚ75�/���/��_b}/��m�a�Ң��r��90�����?���u+���w#AȦX�y����%�U�B���?���N�}��`���j�5:#�a�r��D���         �Z�T�$���t�W��<�G�hĶ�Ryo�&߯�u[�t��k�,קK���<:����t�T�z4>=��|�~�l�S,�[��'t� :���Q
�V��E�/Q評'�~���ں=�c�tx_yf�jA�	�����0����        ��RR�Y��|������8�G�8�y����un+C;����������E���\�=��5�n��K�6�M�ُ�o��i׎(��8_�6�s������#�����屛.�����(/,]+�� �)I7�R��          g����5�} D^�r�UTI0=պ���=g`��￺�룚n�p��wl����䫎iYW?P���Ԅ��e�$���mܷt�N��^]�^>�f����Ѻ��z���w�P�}�BU���QF�        @4TW��M_���x�"�BemH�]�Fn<q�u�N*�~_���5����)t��mf��3����Ց����$���}z$A4��^�H^��w�n�u�hy|�J�������k"eH�\         �����k"% �E�8�yV�����4�o����f� �6=�������lp���Z�[�Yи�m����t�nw
f��c�ɜw���8ah2�	         �C��8�̠O�0�}�a|�a��ٹW��m���'�X)���Ou�ÂW?��a�|���ewY�Q-��S��-�IVZ�u��=�}V�@��M'�a��6�o��+}�~���rf����R6e�	�0��ƕpH���l�:3`         �n�&Qbt��<�`p�-X!�<���=� :��=����ʨ��`�6ykձ��G�ꄁ�u=-�ζy��{u�?\zZ��*jj%�F�;�%[v�sK��e��Z�[e��m�������&Q����         �#�O�$���+�� �"����3K���6C6�)�ʲ��p�g�>�e=�xu]�O�S�����������������'���Dpd�{��hho+������x�A�0�`_S)~W         �C�{jC���ǈ}�w��@O)��/W�ԧG���£���M���B�f�[���o%��w������$�tx_�Ѹ�2�s�������������4�������n�HM���;⃡���#j�;�lLjZ	         J)�隠�O�kU� �,�}�K�T��~_����n�%�Ǽ��pX�[�Fn;��kFlR�oh�6r�C�_͂i��&3]���^uh�`����IO�%�q��>�K;��c�X忳P��WJ,���O�
s_HK���4+�(J����T�X�a           :���ۖΙ�SpH���B/�m� ��r�{���F<�hU�`�w������@ʫk�sg��n]���v���˳�mp`����X���/c6ط��T�p��v�HA�Q~�7N5�� 8�����         �������'�F?�y� ���A��v���ڐ����f/���d�b��*`��JK������?_!�6��������E���\�Yo/�����KX�B���)         @T��B����B��4�}���p��7V|#ŕ��^����ūe���}�Q�)�WQS+%�:�TU[_��]$K�씥[w���;dWi� :v�Uȟ�_$?;g� �(Q�/S����SwCjx�A)%�{��=zز���4�]oϞ=�[�n�,ߋ����K�w?�j�ī�ڵ}����Kq�����4�+7�^E�׶���QϞ=lYvjj�x�^��={ضl�a�Fw�^���5�l_�%��M4��ѓJ{�D۾i��Q]�װ}���X`(9��W�!8H�Y�R=%�l�R���o˲[�Ȑ�Jo�تU+����Ȑ�*oՋ�#؇��i�w̶m���|��Oz�m�b�i�|d]�G��a]��?�.^���=��_����~�{_�Ժ �(���U<c��A�F�Z�{�=@��>)��ζ�y������V�F���J���U�l�b��+����ګ�+�������2�K��55Ւ��;7<q�+���׫;s<rHO�QV[[#���z+++l����JRRR<S/�Ut��^�Av�W5�Ϯ����Z������*z�כ̵�}�S
����uJKK����|���H����JJJl�WתkFl � ��̓}PL��J�z�M�:ٵ@ �zg;����jv��Eؾ��^�P�;h������ݩ�g�n۟G�����%n��zw��e�󔖖Hff��9�k�u���U&��q�Vo�qr�r��<굇��g�������o4���`�Ae�������ꫮn�̇G��n���߉��۟'�W/��@�  {]%S��!Ӧ��C�rg�1O���Nv�G���N��s�^'F��/��u�ڏz�C{e?�}9թ�vg����ݙC���^gQ���v�x�^��~��l/�u�_{����qEǩ�O�6��rA���٧�_z��9�p;ܧ�u"�A�/v� �V�m�����!у�:>�Mq{��d�p���z��V�N�d"ؾ��^�P��h��C�o�;5"��r�^�:s�����u��o8�ׯ3؟�A������o��,+��_����|r�x�ӡ����raa����V���b�>  ��n�:��2mZb���ug^_	�ss�}7;�#��l�^�9]�[!���}��y�k�+�%z�ϭN��;�ܮ����u��Ө��}E��J�zM9��rz��(��rP����k�r�+Gy�xøK�N��ٵ�	�1�81�	nO�}(n��"���W��}n׫�}����4�84�}  دW�����"�	D��=��k��N�':۩�=N��vH&��}���>�+�$j���N��:��R�S�//��D�U9��+m�:U�۝��W��r�ω�^9����ծ]�So9��+��������^s��,ium��C1�=J���s;���}���n����R������ � %�_��<+�n���rʜ�a#|�[�^�d��t����D}�^�׎p�J��땐LD�����|��>ګ�I���E^	�D��Y�N��D���L9��Uvo_��WN��N��g4G9�\e����]�����]�W�rk��0�������ι��J��R�\��M䙐[�~?M�+��z	�y�>  ��T�@I�O�E�I�2Tȗ?G�r��Ë����@(G� ���y��h����a�D۾�>!m�@�W%X{E��A{-h�z��:5"��܈.�uZE$Z����h+���M�z�ھ^m��^�+�r�y�]�_�+o��Qt��^y�7(���i�zF��I���	�����_�O<���̓�YE�}�d��B}:ܧG*��� �!J��Y9s+�9q�$�`�����in=����w��!��z�[�՛��$l��E���O{�7F��u�֒�V�W����2h�'��9��^�7�o|3؟�$*7���y��'/���u�m���1��4/�2��������כ���z�|�  p�JU*�\�ę��!I ����
��\}
%ί=���Bl߸E��͠��k�3��'�[]�ߨ7�Qo|K�z���9�Qo|���F�8"%IFX= ��?N�ջ�*dݙ�7R�����D��ph� p�uZ���_�L�D1ujRm�1O)�F          7(Ȭ�}���(&槪�<��xo�d GD�  ǩ{9y�gN~C@���oD�q         �H)#'�3k~��)�I��̪G
��D�  �)�)�G��5��)�$�r�2��%         ��2�<��?�h�E�Sf�*b�H �,�}  �B�U!y�e����μc�ġ`���"��$         <@�
��eݙwJ�}��H�Ιu������]�  p�R�K�H~)�������G�y��xά1U          /Q��/$/��=o\����%���7#��H� �i�  p�R2L���̙~^���̝u�a�sfmY         x����$�8�μs�e�>=R_X�ǕRi �� �mJ
Id�9�<i��JbX0g֥b��8Y         ��)�z��|�ɟP4s�"�a���7b�M��/f  <�<i�B�aV���Jf���Ě�S}���?3+��(�	   EF3^�s����@���^�Q�}��y�T�R����!o-��:�z�C�΋�zG�����x7���������Xs��Ɂ��{��j� �+�  �
�Z�$��y�0��4�y�������K��������h%����Y��#�3��	O�i'k+3�M�V�f�c�����l_G9Y�f��*پN�^�P�������?Ys�wT��>�&���=3�GF�H��9��u�|�)�+���7�x�L�+�<E{��_��Y��w&�m�Po4)Q�'�9y�d�[7�ʭ��2gzװ�xܬ�dw� �)�<o�ۃ�Ǉ&ͺ�4�
������Ws�;I{���uI�V�;f���}���7�o�'���ר7��U�ʺ$�D���5ē�h���U|{�㫸����R�K����97�M�\<�Pٹ�ׇE�4o�с8E�  /Rj�?I�s���䯺g�}?-iuW~�P��;C�:�<5T:         p̔����4���hHjsJgޱK<$+gN?����u� �k�  �,��G�	�]���mQ�ʴi�n�Q�ܹ풤fJmH&)��         �7J|�?����s��yL�H����J�\��Y=�������Z�� ��>  <N)�f~�?P������tU���w�9�z��ڐ�!F���
e0F         �R���W������7R�sK��U����3�.Q����d�:�� #�R]�/�+$������C�G
7v|E��"d�N�GZ���"���s�5� '
         H0J�V"�����s�_W��~r��
;�.���-���r1��E��uG!�> ��  Ƙ��z
����m���a�z;��{k�}����rʟ����3�/�Eg�'	�u�
         $2%)�>߅%����+�x�
��7/g�1/w�Ԕ���c¡�x�I�KM�I @�#� @3�;���h~��6�@N���*�[+Q+�R�����H�-�*5$Fց=����|\?�z?%���J��Y�$         8$�Z*���+���~	��*1V�>:1�UJT��Qb�>��oHr(�2�o?�!����!�U���#U����W�`  q�<��n~їs�����<SPa��*>��Խ���         p��H���h��h���ה������=�A�}u F�             �1CT�t�h���}             ���"���RUU%^��nQ[�����B���ŋ�ᰴh�B��             8�s�βe�υ�t����$��>=^�.]d��͞���!)++#��1�             ��k�H��.^��B!)//x�>             ��J���P_�W�}����`            �ߧ�M�t)����ڐ 6�p��a7�B}n���y�>            ąkG�_L8Y�geHEM�<��W�˗>���X�V��0�RZZ*Ns�^B}��`            b�w��'�⬺���I��q�IzJ�Lz�mAlp:��V�/��z	���}            �y��1����5X�ewY� 68vs;��T���b�>            ļ~�Z5z�ߧ�W� ����n�W���
{�[jj�TUU�Wt��Y֮]+���,?%%E���S/��`            b�O�C~��������e͚5�,�_�~����P�>ZXXh���п?���S/��`              B�            pI����H�ʚZ�^Rn}=Vz`��L	��Hyu���˫	��C� �Ӳp��T���Ł�R�t�Z��F�B�⦽��JuJ���㓰�ݱ^$טg�;������L        ��t��	�{ʄA�dt�����Z��Pؐ����/V�?>�JJ*���գu�\�����dD�v���R���PXo�!�}�B�-XN��!��"!���M��0.�P [
K�n�1�pvfں�pX^�r�aӻM��ܶ�}��m�]�������j%�#n,�M{K�pt�|��Q]����?���\&�#��+iW���Ր�[�˺��$�����k��,*�uܶRV>K*S2�{��ʀ�oJjU�������b�ل�         ��O��Ni����O��Nm��-���y�5�löC.��kΓ��w��'�}2�{�r��ar�#����{���ۊ�����ɠ�߆I��߯�Ӌ��M<}�\8���렇��p���>�����lp߽�j]�կ.+�uiWw����.�/\y؟)���kF��|�{m��r�C/�z������������\+ ��P��Đޫ>�5��P���!��M��}z�>������J����         �>Т.�W
��ˢ�;d[Q�$��rB��r���V��Kv�<w�r��ɧ�4��h./���V>3�t�N�QZ.��Irr��rZ���s��Z^��w�?=%kv� �FO+�Q�2��F�Ӯ=H�{�3k�]��SM|�M���k�����t�P��]����w��B}U�!k�N�$/��"��y)�aW��
�}���V����_)�֔ ��vay��&        h�ͅ%�����}�Lv�<���hލZS�����^u���㿥6nty�w�?\*�-\��Խ'��$��p���L��-�%���r�ܧ����
x��Oh�{���Y2�wyw�&Gק��L~���r��ϩ���KN�����\x��|����������߫1�/`#/��"��y1��p�WC}:�7�7d9ᾘ6�c�lx_9�Ok�ߴ$��Wֆd�����-�����d�  @��)%�Z���U���R     ����g�nW�a�Y�m�\��d~�Ւ��K�6�2�Oyg�ƃ���;�j�k��C���r��^�W~�]�ů_��V �w��
4���^�d�O��C���E��ȫ��1=БƦ����u����i�߾\�=��`����+墡��)�JK�9W�)���s�=H��&���u�?�f������^�ED3��k�'��ED+���P_D2ᾘ��o~�8�o��)��~czt�.S�8A���k�������E v��Ӑ�mep���4"�2Ҭ��mSYu�UT�ƽ����Y�i��W�H�j��.m23doy������7y/�GN���]���Z�m�-/~�V6�)L�K����4Bz��1�e|�nһm�d������5���M��O����7I>���ʨ{�,)��E�g-R�e��7X���������lC;��F��^R&˶��m�}��~�7l�k;d����}����}W�M���5��u�Sh^V�6����/.���   ]S�t�q��,g�7����m�"4u���o��v���?�O��6zW�F�U5�����~�[����c��Vu��h��7���i�mݾpho�M��>ϱ����2�{Gk�`�~��Nj|$����z꾟<�����苅P_D4�}V��p�Ă��b%�A�/����~pq�/4�؜7��u,s�?^�> v�h!��>R.޷��G���Z�Z�:����Xq�>r�9c��p�������'��ҵu��OX��T�KFL=�dy`������I�D��͗X����;����Gt�/^� ����o�� [1�����S� L}�~�����t����|$s�_$�`d��V�2�w+ �߻г��E2�f����|�@9��v: ����zM?l���w��K��%���#�[��z���{�]-rὶc�>+C.�ך�+=9I���k7˻k66���å�Y��;K+����x��u��Y�[3���?�ˆwn'?=g��i�ө����תjCf��������˭;   ����ꝯ�-��u�3�� �6zV�fԠ�_��z���sO�n�7,�;�_��tѶ��B&?��̻�º�~}�)֧���*<��56ﴗ?��}��hN�/�B}�P_�ءG�x��K�N��9�ܒ5�نٰ�H�*�E�HO��-2�[�`H/��&�n���Er��G�r$ ���㬠Zz���=�#3��գZ#R����V����Դ�t�����_ן/9O�#}���g�k�]n�X�=��ON!m2ӭ�q0�	�<���KO�ז��B~��$��9���=�
�ꑞ�M{���j�;�~o�w������ɋn;�|�'���E����&�s�I�3~T���FpA_���R�������A�gn��P�e���O.�=���Ƕ/��u��Ow�����)/��Ӳ����Z7�4D~{�8��Z}��׮�Oy�m���#��cw��m�x�3����]|����a�5�PtPϴr��^r��%��Km8,   �m=[����J�6�.���? ���ߔ�o>F�,�-_m�e}b�����wut�ύ`��ʲ�ִ�W?�n��^u�\0��C�����|�T D_,��"�%��������j�/�p_l���S�B}��!���˿>]f �����S_��

������}��T+ q��_ ����Q�������#li:���ϖ[mڈ��dP�6��)k��)�O�a���5�x�j���n��N����a��(2��*`�w�e��G_o5/'օ�^_���:�UZa���G��#�k��y����th��� �E�f���Vxrc�L�{r���W=]����@'t�`g#t�:�G��#��0���wi+׎l�����=F�^�Q>��cr�^�����>�`�^��3Gt�����n;L�jk��9U�����>Z�z	�N"����%�rޟ���!��pq�#�j���ȍ�I�=j�FB}:Խpc�5���O5���k'ȅ}ڳ����Y�����t�Q���h��B�uh��^u��P��-;�Mۭ)����jÆ�>�>��?�۸VHs�yѯ���Ѹ㤳���W� �  ��dg՝�k͝%G�����}=��g�0��u���;]������M{K���[el�}��1C:��Bn���w�s]"S��أ��z�q��ix��z
�3/`�X�EM�/�C}M��z�/�
���.7�%��=�M=5�V
�wxN>Z��I?����Q�t'�ۓ��:��1��EA�Ly	����P���_���}�����0ҁ�Q�y�ONa���?X�?�|˼�Z�:�w�C��Ғ�����\y����ŋt�P5ě��[��~��W�m������2aо�mO�i��ӡ��F�ٗ�i�n9e8��F�Ф��R�N#����_&�6R�^�Q]��
�y}��C���6�C_���Mcr�<�.䥧%��TeMm��|n���aǻ�m�,��c��U�(�F��i����߽�����k뽋��z�C�r��}��f���eɖ�5z����.�>0(�G�"=����G��5��/�i����ij��v}۶��f���������[���S�t�}����ٻ�(έ��xB<�� ��ݡ�B��R�W��[���u�
-�P��!�G��qw7�=o��"�ldv����_&�͔��ʼ���{�.��~2w������A�������R���������v�B�KC<2�G��I_�@�e����������:+�/��+�~�g    ��L������iM^��+W��	p��F  M��
 1K����rH����uE��-Г��y���j~��ôm�\Ek���;n(]����;���m� M��>9U�}��S��z��b�{/�iK�ON���:�7�*u�y���������P9ԧ�'#<��������A����
 h���W��������׸�/����7y+х}{���d����@p��-�s��+�JN|���k�z��p�h�Wg��mY��F���G\����ؖ+�u^�_Jc<]i~O��I���p���,L�^���m���x }����q��mWo���x����ly��~m�7��Ә��<�p���u�p���'��K'KZ��K��k�5,��A`�	s�V��r�<�q���וߗN!����?z�Cmk頪14>�_�[���x��g牱�w��<^�t��{¹��e졽O-��9)�����g��K�7��)�21�7&���|�q�-�;ꋶ�\+}���8�:s�V��B�ŕU�;q��_���,��#� �   �����]1>�yy�q�&��D5yր?;J�= Ԅ`��p;%�R�|A�[��m�)Z���*x��=�f���_��Ќ/�Z<�&~�QѮ���<X�[ Z�47m
����ӦP���];rO�O�B}rUᾃ�I���	���տ���\	���q� � ��
4#���南n�����.Ҙ�#�D�O�fZ=��^:��"E;����<���\���q�hߵ(Q����P�߄�f���6[KTS�CDZ6��ǟ>�w�Fz��*�ӽ=˸�!��o7R2i������k������53��w7�P�վ��B��)�㓃}|�v�WD�${v_y[[w�F�O��ܦ#4���h�+�=��*�?��B��	V)��-��_Z"��<J_�P��򊆏���ա�;x#�F�O���DXJ^��K�{C]ch�Ί�IseF@s0NJa8�����&�����C}�?�s��#a���&�c�_��y�AT>.4ɍw��]�RS𘰼�􏧮4)ԧ���>9H��-:��ߑ'8    ����jG?,��(��ڎjU��Ɋ�O!��T�'��+� @���� #sf�������H�������'��L��#��������B];Y����؉6E<\[^��s[��$OC}r����1�'ww��C}=C��������V�۱�y��j��v��vE�`��41��  ���ڂ���+��XE���>~��k�J����J��q�sWǕ����i7ږl:�	`��f��������'�O�s?%�~���'�8���V��2/{kzw�pю�Xx�8��-;?W%����[�*3��DȢ�����d�y���1i��i_]��HXl�����_��P!$v䥭���yc�1˕��9�q����_̔Z�r�Qy�J��s10���C~.r%�i��M�yZ^�xB-��%�w����E2��
���עi�[hۊ9�b�#r8y��%������ܱ��l�|��k�    4Go�N���9��w<�cu@H��7�����4E���v�� ����y�x���{���'���_(���{�i��/�?���yj����k����w��}}�)I�h�����q��KD ��A6�1Z��p_���t�g2�G_ ��|�p�{t E{!h[� ;wK��_De�� �h  ��Z)��i� _'S��3����>��X���6R��x��B{�R��fPU(�9t�o>�:vQ�x2W�Zԯ��}�� N��E���|��U�
�����<X���Q�c��5�OQzn)��cfx�q��%�I�+��NT�w.ǧ*&0ڙK.���H�"���#���4��#�~q	}�2}���V��6U:����
�Zz���ݒ��<�}GJcXГQ�JGPBM�q+�xb�����I��������V�ң�sg�wY3���,�:    ���֒����8g��L���d��7�ݑ�<6[1����3���� ��> ��J.J�3w�D���/>�|&�/�6o�p6&I�x����@W�v=9OQQ���?�>�  j�S�>*`u�]u!Z�������K�rPKҭh�)u���!ܢ\EJy�  M��3W�S�G�;���K��̔�tekj"�`_vQ�b��4�:�R�e+3J�ɯs�ʏմ ���������Ӣ�1��8<%���/��O�z����IJ�����xh����mj��M�/aD���-z��P�[�2nY�%��[Ct�Z&d�*2�<���j����cI|�n�F�,/.
�1�]��x�.�j�d���;��������/$-���3��')Q~uPn�Q��4�-�s�\Q�r�����Tzx�>��m-[����Tέ�|����o��LR��s�3	��>��D��JۚX��    ��|�������\���m'����n����٢*9���y�u 4�} �tP���s�z����r���q����@\9�-����ha��`��w���sт  @�̕*�(J�*G)4bn$�ߍ�Ս��X�����RJ�v����A?[�q��v֢R����[%�TPZ.�ᰔ,
IJ��q��C�"Ӳ�Ƹ���ШgQ��J�\=���P�����TZ!���,��re������O�*�����&&]Յ��w4*��-Ov���l��qK^�-���K=��{@���9��e�h�[�i|��z&�>�5R<�6_��u)_pxe� ��!U�qR������������U�z���Zҙ�����ڤ����~����>�PT�|s�)E�MS)W߳7�H�AGG��W���؈��ES�B�V�#W+3�ڻ+���Z�f7I]Pb�g�#�
���A��{����l���ύ�/>��g��� 盓����{~|�f�   �#��ɓr�?�o�F�l<��q;_g[��W^�����} ��> 	�21�i��*�O�/�c�qu>~��k�`[:�7}}�b��x��������ށ�c 	  @ڔۙ5�E���;�͍T�Xޚ���]D�!�ԕ��OWRiGPD�
&�^�C���qџ/�q��ǓW4����
L�l�P���S@'#�E5U�2a �v�D�E������>4�Fvs���7IW�~~l?���]1�W��\<Q(I��\��J���$��I���h�0��Lp������&o�TB�����	9�:_��M�l{yFx����G��W�덅���9����\TG��M�N�
��5�7��#=>�O,s0"��}TAn-7R2��=���gEh�'�����&5�>w�z����igE'_\B���۷]	ϓ�O_�y}�� 7ڸ|�:u��8R��%��,�׃^��?ZT�7~�ƓbcjLc����snO�O,LUZ��g���"�:6�U��[4A\��V��5����ܔ:~��q0~�w0��}�bl���V�B�7K��(Rۿ�YT^Y)B����1�ϭS��,�k�D�<��љ" .e��i"����=K;�Mֆ/��q���!��ڡg�G�����רN�#ٹ˼�����dW�y��zoc�5   ����O�Ut��);wr��z��ׇ��7?6[q�Jv��֮� �	�> 	�A*�h,��r����s�hg�Ve��c��Z_��ǆ�*~��8�   ҦwW0�Y׭�Z���*�zh:���O�X��N��J�<�����|Q����i�wW���ɇd�{{З��*.�);vK�t�J!�^\���/�q�vܦ����9������I�������#�������g��]��V!4b��KS{u��d�!�i��.�>����l[�T���w'.׺����2nO�Q � �^��ӏ�#d|\v�d�d|v�<�,uv��'ο��Ŋʌ\=n|wQ!^~��!h��,��mm��}����C�d��w�Z<QT�;K�Rhu@�X���+{|�)������G���D��E��rw��O̭�~oGՂ���[Z�M����h�7��ӣ��듇�0#|������3%U��e�Q�:�_��ymv�D��*�e�������P,{}�*���tT7W1)�1�/�p;��-ow[+�!u|��q%bm��ы�����N��?�;�ޝ>��E@56+��s���R|v��+�Y�?߻Y�Q_��[+WK�����e    ���s|�ڹ�|d���e����f�ù��+�)Ɓ���;��� ��} ����mx7\����l�pC��ԫ̓}��W)�hS   ��m-�?2�F�GWX��_��t������lQ����\Q���?�?����n;�Y��h�ҩb�ká��/,��7�AA�|9�����/�^�K��̪�z��@n7�{�J����Bp[>�?�9�ܬ�D�S���دg��&x��[}��Mm��=��wyҔ+�p�����@_�����v�o�.����' �[m�%�o�A-O�-�92�m���cA_O�3�5����Ն�?�)�p�g��S�M���96�����zݸ%{}-װ0�/��z�F�����s������{ϐ&��*�}�����*U��3����������gSt�{�'6W���ھb.�r�fUQeWe�W^��+�i;���i;�-;W����
V�Ý�dD<-�c�$�e    ����X���;|�=���&����O�Wt��ɟ�o:J�����hc��Lyp*<5KL6d˕p�h�HEՅy~��ڎ�b=    ��A�J^��������x��ա�>��b_W;QQya��0���簢e-�@� W��4��pK�C7n��ph��E�>������E��[p؋/��l���ɭ@3����q7����� 
MJWy�,El�?җ=V��	U���m?!*(>?��8v���?��L�����~~nl�&�wKs[�3�מ��<zfL���럋7��m���!��l�n�}�T�|��4�rq�f����+{=�n��rd�U��.?9T����U��ږ�yR�s�n����q%,�Ŗ��ZRM�f��L��̑"���}Hq�uy��^6�3[Sq�4��ڧ#H���F��S���Ǉ��oA��@�*;Ƨ����>>G|敲��^Ο��m����%}���J	_��*,�����!/�����������ˣh��pIo+   @{�]v>1�����G�ci�ݢ@Sp���+�(B}�/\�g7њτVVVԣG�Y�����J�c���un��l{K4�} m�R���I�>.��]�O�!��2r���F�G[% h<G;��݉�KԿЛ_�G�撔9;X�OoG*.�S{]y����8�2W�N��ӎ����^W�l{/H|{A}!o=B�J���"�z%\����EŲgF���g�n9�U�r�Z�r����#�W�c�d���O�@���.qAW��}ȶyJ�.���&S�㹵'H�_Ƴxy�����F��C9o�:Eۃn�
>|^���~��q��g�Ka��0_��U��x�_��ȡS���{@�"�[���Lza�Q�:~��p���5��#u�hLI��}�]$~��:�j��4Z���.�;�	���W���j��2�����W�����(Z9rKG�L�����TPRJ��Ų�M�h}�m!K4$ ����Ͷ.��s���"M�v�M�^8��TW��4��	�����N�&f{%�����ωꄌ�Қ���c�~�.��&z��-U���h�dh~�����^{9XS7��v��j*��fl�OE�e��8�ϛ��t#%CTx�z�    ��+y%m>G�q�mHPB�p�yW~v�6�<��ǔ��?���q�g�1r)����>���۲�nn��CR�޶�`@2��U���[6���5�ҁ���&���!_�IE�Mo�RXT@i""�I@:z���ˎ�B+����!�����.�j������t5�6����i�M����8���XU)�?2������g*�hƾ8z�F�O_Կ��**�p�Fj�}\�l~uKEn���P㶜��%Z��g�(Q��)C����Oi���-���|��9Z�*&�ܤP����#���ӆ�@7G�
$�	a���ᆗ�S|ϕ45�-fcp���*��9�ƕ�Au\��Zx��7�n��Ŏ���s�&>/puv1�}~�_"nR�����a���9D m�CP   @;YU�?3�]��K�������;�Yw}P5o�!@)��rȭ���u���-,,�ל�����Z�kn^E�O3 �І�{wev���-�� h,���xPpp��}�KIϣ�RFG���v��PjR�/��Cn������5���֢@���Z��s�Ɉ�+O�@F`L��`�^�?Hs:"A�̍��ʜb3�S���W>@ĭ�k/�� Q�l���E��7@�����m*����[
������*qX��}�<q�0�t��n�� hI�>�-;    �;[Sc�ىz�[�ʹ\ݘ'
s&���
��)&#Gt�	�����;@ki�������m��i��[kn�<���>� ��{5�:���E�  ����дp������+(ѡ��$Q��C�	�5u{�ueۛ�q������j����b9>�����A9no��� ]r^�b�+�I)�ggv����mȑ�[��ם�ϣ3E;VnI���K��8�q��큱���yn���Z�)�       @�p�<?Ozl�/rw$]�ƿy��R\
�>,&�VTb�g�w��u}��&m�ڡ>9s��}�٭[�����>̀�z�6�daJc=��g���'��h�I�Y>K���=��g� �L���=($4�JJ+||^�f���Dح�=_ץҲ��WXJ��	"䦉�������������\�\R^^���w���~��rk[�I����b�B�����x���v���lQ���~�r�<Մ��<پ����o]��N�~n�}�>�N�hw+5�6S�����)��~n���     �%�yk_�9���<�@W�R�)(!�r�����]�wu���t�j'�5�@w�ŉ�����0��'�����,(�Фt1&q4<V��hwksZ�l�Wi,�w���G������� @}mr�33�jS�Zᾶ�^����>�6����5f}��I��R����	��s�0�q�nt��- h*n���hM�i��O��&M�|��ꐃ�%��&5�ش���5j{3K�U��ѡ>4��Uʶ�ѿ�h��r5��[$��ˬ�b�rc�Ӟ�I�9?m�-���|�y���7%���dy����B�9Y�JC��L˦��"�&����e�j�����e^���O    �vq�2��d���x��~�K�啕t4,�>� B~ �:;��ǉ�+񩴡��C��ϛ�iD�Q}鑡>�`������IAIm�N�
l��t���}O/�N�Ɗ��VT��z�Yyb\�;z0k��h,�&�v���ՎL�}=l�г�h֪������:�&��>�4��Ӳ�>�l/�}҆`@���Y�g�/�7y}���`���  4^_W;��׽��m���^�6��Qb��'�zr�fP��t�Nϡ�7�H���f�x,�����fZ�|�Ϟʕ�T��Df��F�V����&}ҕx;n��3۷�X�q�v�O��b׆���1�D5���-�׶����Q"��*ޥ���ҧsǐ�����߲�V�F�V    ����o���U,?��嗴�߆��L+�����<Wg媑�\h�C���ذ���d瞓zva�g72m��\����#���Pz~]�O粚ԅ�+�����9B'"���U�B{k� �/!'_#Bnr<6����*��Ɓ����~���]���s�$U\x��%���[���ɡs��j�0(_�D��������!��_�L#?����� �^I%�&gn^U����}R�^����>�6�'�];Y*��g����M����i� ��N�y�H��..  h#C�ݵj��Ah�&���'*���^um`����ͺ�����IJ��ɍ�1kxLw7�ֈg�*81�f��J;��+�����|؋��r�ζ���{����.6�biF=<]\08Gb�����J��&zdkj"�}]�i��k�s���P     @���h#&�����ϒ���1�����j}������g��ѝIrEe���I%����R����?,�(7щ��&x��;S��y����aH���I��t�>���n�N�k]xd.��E=�IOW�"R�D�Ty����Eӽ=jt��ȡO^��g��ߤ����+狀�\J^�؟ܖ�K'�61R��W�5:O�l�h���p�\~~�p<u�hL_�@R4��E�����e�ʁ>9�-�݈�/揥�{�*��{u] �q�r��p_s�u�.YR�^�qW7�� ��ҁ�j|��J�Z���b�Y�O������¾������O��l����Y��Ĝ|   ���M�;;6:�V�՟�xv}�g��-�}ܮu�_7�x)�Q�#9�����v��'�u4�b����i;ns3�-�i�,�v�$~�liFK����
��).�     4��g�R������=��ǹP*�>�s�q=��sǈ	L�=f�~����[_~�!2�}=y3��so��{e�@zc��zC���j�D�ő^�|T��?qYt��I�]|.�������~t,<�֝�&*ʗhx�������AS��=;ӓ��Ч��ω��9����]-"�X�t�hQ�r�{$y��A���J��w��s1I����ř>�9���ڋ�a'#����~�������0_��}g�0���I�dǁ�L��E|�n+�>��P�2������4ɫ39Z�Ҕv��������f�Z1��neeM�4CC#�k.��^�f�^P�} ��?���V�g�.7�km6_	S�؃��U
���)�`k��)>�  h��^��攡-��o�_�-W�I
8�7��C��s���J�����RT<c�Q�$E{C���q��c�}�ci�4��ʹk�<q�A�x�˞�H�gn*h�VU�l=..:� mII��㓿�DO���G�����?}w⒨���`6     ���\�)|��Tv[<�KL�Q��o���V��R8_�ixR��Ț��\%���[4��Mt���A!��6��������hWz4<���,س�XoOH�J���di&Zx��_��9�ձ�$e��#D�U>���!&�qy�1�Pȷ���v���nw6Z�.r��g���>��6i0����篋���P?_C��E@����A1����^�v���_��\���kv�S]�����M�n3mX>��y��W�ѩ�16�c2�n;A���_:U��EGd�i����XU�ג2D�u���HXl��6���'�e>���J+@c�� �m��he���QƚKp_�KU{�ۮܤO��gX/�ɂ��]MP�   ���;S���pfk���QK���yqk���DD�X�MRt).�~�����hebDY�ō^�]��j���`��K�y�j;��5{�m]��٤	�������%�Չ�z���_���Xu4����Y�챙Et3-[T�;v��D%��     ��tw�u}4s�=?��P����EQݍ۵��S�����M��]W������s��|��wBa�zm�	qMH����8~���a�W&���_���'rź���.��oцV^����P��o|�r�aM�6�����;��+ح���R}d�7�v�D�M"��Wn�`�Zu�
WW*����|�����x
�ޗ��w�͘�T���MG�m�!��6��7&}���SL��ju�ъ�~�fmN�d�}�J��^UD���'TO�4�G�  ��Y Z��z�����7�e��E%t4,�F�=�]݆`   @K��L��IW���́�}����@�x �dD��     H	O>�[x���s����U�|�+�I��UUE{9q���M�꬘��ݏ^�O���-��T�$�g\���s|�K~�Aڎߌ7{3��Ǔܻ�>����7�ײ�����H�N2�V����\�z�������?�gј���i������/&�)����SW�~���	���C�}���I�ku����Z���g�QXJ����!W��N]�>�������Sv\r8�9�ps��n  ��`�K�>_�l���hu�?��M�R����ǌ�j���>/n   �Yx��9>'�w�����h       ڻ��zR�[�T���*g��_r�S2H�py�!����ϕ�oe��h򀕔8Y���)�����tv_���v���1ʸ���a��igEC�:iT�OYJ^��X���+4��3=8����h7��@߸j���m�Zjp'��6�'�X"{N����hmil(�#�t�j��[/{�:q�[�S?��[j̪�����;9ť�����; p�MnO��,5\���rUɷ��7v�Rk}��{��mv6FZ�E @�!�     b �)-Z��Z��S��L�n��:�[}D'      @{�-W9���:�X�e|*�����4�i���7w����.mHyukϢ�2�RE^IUp�POz�3�*�u�ݴ53_��sTj�ʹ�3Q	"���%��÷Wd�=�k]<��"��8�򄁔��O��	&)q��`Ǖ����I�e-���,�~u�`g��o�!7)�_�������k �*�Fw���������2����A�)B�O��+&(��/@����Ĉ�۟��W|_TVN[.����ӭ��d�	  ��}   I())%C�>��̘�s�����
244k�q�f(;��Y�R���Z������-���5q�����D�x����EkU�      ����D��:�r�X�Ý��u���n��=��ǹ��3�&<5K|554a����PWW|�b�1��MG#^�;�YTZ�}%�o���2�����6�+.�5gCĭ��5�?�'-؋:�J/�%��@_|M�Ϋ�1<ޕ�_(�Y*��Տ�h`@R��.^�\,�hJ���/4�������=㖼��6�,�Pz��5��[�ѯL����Is�<)�V�G%�m��̥��2E���@OT6��������hd72��U���8&K��^]h��  �	�>   �Gjj:UT萡�Q��uur��
���,�T)��TY�';	o����Ft�ҙ�HS%�����&������<����j�ϾzЊ=?��h����<'Ɂ����/�@+G�՘�΃���D?��R�Lem���ut�����$�۫����    �4���e��|>o��\������6�*�o� w�?Sn��ˢU��e]]��SR�H��cH����O\�q�|�v�� #=�{�)����Z|զ�q`��=���gij�b\��Bz)ע��C=��x�˫љ6�N���p�J��IoN"����&�}���k}�.N�����\���1��ꪇ��W�l�/��1�/�U�R��Ύ��X����9��_3[h ��!�   5p�����Q���Z5P���>����x�g��lN�eK�	�ix{���$�RM�ަ⁜��x7�8�T�O��j�����=1�O��,�-�KJ��3�����b&v{�ǲi4��]T(��p5i��M�q�n��G>a{�͟N�D���    ���Wo�����!�L�=����%b�'.i]��G��?���;�`���ٚVM�L��xʾk�TXZF&���A�7$��6m�FoO*�t�/�p�2���َFz���Uڄ'���o����0������RKm�>(�����^T���<н*0�J;��v#%��^�I�z����YH�e����[��G:::�=��4��]���1���v{�u��>��&�k^�+������R��ʠ�8�w4����9���[�R1�>���ϯ�  �:�   ������\��WM
�%��Piq5�޻;�CJHԜJv�1����D�����r���&�1[�g0sh�(���       �^�Y���2}1�h��������ՄTj/��!�e�gZ�$�{�L��x#Op�`&�5�ۮ'��c�1I�~�0�{@0=6̗ޓ�gnɻ: DTH�۰�����)"Tā��W���h�J	��>�Lˇ��}�ᬑ���5�g��ߘ<D,g��2n1�A����,����FR�▣���I�;9����i�Lj�6�\y�6�}�)���=~��N��#ZCO��L��E�]�2ʕ�-3�o�l�a�X�s�fj&]�K�}��1�;Q���?��󛎪�>'[:���  ��>   �	����D���m�K� �KM/�Rrk��ѝ��3݊�ER��P��b{;��Ɛ���#a�-���ƇH�bJ�.��̑bPK����֝��u-�    @::�XPg���MQ*;w	MJ�-����!]p{W�f�
W��}���?���?yY�'-Q�e�q��6�� ��
tq�o�p?���Ҝh���+��٘��biF{�^@�nܢ�o��l��۟��Z��?�7���_v�d�Rye��7�Å*�-�c 1G��Kۓ����?w4�����>z��g\=�ߗf�v�'3��}gD;���!#==��\�콧�ý0������ER���)�m�oM��>�>�Xx,=��P���_�8�x� =���_�.nچä�r˯��Nv  ��>   ���B:z�yx@�Ļ�$�dɶ�f����JILL�c�ͳ��J�js��q��U�tv�wg�_��9�3(���@Q��     ��tu��eSh��5���r�!q.��f�v���D��U�u~��J��~B�c0P;�p�e�0�v�x��dI/��/�4uU�����lqk����E1+�������--�}�}h��=�䞝ōq��B�@W �
~u�N����DR�?4��|�A,K��jsኌ�?K��=J|��խ���~&�֟�N/�H�Vf�ټ1������%��z�Y�hY��^n{+U܍c�{������F�����X��Ɏ��q)"��P��}/�W�_���1��ц�uuĤm  ��   ��WRL|��	ZVVN1�)�^��U�����t��MDs������q���Ӓm     �ቑ~��c&��j�D:+U���@?�7Q�c\�,8!���h.��7����ԡ�b����Z9���yEF�r�bMP\VN�~�!�/�3mY�)��e�����M����!�$UR�[{���r���>9�O��sպ�U6Y�����#B|�����ުh�9��c�	0�Y�'��`���.u���kI��  U�     �+_7��[�2�;�D��=#.8h��,'��^���1�33��"L����^    �7X�jxs�E{��I���p�D�h��}�)�%\�4��^�q��\	�o�'/q~��+�9B.\�����f?W{���"Ҳ��W=/�����~}]�����I�v��5�z�E�笼���d�$�؎�n5���Ͽ�_����mw�H���=�wW���l�V��[M�+�j�	  M�`     �8O7�g�,ъA�J|*}�/����"     ����Ѭ�XqyE�5O�����p_��\�}\���&М���%�����6�K�Ң~=?�@�Kc�������e�Q���dal(Z���SAi%��6��x��*�]�'gЄo6�9��� �驹b|������R%ˎGv#Y�j}a)���?  ��     �y�[�jn<�z�f�����jG����嵁�(������̤F�/)'��&��LqS��+�b�9     �*�=~I���X4�:�>vQ�*%q�w���1���ҲA���shɫ����Ίh>�d�jV������C�c���D/w�7�H%et-9���FQT�j���oK���od�a�V�{�$R�-��7�  � �v��Ҍt:P�(*+��|�w �~O��+.��i�W���1�J��ꁚ7w��=!�u�opg'zw�p�|�z���}ws�0��{7˺x�T�}م�U���D�>_'^����}hXWg��,��r+����U�'Ґ.N$U�����&�Q��C%��   �~䗔���i��D�Cu�$���ϓ&����>�9����%/h�v7���X��Q�h�b8��M,_�O�mA{h���1��˦�:������l0���_�L�����q�˶��  М� �v�PO�ł}eh����5�su�3.���%�������k*���l=QX�^���˶�[���v4h��-�����ʛ�ަih�   �5��I����h�?��S^YI�l<L������wCK^�F�V�f�T����'���i�H*߿/m=F��	&�nJ�ߗ��_��Ԙ��'�RO�Z����@��]�i�{("�A  �6�     �p+�^�|�E��䤂g�sK/��lK�eۭ͂RiA_O���܉.�j�����¾w���ooP;�^   h���/Z�q������y��J�D��wCK^   �}8s�"�ǡ�ף�8������J��}<Ax��i�/��8  @kC�     (2=[ܴW8��q�%m���|��H�)�����ζ   ڟ��rzj�!���Q9����G.�&iL޻�%�v�bcA_.'�W��B��Eh����髴/4�@{p������ϲ����M9Y���A��2waZ�Ǟ�^Sh��}6w��u25�]+�Ѣ�vJj3�6���nG����|kN�m{A=�    @�q5>U����R�p��*U&�}�N9���o{�^   h���/�Wi��>��=Mm���-x�ڍ�F���*�wGh���'�Wۘ�+�������o���˟9_kP�td<����N��:��'Y�����}����g���di*�3
�(��� ԡ��O%%%�&E�e�MLL�m}T\\,�����M	��>     h7��J臓�E���r�/�=�v/���P�D��e��51��N��3�5e{����~��xn��}�Oi�   �~���M�ٹQ-y5��ۍl�{7n��� o��\�&��eo�l��
g ͽ���b�_s��.������Z�Ղ�?~���q<��غ���[@O��+�_6=6����M��cIqu��7�&z���l��x���L�!�I�2~�Cv��z�~��ʶ���T��᜝�)!!Ara7����5k�O�����TZ*�`,W,((@�Ob�    �v��]��m]%e$uo���6�&lo{;�  �}��O�?D��V�%o{k�{�g��#a�ВZW#[u�$�4���x��4�Ӎ~\�~���iU@'9�@T���}�&� ��d��G��I���C7n�&�ҫ�Y6����DDxrl7{q{l��2��0����䡾����"�pW��PH�}            i����g���d-y5���j�����ց�~ގj�   w�O�P����{FT�{c�2�ӥ��A����6�R��ԉ�<8M����jeF���/��9�ʿ�6��k�P��T�}�I�}     �0�����Ս�L:�x�cܛޟ1��u��֬��     �}���:S7ۺ[8jb^k#z{��f]'WO{``/ZJ�68���0�f[���!I�r�4����
��Z���.9YH�ܰ�δbx;ڿJ;8[���ܿ�����+����ؿR�ʫ��t4&]]�'|z(P��x\���?�F���OQ�9$u�.�����̥������@�F�>3��	K3��ա/�#s#���%hmݦ��B}rm�"�'e�    �`kjL?<CTw�/)��_���qFzzd��#����P
K�$      uqKާ6�ݒW[𲾮�djh�����	��6�feNs��S{���X�EOʞ����؉�_ZBR�fݾ�o\֝�î�zv�����lK'��~�*7+�v��<wG�ʷ��q��S/Jw��H���[;QXUv+-����-B��/�J_�HR6���쳆�X����n�ԼB�����3������ܘ�ą9�ȟM8 ��*��ڡ>���^��4�}      �0v���wv�St�z�M�tt�Q}��MG	     �9����N_��k���sMm��ne�L���i��ZB��E�gnmɡ-�.��i�j~��OPB�ڿJJ�ywmT���:}�Jd�7>�7V�_�0��l���b��'k������ӥ����Id��G�N$����4����U��'

����fb�^��4�}     w��1<Q�}zJU!��?��;gt��1�no�	x���!����U�?\-��ݍ�.��{�\?O����bp     �9��/��;� wG�=����yJ�Z��E�e����Ϊ�W�Wt��L�C7b�Z���)��GR�W\J19Ե�%���-��5/h�*��{&*�^�Qk}R߿�^96+�ܭͩ��M�ڗj����!�ע�Z��yGZ9�I?9d��Ƃ���~���I�x���C�铃�DU��XB��e�����f)��,�ml�hGP�h���љdb�Oύ�';t���'k��h-���J}m��6ĭ�k�#4�}     �P��,n��v��H�fU[��U*��T��r�K���ݾ?qY�̍hxWg:v�      �O����Գ9����ŵ��d��=��4���D5��Rߑ��:��	���9&����+5[5rkK)�W��`�\z�����۪�z���-i7���}���;����L�rv���_o�N��1޿�����\�k����t�z-�S����I��_k�z6]�
����K&I:�'�N�-Pi��dD<��emZ>Ktw�cWOW�^�v�>hv�������Y���~�U�S���ݼy����[d���m�uC�@�     ����by_�z��YHR�����1p�G�     �_��I��r\���vO��8���lG����u���S�`x�U8y|Ajn�*�_�o]ʂd�s���X�mV'�WTzg��Kr�f��f��z�g�&��,�nb��Y�`_QY��󷐤�3A�\ݒ�65=���J���8��]|-Yz�(9����щ4s�VںbY��c�|Ew��7%��֡C���a�����Iz�$�^3��=<IWW:�C�    �ګ�N�ۻN�Ⱥ�JZ�T���-�s(*=[����͈�,쓯      ��(����I��Վ\�����H�7�f/�QTF�XS�x����4�$U�����L���֞�l���"(�������%���ݸ*c?W{rn/�������y=R޿�bl��5�h ��I�U�6�M�E�>�2�
g��im[1G<��M�t��W	  Z�}     �x&.��#��F�kRNA��S~��~       ڛ��T�b>N�D{Cm��'n����V�'nƑ6������+Pr������������mO���kv�@4��3��R�w�y���v<1OL�^2��h�-���DLવ)y��+  �}     @�Z1�6\Yp��p
��$�K��|�nf�i�       �-��lߪִ���
�%��ӻ{�Ų���V��kk�V�����I&h{�孥���N�/%�@�������hx�byq�F�ص����fڹr.9Z�� 7���`ޑ���BS{u���"�'�c�ג�E5�5gC(�X��@+G���=��q�ɡ@ �C�     ��FԐ��"qk������[,�6�       -��s����<��c	��W�����m)*=[�G�aoMӽ����)%��7j�>{���#wks�}0c=3����X]���d+n+�����79��igE���Fz����$� h�     ZϺ{a� ���*E�e�TeV��-MI�C��}[�u�ZU�d4         ���Z������#C}���^ǭ�\�����bcA�{�P_iE]�M��񩔔�O���4�͞&��"~�Vf���94��퍮��c��,_#� ��>    �`kjLO��'J����gCH��C.����F�{.�f�ٛ7%h         �f_�Hۯ��%eM^O\VM�n�t�߇�f4]|v�v&XTͨer<������lcA&���}i������J����!]����o�F���  �,�    4��}����x��{��;N�����z�YwD         @��*,�搒W(n���Rdz6UT��9�ZR-�m'�~i	��R7[K�ͅ��Ǫ���J�L*�ם�Fщ�h ͹� �&3#272��������J  ���	,�CC�8���	啔�vG�n��{��5oilH/OH������Մ�Zg�IIpb��q�'�����5�u���)=9��XN�/��l           ��T�vȏ;q3�&z�����mU�}9�� �[�N�to ̓` �z::d��K�Ai� @�-ؓ�Z0N̂S�eoM�{v�G����_v�R��O�Z2��M�j<�Bl2��P �#J�KY�������d�+nxt��q%�4j=��w��3�¸*L�݉K��           �aI9��e.d���z҄�0�ێ� �C�    @��.N�ݢ	�ӡC���aoM>4���-�[� �6:�>=HGU�9'�������I���i	�{�?m��`8O_W�f�t��g�$��g�J��3A           ��݅�RUh�lgf"����H�A ���    P��Q��^Va1�;�B�2D��>.v���u4ԧ~���������!��_�=�'�dD<i�Ҋ
Z�f7{�>��h,nr|�:KW�SE��l�߅��@���b���"���KJ�5{����           �q\,�hXWg��щ�ΧsF��B9E%���� ��>    �j�j����X��ȡ)�o�ъvm`(}�2�{zٛ��[S���s���<K_�@e���b3si�l��xp�t�?�A�}=�M	�y���}t#9�           ��ޙ6�tu�
��I��Ĵz?�ۃ��u�o�>]�� h&�     ���X~c�ZOz�ҳ�}gD%;��w��U����O͢	�n	��!cC�~�����<J�
�         ��>]�ϋ"ӳi_h4�-��C,��W��{\d�.<����1b��
q� �|�    T�bc�X>W�㎇߹/:#�~9Dچ[辿�}q����JC�:�@7G�15&+C��#�{Et9>��D%О�(�=         �6�*j#=\��!ޢJ����k�	h�Y��&P��b}�ڎV��p�r0�HEe������ @s �    P�ܨ�2]Z~���%)7�J+*�@W���J��J�=C�/)�o�         @{��`C��{�{���14�^�6���9db�/����ZR����BK��8+:�v@�    �������W\R��8�WTZNƺ�RK�^          �6�ia�������d{��\!������' ut���m+撵�����3A���������}�p����U�~<y� @{ �    ��
Գ       ���Ȁ��m��ȴl�,,��1::�,�n4�ۃ\��D0&&#���F��1h!(qFz����D췌��F����p���Y���O�=��ʑ}��H��D)�ڝ��UtoQV){�
�mۆ�i��p��@�,i������D|�^vl������/OH]l,������p��++	 ��}             �6�j���4��g��d�ߖ�"�ŸџM�.5W��U�h��$��k�Q_�3��#�6y�<q�����Π��p�XnH�N����b�����3����Ԅ^�_,�g�i\������̷���U��v�z=��0��p�k����Z,�g�Qz~ソP;7ksڹr�ƲM���1V�Bʽk'K�������b�+P����qY�4�� ҄`    �]�t���]���\�칆�n�dRqY9       ԇ+�9X��q���B��Ԍ�uV&F���y��`s�}�=�i��h���PrNmy|�u�{<epgGڵr����)*!��G�z��Ɖv��x|��ᾴ��=���h~�Z�ד��U�kS^q)����d�8�J�n��>��֊���X,���8��D�'�{��'撳����_C�\����|����P���5���"�~ ��}     w�h��DC��S�2��ut=9�       �}���\����`Md�E�g��kѢ�2Ľ;m��ᦨvǭ\��O�ST�����Y#�w+3Wlc7[K1����ޚ2�NG�+�3i��݉Kt-)���D��#�D�V���g��7%��
K��8�QPRFa)���@%�*�>Wjz�p��6�	�ER3��}>o�=�>efF�ǲi�ّ���� �*\����ݧ��s�m�����׋��پ�D%:eʭv�zZe�mE�����Ǯ'�Qg���HZ�n���rU�?L���s�j���ї�R�r�.H�}��\:���*oc-�������)6��nkƤ:           hSzu�O�>e�Ao�:E�N_�O�ٙ�<8�`	����>����C���\��hQu���l+���o� �c�|��9ch�l;�T����ܟ�Sai�b='n����a"�3���� Ɇ�d��Ù#�ѡ>"$���S~�?��8���!#C���],s �HI
o���)��bl
�%;~/�&���>���JϏ�/#��W&$s#zm�	\��U���py��q�j��>�¤��2��x�6]
������~}PW'Scіܣ�����h�_���B�P���e�A��=0����*�w*"^�� �ûh�����X������+Nd\���O_��2�fh  @��ʣ+�-�n��      h_�tv�?�����L_W��;g4�d�RHb:��t�"4����DhL:�u������H��Zf�B�{wU��>;X#���.n���lGK������S����HɤO�g������lI������t���^����j�8�Գ3�\�r�KISq5®��>^g�ڪ�w�*�����H��p���wpQ]i�_�ޛtT{�$�DMli��kʚd�ۗd[���l6�h��M�{Q�)�{��{��3H`�3���0w�s83Ý{���c��u�X��hIO��a2�;+�(��bc�V�2� �S���ݖUX,��ˏGҡ�dhm\�v��۩����~gT���F�+�v6����*붵���R��F��xm���� ڈ�����i���������l ����+��K�Ey-^W~Q;y�d���N��xe�y�D�O%����ܩo��x]������{~[��mG�       �%D���S����|�~31;�ܜ���DE�����1ɢ2�>�y�>�u\�t�w�NA�q+���B��墳���:����y�c����Y}*J��@�u��e�tC}���H|
9*s9"�G[��@���|���5��;M�����/��[g �Ú�?Mg��i�����:����66��$�-~��Q�
���v�/��K���s����R���������}��c�$�ӷ�Rg���/�n|iU��?77W��������M\Z�l��!���\��'҃+�Љ�Y  �FC��x��s�TT�����Szz
����CYi̫�{Foqƛ_dFWIv�?̋N�����7=#�        �a��)��
ϥ�,���JQJ�!��O.���}DЏ�������z�Ҳh�7�Ek�!ݼD���~���L���)�u�\��;����CAI�[[Rw7'��U}R����~;@�:.���-�?�/�4}9+�rxc�c�h��kD5FS�Q]�����I.ˡM���Os�����
!����-Mn/	��8T���)4p��ַ��%*B�hj���� �j��7���v�`��Z���tvv��sr�7�ơ���2jM<^'��m+��L�} ���ʒ��;�&~��  �ƌ�����Ԭp��Rӓ�������3�Y��b���S�xe�f        䯽���p�P���C��8J��uy:�Q������RZQA�l;L+�M|?9��t�>s����_D��L�/�70p���\�+� kr��"�p{`;+Kq������cz?��W�N� ���m�9���yt�W�)��iHw�����9l�h��寴v�\�Nz΀����?n�g�q��g�4��l,�>$�;�&>��Ѣ�q�u��>%��q)�B����bn�5f�**_�R�S�h��b9 h?m����T}�E{��x���S�aF�p���ފ ����l�ɑ���}  ީ֜p����T���hDeB/o���掷�c�ɍW==\��a���C�%       t|j�>�]�+*��eto�������^�"�Żf��z�l2��W�dW~�b�����R�}��jW���G�]������*�ᾙ4�Ww���H��C��.��ߊX6���E*t+L5&25�f|���?r����aȥ̢{��H�sS�)k��p9�z�1?�ts���Oy������>�.^���]�[</�R����=0���p��U'�D���y��i��Ƕ���yq1m�Sq����eg��k��Ƌp�i@��M
�F� �#�}a�q�\وl�����RJMO2�P�J���x�Ye�ee������:�xM|~��I����U�t_y�"      @�V8�VP$���%1�zK�،��r�/��X����l��
�W�'bkia�nE�����РL����׫�t%��ֺ���绍��{o�[���ف6>z�h�{15�LAbM�`���_��s�'�r�Q�q���}�n;B �s�T^YI�h��Y����cĥ��;�;�-�K����HOMBONBc�h��K ���Bn*GG'q"BNNۄ��{����>�v�f/߇o  ��/_W�����i�%&�Ҙk��ǅ��/��v�����o[�P�� �[08Tێ      ��B<]iz���N�����Κ\�l�BcF�U��)�v�X�R2h��X�>�V�k(��[\���gH.-�@���kM�ۥ�Gg:�r��冼���]�5q]|���s���$s�ܰ��%�r������4w@Oўv�#��p߅��Hv��[?�suL�?�mB����|�+�d.uq�)��)�ݙd�_r����W��J��5�d��W���!n���֖TP�6� e��_ٰ���-�f(�އ���.���'.*~��@q����LI{��TNNN�kk��d/���Ra[��i�hG�3  0y=ܝ�Ρ��a��Y�����O]��|      ��.��_0�8m��qopYn�կ�V��HΠ7����������0�����֩�z�[�x��v*1M{}L�_����k�U�� �`��*_h�õ�S�_>�cH�ಊJ��C~|b(�w㣷Ӝ�ג�v\�׆P�֧I�>�-�o�|�[<�z{�����"R2��9P�������v!ٝNJ�>~>�yw�#����tcD��pxo΀���a7�]��9��I���Ϗ��ꡌ8���`��Ej���d	��8���Z�-����6��mwuv� @��;N4������ ����ԧ�?���ծ.>SswT-?I�E�Pi��     0���'XqX���B
JJ���\�����M�m��=7�6�������%�}�yK���$�Ԛִ\����Z��q�_�[�6�Q�޷�jwm�N+ϱA����3-Z߬�A����I6j�L�G��ۭ� cm�U���m��T�;<���mE%��6��̸���tѦujhw���J�қv�?-�P��]�x.���t���5��y@M���;����!��u���2��C���T�+Rևߗ��wJ\F��=�k�+nrP��{2�t����z2��?M	:Le�'|�hȬ��@������wɒ-ԧrttD/	!�  �� �Tj˅{�����kw���������c8�     `$X�ӿ'��@�^nden^��Jˤ��cE��s:U�dei�A��]���q��ݗ���+i"`��S BSj��\cF�����$B'{v���-a����Ь/~�I���bj��z?_�z�i�>^n��80��qZ^�!��V\VN�.�&���b4�&� �g+��j��9�pU{}Z� ��}���=�r�8������Ά>�7�dǡa|�>�G�����m�:��h��޴�Os���dÙ���t�/��_�:;t�n��Q]񵥯a>�Ԫ�ԑ�K�gW����O�����'���\�z�i �q���L��)VV�F]�U����� �'�     ��_��[��pw���|6&�`�ZSU�ĕ4��      ��+���ֱ4S�rWc8ĕ�����a��ޫ�Q�d�st=9i�6���^۸_��R���~7�	��f��c��У�ҧ�O��ִc��Z\un�2��c�RIF+O^4�z̕q�����zai�Amn�o���YY�p�g{N�j|��!=�f7��W�c�i�Vf�8&*������	�5g�Fێ7Q���$U�;z���g��*�3�N-�z�/�.4oP�hO�{e�_\jp��� ��3ɪ��&B�    �n��g^r>�ڼV�nށ��\�h��=2���v��      ��&��J���r���BFQY9��P^I��p�gk��`+Z���[��Pս��&e;O�� ���V��?[٬���{���d���B���$֋`_����M��s����l�y�B�W>,�s٘���n0RF�9��29�����RhS�\��~��<)��'�qظ����qC�K���}�I4�����foӢu�*��s�^#�_R��c��������-��UoSB�m���  �	�>    ����Oc��=���J�g���@L-;~�֝�,v@     ��uss���\�-W��H;.�Ӊ+���]}8���&�t'ky:ډ6�K�Ic��Y��P�]��ߥ��ϧ{N�����������jX~ʺ��嬆��q�9�W�2ʺ8�ǧ�B���Sj�h;ܺ�+�1n��\on9$�fsH����ߦ�hq1���AP�8\��B��   �}     5�@�ӻ���:E��g�B۳27��wot9n�YP$Z#s��e׹�g��=����e�����P���y4��m��(z�����҂�����-���\��e[���"?�7����)�>�u���V��.��09�
�n8M�~��     d��ͣ��>>��U;)��m���s�Ψqyk�!��m���Q���֚^�y�������A{�Pl�Q֩�_g{�: ��w�g+�3�ϵ~���E��z!N\���mGĥ��y~��Lu~���i��'��ِ����M3y�"���N'����  h+�    �!:#��\��÷��H�2_���m���Yc��]��_ۏ���1I�`����Ft����<���kl��h��U3���6��£��P���nr��C��C}     2�����}��V��*N��JV��-{�Y����uѭ��)e��[hʢ���	n�k������h*���L��>!�È �l�T�&�!�վ��)�s~��-�x�従��v�*�+^���}�Lb~��G��;�PO����kO_�/�����b   cA� :މUTVA�A��@s��V���c��9+�dg���++1l�N�f���y��Q�9�e�jZs����v8.���_ڈ��9�0m8�󠻿�(�b��k6����c|�0�Ӎ.�f6z�1�~z߇�����&B��z�Pw�C     �����������t��i�9��D���ڒ��9���V�s�ק�v��F��79���zJ�
A۰S^�o�C7��A����b2���.~xa�zb�`�^�e쬪�w�2��c~;[��=�w��M6���`zv�0zd� zq�^���y2zv�Y�H|
�O�֤�s����2���U� ��!� �F^q�� @��2J��4��-O1u���ʊ�t%�
��Դb�,��6�lW���S�kxG6)i%��W̯i��)V��$}�z��
l|���#���Y���HZ~,R����U�f~���m<_^���E�'�!ݮW��
�L����JV%d�R77'��� ���:��W�� ��n����A׃})9��(�e�v6������uuu�q�Տ�϶�U����!    ��<l��c�5?X�+�Z��ze�?W���)��?o���?O$N8:����}}��K3F���h؎���YPl��W��=��j��ǒ��
�޿,��6����m�I��ϱ�.�*B�*��dњ�kkeI���!�~�=O-��۸��?����ҍ>�7Y�?�u���`����˯_���5}~�����)��[%w!�G���fO���Ҋ
��S@9�%d��ǡ?og{�2�~¯����:��� }+m�1.{`�x���ȉ-o�:�d��}#fР���1��t,�* @�B�   �p���0W�f��*��Ǖ�L3�ǡ���\��������wL�b؍C}e�9d�*�oS�J?G�?(��O�#���z�(zy�H:���@�NFQ~	B�2��I|��+,�?{�>�c2�aD���K&�?ruB�\-O���]=��E����Sq����1�o�o�i���G��~����c�����ҫ�������sho����p�C�    ��]T��������)<o'���/,!�pe���Na�����s�l�*&q��OJ�
I6j�����gZ� 1'�e�Q�P:�X��g���F�����&�p��ȫר����|p�$��?����!N�k��o3Ǌߙ��Ͼ�o?*d������4�ϯ�M�9�B����� ?֏�M���2�|�dc8��[�ѽ������mGh�Q���M�N��G�/7���r�(�Ә���ڽ$���)z�_ޯ6�OZ�b�����[�����a~e�f7��7��q������:y�N%�QI���7����[�+��0qR8{i�H:��F�\���ȋӇ�P㪪��(��'9?�t3z��4��3S�ҝ��H  к�   ����T��kj�O��KLny�����P_5u�Uʵ$oK$e��G��ӧ{N��n����a��+�F���[��ӆ�Ѩ�'>���_w�e�B���m�u�2��uZD�N�7�;�+�7���yC�{k��b�)�Gyn�N1���;:�yp7om�?�a;C�N��D��Ά�+�7FD7x~,����c�IC    @v\����Zh4"4�۹hji�$>i�q� !���Z��U��{��^�Ÿ?H\.�g���񙹔�[ ?�w��"+y:�S7WG�ՋB=����v.�~<r��}���}O�Ioo=,�14�2?7����(��l��2Q1�����\c&��~�zG�'�O�[���P<2���\J=�|;�NJ#Yk~��l��h�2�/�)N�����{G���������E�e�IJ'Y�޹��뗫�u��忙�.�"���t�w�"��a1��Ý��;��}v�.�T8��塞@��.��0�}��b�����빚#��<M�����  ��   @H�(mf�O��K�'�57ԧ���'�?���T<^�_3�5����/.�Z0��;���t?�
o�����ف�������g���u��KԻϘ@��}�S�y|��/\��wtr��^^�t��z�ۆ���>����x$�0m����a���V����Y\窒<n�    �pž��	-x��I���}T�Hu������h��x�y��U]����m�Gu?c{��KSq�!>٩J�lA�RU3\A�chF���/ۛT�����I��'nqŤ�㴩6���J��O_,�F!��b�	��&e���?W��[M�:5����|�Izs�!��շc����Ub~��_~lol
�M�b~���m��jfU~�UU���s�Aq]V�������5�����������b�A����W��e#|������'m��je|�,e�;��@�ϥq���}8Wz�r!�d�'�s%F����-^�Y�`og��$  h=�   �����}���.��Q%�����l�M�P!�
��r���g]�0���;v��+_�-Ţ�������r�Ν@OL,ڧ.=r�(�:�y�%g�}��;]\��wܩgL�N8�R��t���״�=�|�`�ܿ�`���:��܄�ˎ]��;J��Se,�E�.��>����\���2    0on9$*Aq�7����p~T>_q��tbz�a�2�'c��{��i�q|�n>D��v�y�8��'�p�q݊ߍ��.������t$>����~o'{z����J���t�������Vnw�s!W����t15�dv,�*���gQݍ�C����Õ�տ8�[{|\�����D�,���̯O'�_~��>XF/N���Q�/?/�uq���c�O]�]�_�����~�u�U6M���t�ZlJ�O��B�Z����p��=q[�`ߐn^�+�$�'�����}��7n`W/�  Z�}   @e����J�EiYY�oi�߶y��8C��-�hV� Ѫ���hjNO�����+i��D�hQPԌ
�|%��Y[�����rH���%�Į���`��h5�w�u�������N�a:m|�`���:���$Q��n�B_��o�[[�������@     ��Tb=�z7}p�$���~0�W�涴�y��-��A��p�#g{������U�L"l���)n��U�{y�Q��+��ۈj;vVT�|�/()���q2Fݧ|F�	=r���G�����8�j�t��硭�usX�8�u2 Wq{�V�3����v�mM��M���jVj��?���..z��>�����7S�������:~��_�9��ˁ��L�n���Jn�2�����������1�\}��S}��%^��3>6"�W|�m��:x4�+0@�zuP�t����5ʶ�u�}��S;�  @�A�    ��x����gZ88���Wo�Ơ����ҕ�����T�
n�p�쳶���|c�\>08��`�mΕ5��c��D��������y����nSq@otM��;���7�7�O�c�5�@     S���J�ɣ��L� � �}㠟_����p��5{hgT�>��B���i;�r��|�=>~�r�(q�ֈ ����7����'W�Ⰴ�p\
-Y����L�# ���O�N�/�P��T1�OK�+lr�T����P����ch��Ӏ���������;���N�����T_���L���|\���W���{9ډ�dq�n�ǥV8t��&  h]�    AJN�8���Q�a��CE�h�CU��:v�֮�7&Я�`�lj�yW��(!3W\�3�O^Ig���Pw�:�6���пkn����	�95�ϓz{���[����c��tN�    ����v�����>�oM�&���UX,�|�m��&UA:�����_�Y��EӨ������������	����s����v����t�'��s�������|��;�����T��ru�/�{~?��詽OG�_����%��R�a���t�_�!����=�V���M�߯;��r�>S|��kT�r<�j��Ǖ�U!^n���9̬-��X�����Qe ��!�    `D���['�嵍����!�hho2�]x�gbϮzDخ:�j�dd�P&W\d�x*��ã����V[mp;޺�}c��?-���Қ��3��T����S���1]\-rT�����ˎG    �)�v�kO_��h'Z��W���ճK+*D{ڌ�"���EWs��e8�.�n5�����#iɄ����(����%���;�U��)��l2uSB��'�'�U�䊔|��~W>4�~8A��a�^{mS�U�;��r����O!ߚ�*L�_e~����P��i?�u��������g~��ӊ����rº^���r����hZ��l{��\JN˷Ru�;�l�`�v1�v�'c�t��Yw1 @�B�    ���i�y�33�6�dcE��G/N�=�q���� ��D����C���\5@�n0o�j{�<T\�O_�;��s�����=Y{��`W���o�z�G��G�\�vGjeA    ���O�I��NKqŧ��c��N�l����t�W�	��U���NG�R��g�}v埽�a?���i���Ο��6k,�7���s*�'��V��?�d��x��{�ӿ���Ő)3d~�9p�䫸�5�9E%��2�������tsX��2��w����K��ו���;�������w̔����J{=������羊w�I��_��9Qw�����\��;����< �օ`    @�B�>�	��Bk�ջ�w�z8�ROOW��h�~�g���vO����z���6��[��T��y���;s9\�gj���Ew� /������ކW�����v��I!�h{d����w�]�C�      �O�O��I�������ߢuq����'&��,l��������BA�?����U'/Rf��VA��U�jU��q1�����j�N�-��\E�?����,Q��~�<~��u����J�xb���rH���/�j�`Y��=���~�B���_�����zD���mu��`mI���@/L.�s���n����4�e{/'  �.�   LX��|[CU�N�
s��vks�Ҽsl�Uh:�8�x��Pn�k��lz���E�������ⶻ��>�`�������<�9��N�=�c���A��Ҵ?S��o�M��������"��A�m/     \7�����J2� š��Ր��{sp�ӏ�O�~. �����;s'hO.c�Bz��+t��Q���ޓ�3Ʈ��ڸ��_g��T����tr���'=ru���Z�w��@?����)��Vq��}k�8��O�Μ	�pH�����M�:#����X��������	V'l������E:�k
�_M+�V�Hض��H�s����h#������	���/YTVN��� hm8�
  `�)�+�<S;pxC� 4J\��@ιW�9;�:�J�9E�#��%��l�*)�����F���.\�F?>G�+��Ҳ����MWs���L���^'�����P9��>66�O?ا�>މv1��Ĳc������a�b��h�6��ug.7:n     Y}�h�c�!J4R{7�� ����$���|�t���y�EKC���Cp㟷�����j������~�@<�<��gO��.u�:r�>[0ET��e�?x��~���ݢ���$��ߦ7>����ʝ�j���;�s銨r�noK^��ۜ.?I/��K�Pݭ�����9�l�T�5����I+���Qm����@��le~/�*B`�)���8�:��G/�K���1���wL�%U[�1q�պ�W�^g*��ߏ_��o���*���=���6��U_����_��&0�]YE%}���y�8������C��������̯]���7�v��:���*e[��nk�l�5�  ��$�~�k��)��{��<�.ڛb�FR���s�:�]�3����w V��.��J�#�w�p����������4��l�	�۸nnq	������&�4�I�;����|��ܜJ+*������z���$�c�������='�un<���6� li[�k9t06I�������Bh��(��_�v��Gц    L�Đn4{@Ozg�a�d�	Q�����G5-A�4����k��r��y�^����O��[�]|��Ǖ�ߨU��0�o
כ�]Q	�z��g�ի^ǟ��]�[���a>��P=^ݰ�~8a�g�5�/����|�%,P��U��b���m��	rV�4t~w_�B�Ly~}ݵ�/>����{E�P�����/�Ǳ����ɡ����m��W�HF͙��F��V��OϬ�%���tћ�W����3��<���E_u~��Ĥ�������ɼNv�=p��0"�zy�Q���?s��:�G�����ʆ���yjhwzw�D���,nK�+��w' c������b*)�3�A7;;;2oQQ�����T����	�!�_   hT����S���p�ڡ>��4܇P�DjnA�[S��N���҂u���q)7�£���M+xG�7ט��� r���F<�mxuqˌ�5��;��"�ajw"�g��    �)��rSL��UT���մP����5{��= �mt�����i��b�4
�⢭�7�oP���j�X\^Aoo9D��9!�X;��k�D��P�[�6�q�������)�:Ws�����_ �J�2��;����]��(~o\͵����n�R��_�L�D�ߝ5�Ԍ���ɢo7�0��&]��W]Uy~�T氮*�uͯ�������~S��o]�;��7���@y��W�]����m����_�9]lKl����W�RBf�8q��!x;�Oy��E�{P��m���\��|����GIII҅�8ԗ��g�`W�������D��}TXX�`�dp$  ���P�B}���/ԧ�y��Z�(�A�䲿V`ol�����xttFv���*�b����8 �-jN\I�����h��֞�L�Ι Z`��%/���?=�⪀     �������)��	3\���3w��mܯ�nX�/��zݖ�����%�l'��c������1�x� q�W�;��=z���j	y4�*�y�v�sI&�f����Y�=��}~�Zy�b���/�ܚ�������_Ϯ�E�$���WRF�u�x���3)���(��OL-�et[����=����˭K�0��-.�'W�lR�����{����x��/�~�o��{����_�G6z_���<�s'ҼA���ܚ�b��QC����m�:����,��vV	��t뗿��s�+�1_>4�=D�Z�Z�Y�1��q�O����k-����P�GS  :��3 ԧ���B}��:H��>�UTZ��1�Ys�oL��������M�>6V�?�t��;�/\�f�Ǜ_R*ڸ,�[�S�`���_8�      �����b��E�)�ӕk��-ҋ�e;��s�M]-���[�L�"��vm���V|R��q����L�b<��o>H_�;E��'>K����˯���Vn��O�i��hz�����W����П~�bP��-m��6���J�o։���$���|>V���:�)󻡎�]�l�A��ďӘ�����YK��G%e$��/�zx)��ee~'���<�}��K6�#�?�w(����~T����MBV^�,�;)XQiY4�_�#����{YC�]��S�ĉMy- 4�,a7nG[P�O�M��"�'7qDu���]lmm��De{��I'�WRUQ�o0f����F��%4�Ñ����M���3J).������<L:�ׄP�ʔ�}����˛x��>��/�A�Ft�!Ks�^Ž���q0&Y�f��|�I���WY�K�q;^����Hq�r    ��q����L/�IK&��F���g�w��Ov��۾��%&W���/��Rz���4⽟�o��j������[�b�8Hr�-.ի��>	W>�}8o2��$ns���΀_�-�ݵ6c��wLU��y;���8K�2��r�E�ߤ?������A9��/��i_^�����(�*���M�vd�шex�2
��TbT~W�NE�� m���nm�S��xꓟ8�jkk;����;0�>����u�i�����=Z���s�t�3R7�g�/q8��L2�׌P�J��. ��T2M�i�g��>�������-iHW/�`^#�����K���;�^�Yk�6�*5�PS��q�    ��(.��76��jg_,�FA]\���BT�ѧ����լ��!�=�ޯ�J_���P�����yҠ��z?[�l�?��ߔ��ѝMN����h��F��Et�w���]��O����/���W�2��M�i����{�W�wH/zg��ld�߳�F�߅�_�W�z�iqQq��\���b�&���
��u�O�^㭪�D����*  @eR���T1=G�L����>��M,܇P��}��w����q��ƪ|����k9�-���=��_W���}�sm�g+�Zfp�    ���+Ӎ�p�m�XQ%�̌D���YDe��jg�]v��DZ�rG��d=�Wwт���Ʈ/����W6쓲�%p�+����@��KW�׹sW�
R�LF;/&п�O�LZe~�G��=�ߥs����>������B�t��Υ~����N8��"㤮���� Y�uح���]B}*oRR����ɿǡ����/GW  :0��!ԧ2�p_KC}���H��>0%S�QF~��u��"�q5?C�R�v�=j*�ݦS1$���Uv
s�    �3���3�wц��鳅S���Q�P�**+��E�)r����g���T\U�[BN�.*�s��[���?��ѩ[
ʪ��;�� ��8qQt�1^���%+5Ч����@�i���S:����/u~9�%�^��ބ�m���˭� ����}���o�������$܇P�i�V  �N�p�C}*��}�
�i�'y���."�&����M��4|�������&�]�z�p��1I�Y     -gomE���7����9p�䷻�����M&��l<�'W�a�����9g.���O$w{[
��B����?��}���)�F�Cq)>�Wn��VL�ʣҊ���@ߋ�GД��$���&�� 1��B����yh��0����}A���&0��e�l� �o������Ӂ�d�VPD���2��>b�|�_|"�l Ж8�v��e**j�ך��e�U�3���/]�t���[�fee���cS���   ����V��d�U9ԧR�}��n#�Ry*wq�/��t*G�LLxt�^�>�~�vC�μ��G�    ��ۻs'�C������Muվ���ipW/Z�b;�t�L���5�u�Q�O�STB�o
��E�-���%q`��;&�̾A��}��6�{Lp�б�	���с~di��q��LR:���(m���[>��E<������Fy�o>K �q�����__��T�oE�:�G�s1zˇx����9,P�v����Q�ݤ26ȟ��6\��W_��oOe~g��[�_~�n��"cs�9��{z9�����\~���~����Q���o�2�<��c��k� 73ec7''G��ZCHHYX��,��r��5������<���H+  @'!U��C}*��}�l�P���}���I�C�Lپ:*�q{ދi��?&#��������}�e�     ����}4o��v6�۞Y��u��O�O:���s�ϞZ��d8��?��5w���s2���E]��
���6��oϞ@N6V��͉��i.���D�>h&^��U��U��?��������C�c�5lky}?Rye%�:E�+�\J�"������O�Z�K�3�~�������wT��!��������<qQ,s9=�@���������_�M~7<r��r��1,��)��]��ICD8�.���{X��ۅf~���KZ�]hsqu_]�xG���.\��O)�}����3�z����w�  	��  t"�+�wk���y�^Th������<2�HS޾.�����ʎZ���H�Q���������`T�C���~�A���;�t�-��kJ7���n&��|DJ���?������_%c�3��j&)���    �[zo�D�3���6�>f�.Zw������4�_K�����#{��_~�E�ת,$#�P_nq)��q�U�������b�Vp ����O3z�0��`�8���'�����h�x��箺8����x$}���^�!�K?zw�Djdz�՛Fі�4����$���J_<��r���!��66��(��-��hhw/���:��<Nq��~��lhT�����b|��>n1̕�tq�-);_�P`ge)n��I��4�^Z��d�U�y��m��k0�7R����߿_�1�^^���xx{��ƚJ����Q\Vn����������(%��
Kq��)�W  �N&�Տ:��.�Yp�/�3� :n��7L��
�nYu>ݵ�xw\Dk    0���[[�m�U�㖵|;����W��˲f�mk�e��x����;));�I���ǝ��@���K��u�8h��?Q~���� ��ӓ��UMk7�����h]Z^A=���C����A�"`��m�hhwom(���ϭ�#*ნ��2Lۚ���me~�&���۟�
s����4<�G;��n��5��|uf�L��_־��v~�������5{�~}~��̯�r�����^y"��e_�i�v��zZ٦�E��̕
�L$�ʼ̃���;��B���N�J{lE�˕�^�K�G��K�GV�WyN��������՛�z�M}i��7���F�3n{|.%�V��(N��+nZ����{�ʚ�B���N�Y~��Wֽ3*���w�$�`           H�?w��յ�"z~���TT���r!��}�3}8o2��$n� �~r�Nڪ�\Fy%���C���&U���ヾ|���SE{A��ā�[j^w6���
Jש���WH�b�)-���0H��d|��k����ȋ!\�%��+�R�7�x~9������46��=����ջ�ۃg	���{sX���"�w�^�����_H���7����Ӛ�~�+����i}������O�:���׃q\M�ۊ���ң��E�=r�B��7p�ݕ���K���*�*�ێ����<���*���0��f��%�[%�Ø<w|�Ә��O��H|�A��uv���N���t���с~����X  y!�           ��=��)"ZT��vd�� �=�m��Cz�;s&��>����D�����f�g+�-���K��^C��ж&h���Eȃ}���^�O�;��Cc�k��o��/̧����g{N��t���=8���r�?7B����q�>��뷾�I\��Q���r(��B}���N|M��m��爛ݴ�����"�_��v�+bq�Zق}����i��WuS�y��x�\��}����:�E��y�Z�n+�W���TJ�-P~��ݛ��
�g�ļv����t8��p��6>z�����++it��*N&��̼�� ?� @~�          �T�����E���
3���y��U�f�	�gV�t��Sq�/���5�/���9����h���Y���$���3I��.�[\Jq����]��j�>�q)"T#���餴z�������ÕJ�+�������ߐ�?��������o�g��rOS��&��[��r�}��ם�\oU]�hȡ��..�"�.����x{\��F�����c��ה$e�p�G�չ=ȡ��%�)�YY������~a��pp�����r,�*=�|E�eݰ��̌F*s��� ��}            ���cE��h��w}���Fo�6�:���u}��T�`�����:W�lHBV��%g�S^q)�:c�/�6�-��ds}~�(���9���(��[���{~~���9ؗd���jg#�V��R�歽έ���g�s��"�p�bV��x�_��ƛ�/�cN5놦{�Qzty�2/U�.�-r����?s�����B��띟�cҠ������t����z_�|"ȁ�$ �!�           �xj�N������p��t�^�>�:�.u��ޢ�!@[�*A�Ҋ��#\��]+(&0��-�hpY������ḫ�o���k����r���ű�e<l���E�gQCr��[ܪm�eRd�xݯ��rzv��T[�Z�k�碁}����R"M��]|?�ϣ�`�^2a���ۿKV젎� �           @"]]�\����2Qu���أ˷QG��LOM"�r5%��p�J�6�a\	�a���'�^�Oj^uE[n!��M�������w��t��U]m�� �JX�4�f[��š���/?G�Us�k�T9��]rJhw�9]�V�P\2�J��m: ��     @j�����!��dO     о��Jh��h:�p����mK��nɻ������VN9��~/�M&�0�������v(��S�}Eu��C�C7,s[�`����Ҳ ��jw��"o����ab�������o� �uC��E��vD=��<UZ='����^��\���,�5�`mE��%�� 9!�     ��k�/�&v>     ���8���z���v���u�T>������hmE�����M+�_�#�)7,��_�i�W>;�Rd'��@{xht?�-���YpM ���NRí�QyH���`{G5����`���J�3I�r�����@65����Lu~?C%���^�e4OH����� ����`ߚӗ\�������H۫����)�[=�7f*�r�"�3�?��	2�9��x��9I=ގ��_�����4�mH����b�Տ�F!�n��n���N��\����F�^ !�}����*-/�rM�<àgV  @�noK͛�P    �d8?�������X���|�;}��x�@��ϣI!��Q�����u{���z����3ǐ�����[/��{ۏ��� ����CZ��ő�P�Íya��$���a-�o��敔�}�xf�q�7��L����/U��4f�h)�����b��P���hëV�����h�[���e|��6�?9'B�<ޝO.�a�����s�J�뻥O��Sxonu�w�(��O�o�[��_Ee%�zr��q�[�������<8����F:��9���������� ���K� _�J�Rr��  Ӹ`���$     ���' �>#yz�0zd��zο��cPbv}��}x�d�d_��9�����"�  4쯿����"��-jo�	��8H�⺽��.]0$T|-�����rV�}c��G����=����ZR^�m�V6g@OQə����ջ����q���^�b�4���Je���T��J�����CTy���UU�=2�&~���� ��x           ډ��=?m���+Yy���%J��#;�س+���+~�d�`�ZM7�Ǖ�^ݰ�Υd@{9�}��x�����w>��������֜_Y����ѭ_��OLѫ����Ϯ��h��	���ݼ�u��������ق�u�����skv����*�z��;/�Sa��������j+9s����/yk+����*,���^{��P~��[<���:���5}<o2��z���     )�(v�j    �|�ZȖ�q-7oP��-���7Qqy���oo=,ڥ}p�$|e�(q;��\��V��"���a�:.� `�qq��t'l�y������F���.B�^��X�pv9=K�=�)*it\��M�����D�� ^��Q�oB3���+�x�^�{��,̧���9����:N�<[��]^VY!�1�^^����혌lz�ʹ���E ���<	-y�`     H�w�=�j'}�pY�k     ����zmx�dd���Z\VN���M/ԧ⃹7�Ҵ^��AXn��UX�ħ   4_��k����Ǌ�)����B'��	�r���璛�����g������aeW��j}�N^�wY�~<�Dc����S��K� �`     Hkŉ���������=    @��.*��g��X��V��,4�"�X*��(���d��*��T>�p5��l�'�}���I����rdm�͗UP����2u_�h5
 m$���h���`+�_v�=�f�8��1���Z��/����0��zy� ��>     �ZTZ�h=     �W���b��/1;����$g[+�56#����r�������Pըc㶕|��i�2�[1� І��9цG�jOn_u2���b�81�������~�����S�
��]mm �`           @;�4�n��S\��r\�E��[@    `��\i�#���lݙ��Ȳ�TQiX��q;���uK�F�����^/*+' ��}            &�)z   @N\�o�#s�����~SD4=�t3�WVRSl���''׃=\]>��]{��Z���           �l��6���Vf     ������-�KA]\������?n���������$J�+$/G;
�t�P/7���Y��V4�o�����	 �`           H�+�趟��l�(�ݹޟ�8��]ohYV^Q�
,    r��P��"��v\���~��J+*��>�������Μ	dfF���o��䟽�����Z|���K�#�Hv����*붳����>s�����x����            �������!�{�M�.�j���   �\>_8��Դ�����E"�ט3I�����u��o_4�7��I{v�UϦ��~�N&��#̧=?u8��?X,�Ŭ�_��Y�R^^������PNN� ??�ƛ��7��4 �     zv/t&My�������pڒq�**+�?�7��܊����ҁڃF��^�;�?��7>��r+����           Z�������̌�e��6���7���E߮�M�ͣ`�г��p��/:�ɹ2�k����2�[YY��wr������>1��x��JyNp��`     ��4G�믬��J�ÿ6��7�2�.�;$�ܩ����i����     ���d�Qa���%��    t�y�4��e��M#�a}D�]�O���I�-{w_J�n>D'����8�WZZ�f���̔�Svv�T�k�P��ٹ:̈p���     ��]���(r�*�Jss*Qn� ���m�L!v^doaM      P�)��B    �y��le���Oyy�>zc�і��ف��5��WH��(���d�֡>�������ᾶ�LX�}��>    �66�����~��r"E�e���H�O��B���^|_EfTa��J�9���Z�)����m           жJ+*�p\
���
��8�Ǎ�rr�&����E�O~�    ��[��)ô�/Y�ä�}̬���u�"��
�
�B�TV�O�daiC2����WE            �������+��v�O��"�'7�     ����2Ң��JCs+��s%Gw�h4���
rc	     �7��d�|~(*m�vT     ��d	��Z;�'�x��}     `Ts�8{SEy���QYQ
�姒��/�;���c*ȉ���p     �]��#     �


�
��8�gff�uVUUI�Sq���4���     �2#Y�vQ>�V ,/ͧ��t*�O&3�9��9��c*.L�i�           2��[Y������mD�X���Q�-�`     4���3Yڸ��ƒ4+Ҙ�WK�z���\oY+q�X�PAnYZX���          @��قdU�A �     M��H�M����UU�Svf<�{�FcN             p#�     ���:�See,]K�&w� ��             �`     4YsKś����S UU^���K���I��dV�wp�             tf�    @�23Ӑ�K0ir� �
U��������i���}vvv            �� �     m��}��=��:��s�[*��ы��D?+�\ii)            t6�    @�1�r kW��s%+�kʕӜ�#߮D�            �3B�     �L�]nK��[�K�q����,�˨�����8�            0E�    �,��H�� sM%搽�            tF�    �$��ͳ/�e�QvFYZ�Rn�G            �|p�     �anaM�n�TQA�����=�ll            �3A�     �������m�1'W��D���EN�����    @�f����n^49�;�z�Q{[r�����*�*,���<:��J��)25������%M��;���ő<l�m�E��WHg�3h��X:����u{;����7�~�J*%d�6y}�8�l��n��[@�b���-a�dea�w��@LR������{���"b��������/�̕�d9E%�+*�����`rS�_���ٻ�6���?I�{��މ3�	$� a�U�
��-��P
t���.�-�B[F��a��Cv���޲���s$d��Z����Нtz�;�9�������z��vƈu�3�g��<�j��ŏwΨ��v�>�<���׋q8t��A���~�1����=j���t�q^�X�m������t _�a���O^Mm�q���J��Q0|�}���X��q1:ճ�^;�
�bׁV�i��3=�hλ��e'%��9r�Ku�s�/����n��5�O�d�ֹ���W�@���x��2�[*��   �}    ��|��t:�Ŧ���l[�ּ����Y�	   @ג��M�O��&׽l��҄��t��,�`�xZ"�3���8N�?Jq��o�f��;Κ����o|�7�nm�'�>��]�^ߝ�ZÄ�^��kV̟	)�~ln���ۥ���*��s��Z(���ӭ�W}��������3]��	@�x_�}������{���	��}��������Ԓ/Z�x�\v�4����O_Y��zI�c���LH�V��bct�I��zj��f}�9֗��g�/.���cݫ_F����y����^������l������4�[����������z�&�ٗ��u��[<�9�~u�4�<�o���Rm ���0��m�����?���2�+��ooa����oUTר%Lx����[��Ǵ�`   � �    ���gWR�PE�Ta�N�޾\Y=r���    �L���.=ݪ�������8F7>����;�����y�Ӕ�L�ʟ�V��5�h�����SoY����k��/��*�Zj���G���*%.Ƴ��Z|���IV����gL֋�7�8|
��⃳O���	8��;����9�j���j�+&���3F��1���jO��E�ݦߜw�n�6�mk�Y�,��?m� �����������{y΋kO��,   �^�    D�؄,e�$��h�宗#*Qݲ+:�
Ng��ˊT�TMM�䮑ۚ\r�j�h�    "õSG��N��:^�;;����vi��|.���Մid�h��A��U51P:mX�&�}��ֽ�R�qLH�5[�Ά�V�ߒJ���tl�n:��:�tM��/�E�|E�mh�i�Jm_;v��_�����j��� ך`�e���g�i���F�oV(|g���k���OSEn���VpԴw=\Zn�z�y���T�u�@�7�o�Nڷ��>3�>���<B�^n8�g�/��jrlӶ���_�h6mn�i�۔�v�c��(�U�k�s�������MVu�=%�~6����oz��y�b�uOIԏ_^��
�^�Θ�����   4�`   ���JPJ�0�%䫴x�r������ԞJHJ���H��e��(�|R�%w�M4�   :�ӿ=������O�V����k�@�m�N�c�6[��T�{��u�3�_�����׹~cn�nݭ���j?{��~}�jA��ًמ��|A���gBR�{dZ�f�[�߷��~�}���R�LUkm�lSNv���N�O=R��Z�
�`��vt�͘��|�E��WWO>�jo�ϴS6���&Bz��������c��ZZ����!}�V�^&�:�g���q�t��\j�X���7�۴@�t׵�e�&�<�`������
��z�S���ժq���#o{��o�-�-��׏N��Gmn*6��_���M��T]������   ڃ`   �#&.]ѱiJL)Te��mSa��?ϻ�+d}�ɭk[    �랡������R�f^�B6_�;�o?=O�`���zf��*����?���Ea�w7�Й��7n����;�j���?TK� �gM�*�M�Ǫ$g*6�?T���/54;Mm�+�ت�f�<�K'�_>X������jEl���+��� طt�~M��Ú7��M�߿�Y؞��>��uC}����9��{P�<���|���j��&���o>�o�Y�w�,k9=!�j����(f�f�c�J+���_�jѶ�Mޯ���j��~����YV�>���p�}�ig��������c��OV�`��0   ��    t(6�M1�i֔�R%gU�*���������X   �8��d%�D�����������s@'?�r�3��W�N�L^/��ت
[&�7�����+U[��F��e�lgn���WT�7�ԩ��[�.?L�������Ǻx�0��K��s�����M�ϸ���>�`��5[U\�1Z���V��ڷ�7�4N��t�Q�C�T}����:S�-A��ru��X�oCݔ��X�7j�o��e�`�.�+,Q��$�:��(�>��P���w��l����k������[��|��%�j�=�V��բ1~�֧�{Å2�M{��N������   ��"�   �ò;b�Mnw��K��}ll�Z�H
   @���c���-o;\h�mڪ��J������Z��~-;M�͟�!���@�����q��u�?y���7[<ƳK�[�>�Tk.�w���J������+��&����� �i�;�o�V�:���&Du����N���RGaZ��{���W3&��s��&����{��=}�[�n�sk+s�4Pz���	����7Z�j�x.p��zӚٜ'��t�{����ie���-��х�tѸM�W[u�oz���ۄ~[���7��j��6�5�X�m�
�nAN  �H���84�9�   ���xEǤ��r��\�j   �x��6���#��*��5Ǐ��4LKܶ��4a�[gL�Bb�	�������ڭV(�TQ��N�BE����k7j��	d���Jw�_k��&�h2����C�W�����iWڑ�}f��	_M��?Z���'�=��h�*��y/{夯��.޾W;���>_����̦2�i�����=�`y��q��z`�2=}�9��s����߼�Hg�d��(�~v�q�ޜ�  ���rUUEfhtKHH�x���.W����A�   ��=3u�������m�T�A�[tl�5y�ݮ#?�����N   ��wJN?�|eu�\o+V/hj+��+7���c-�@���cVx�����SFY˦�Xc�>�&�=������3K���}����-TUMM����6�0TG�y�}�+����g��^]��A9yh_߲	���y�`�2N��ݷ<��ۘ�gU���n~����T��#�J���6yՆMw�y�y�)��Lݓk?�7,M�քo[b�g�}�mWm���p��o @����ݻwG\���r���$��>S/r��Ƴ���"�>    �n<q�5�։�=�5{
G���9be�L�p��8   �lC��}aü�ii��5L��}�
6WTi�����Z�y�/�gLԫUaA��7�w�ء��܏�`c}�On�ь϶����
S�ʹ=�����x�>b�UI�>Ӛ��#�H�jO 2�6�?��o�B���|h�r+�
ûgZ��k��!���U��
f����z-k�_����-MS�֧_�Q�:n@/�w��d��v�].k{M^��ܴL~{���q�;�����w�9_q���z+�s �EZ��������P"�>    m�p8�o�E"��v�U*   @�]��kS�`�chv�U��˄��[unٮ�:ˣ[ٚvɎ}�t �jś���#��z�+��Iu���7���3���Hy��  ��IDAT��8��`�	�ُ��;�{��L��*|�3϶#D�1�����9��3�g��[���6�U�Y�����N���qդ��ի[��{��HS1��3���nU��T|b�Z}�Hk����}�ky��  ��H	�;��)�[SS��2B}��`   b�.w�-�Z#X�b�)֞��:՞�v׸��L^&D)�o�z_Br�Fׯ�2L�   ���`f�)(��d$ԭ�+ ��+��
�y��T[Z�����γ�Z�&@W?�g������i����
$�3-iMp��m8\Z��l��~mxM�ގlg^��\�V7	_}��!�دG�m�)���;H�z}���WsN���*����:�����1C��W���`k��;�w��|�;F��-����X��bc�sǜ۳}Y  �i&�g�UV�rwK�ݡ	�y�;�G�/��   B잷[S������W�K   �@JO���\T��R��?N�?4�q���Sr\��ܖ �s�6�3�X��N��jK�[\���I#}���6�&̴p�M�Ǫ�v����U�ۧ�m��5ʪ�ze�utzo���_�b�����q����o�k|�m���z�~���K����}O/�� gZ����Vz��C%�z�����铭哇��I�ɴ�  M�ݻwX�}&�WR�P�W��}��:�}         ���~dQQ]�ǉ��8U��n�;�}�>�-&(֚B��
K���:uXE��V�ؿ�����[�>�4pmx�=�t��3��4�N��ʉ_����ZÄ����*��I��)9����h��>nBL�c�2HǺ?S���|˦�ce#Ǿ	��웬��ʂWM>&b�}�8�+�u&��-X�kO���y�T��e��Ԁ �N%��p���B�#��q�        aW�JVrlLP�~%�Ę�<N�_�0�-m	�v�&�g����`�����B�& �`Kp�~��ޟ/��*؍퓭�=3�n�a+�d��׳���?\�oO=����sNЩn������c��e�[���,�����^Z�Q7�8�Z6m�s�ӵ�@�"�Q�s �eJ\�1
�+�4�yn���\�>w��<�_w�s�`���%�  @��}��y�*�G��c!�        ®�^ة~�܀=NYݐNj|��@�B_\�÷�_ֶ ��k�Z�/��{g阞��žCV��˴�5����b��ɵ��.?\w��U-01��j��eoga�W��\�:�߷��>f��b�*TǺ?�V��jɎ}M������`�a�����T��~�.���em����~앚d-��)zkݗA;� �lL�oӦM*//�������l�k�`0�`noLL���B���C�        �]nqY��A�҂�8J�~H�����1�w�;F�mi����o�f}s�(k������U:�H{\#Xmx��Y��`߄���[���I~�����Վrv��t��j�����?���z	_�1�x�b����18HǺ��~=��/,���~[���*5�R��~3oQ���ۗ��`{�Ygy_Q�+ژ��|w��xƑ�3���� �� �U��v�йi���A;''GQ~_Љ���ڲeKP�6,GGdm/�F�        ���������g���d�q�.С�ruK�����Ȱ*� N[����%ۛ������f��rg��Gv�g�q7n;����Z�f��GJ��q�(M�ۺ��|��k��J��k?�J�i��TIG�ŕ�oUf~��_�ȴ�}{��1Kw쯳<�op�u/oP��'�O���0ǂi����$��̭�<6 �7&��{>/�����xj����q�����8^�]�I��5 N���r�,E���� �D�        @ؙ�ݖC��U~������V��@2��w��̑�e��~z�/�<�٣�Y^�mo��2-R7ȷB@��	����ۂ4��������ߝ?����ڣ�����H�o���+(L봧������z���8�
_U�>|���D�=�q@f��l*ę
C��@3!���d�+'���`��]���(�H�i�{+!&�j+�	q:~`/�r��Z�vl�s4U��gz���ֲ�����G鑅� ���5�{�+1�K���QZ|�*=�������҉a*vONT���E�oenQ�U@�B�        D�w�m�Гj�}�J�׏���[��y{�6_�ϸz��6�Le�����-WTi��=�z~&Xw��S���#��̇��[�I�`��gg���Z��6�����K��iu�-31����kwA`���.�~7o�;�ꗑ�oM	^�����uô1ּ����c�T���b��@8똁��?\Z�Ha΋��춪	I�1�5fH�[�^>iD�c��;�|y�&���	�;�Z����z* � �����7^�lk{�>P9���j���֙#ir�JO���fB�_�;��oԓ�ת���;v��9~���K�~U�͘���K+6�_��i՘ `        ��,\�N�k�v�	��ا����4��3g�F�u�	J�����9P��i��m�_�7��*�h퇯y~��r�+�����/UT�`M�DN�>���:S�U[�=�ҝ�u�߸�1�x�����k,�޾6��^^�Y?�1A���_�vꤠ���x���:��3�~����-.��*{^&t:���٪j=���=ߚ7U�.�q���<o����i�����V��5L%�[O�X线-X��h*a���O}�҄S�7}��JSq �*o�ݖ��.{�5}y�@��W�N��'���K�:��7��"���~KKw�orLS��T����J�1G��fM�5��O���{�W�@��        ����r�f�f-���×��K�+g����M��]C�ҏ
��������!���%��_hUx�I#t���eS=,�'S��T��V�2L�+���ɪ:��l���.y���w�I#[��/�f�߸S��r���7�
_�V��=q����4��f�.3�Z6���}��x�u�z`kM��S�2��Ҋ��:��H�Z�z��fk�[�}�i�����$^9yd��LU��y~���iq|��'��//h��w���6LK�@G��<�O�ܣ��j&7�4^~�L ��ii�]o�ϼ���Z�7�g*�.�u@+v�Z�rv�&��Ӈ��x����7\�Y���%;�w���Ϩ�3m�o��y}]dU4_\���;>:J�Ӓ����t��������       ����W�A���9���7��7�z������M��/:E�{{q�����%:��A�0����u�t�^Uaye��q��!��%�ֹ��s?֞ ������+�L�L��`�.m:����ږ˦�eG��ϛo�jBp���2��2�p��>��᫛O���֬���?Ԕ�����3F��q����<+$��X�z�1��'��7>�s����_M��[�M�д����ڶ�&0�w�V�9�Ha��}�]�}�%�v�V�4��T(�ͼEV������_.>�NHׄX�7罀?׻���z��	�^wd� Z�#����k��>]��,�B��ӳ����VP�T�3_v1A��� 0�_���O<��m ����+�
�浇�R��=�s�x}� D.�}         b�U��ϼ�Wn�@qGU���ҟ\m��LE��BO&�s ����)V����1��<�;7_bU.1�}>��U��k���[�h>5mrM�S��i���lUDӼ-IMX��٧�Gr�՞���rq���iCg���	s�U/�(�j�<��U��
9�z���^w�b��&l���W����1�Ա~��>��YS4�o��n7�>�6����G[�j��}ƕ�Gh�ˑ�3��ʵ����s���O�d'��G��<~@O�~�I�'�w�9Fo��Ai�h�}�[��WQ�T� �Ng����R��|�j\��Ͽ�wH���U-��
�8��fU��������i��h#�u7�?�_��X�]5�Z>�s?�}@d#�        "��m{u�#���ל�k�'-Y_z��h��lߧ��u��\&[g�g�j&�����:c5�y���=����?=���|-8Mp�_W�ԟ.��>85�TL���D����
��WA3�_�A7���^���hB|�9��6�n�Y��2A�|�G����R�	��-ͪ�g�2�3!�6������W�d*�z�eϱ~�U9�0-����5�y.[��pi�u�g%%�f�H3�{���JәJ�f��Wnj2<���oG^�u����;^[��V���>X��>��s,y�Qs�|t��V�ȥ���SPbU�땚d���&/���/������aK���EVu���G  ���>ccn^��3�~}�y�/�g����''��W��mr�~A��D6�}         ��V3���0�$�5r��:���7}Hkj��@�����_��jr��w������/������]��g�~m�	�����pY��>Q���~��E��㬩V��0�ܿjCL�ʴ�{b�ڠ>�P��m��9��XǺ��T*4Ǥ�qِ�*����R=���}r��u�yiŦ6??sl��b�U�0?'SY��U�i�p��,��ϟ�~~�=������1&<a*���s}���y�?L ���,����[X�On������Ws�]�o7��D6�}         "��/�O��q}�u��tJN?_�Ƭ�X�}�ު�w���E���p�U5��a����&4��G(�=뿾v�U!�PI��z&,f��k��fLЬ�C����τ(_\�Q�p����-��+Sτ&��n�&�׭�c}ݾ�z�s��Y��j��������^�k�����`�a��Fb��x�/����֔cu���;[�eLC�o�]�^O/Y�j�K�`*N��i� h^KC}�,�g�L��7��ִ���+���L�z�O��+ ��`        �h+v��Ͼm�sF��f}������8U���/���Q+v�*�3�V&d&�;n@O�]�	W%�D�pi���b�!m>�ߦ��Y�]i?�����o���G��oVXS[�}��9���kL�,�iU�K��QaE��J+� ��}[�J� ۳��1g��2�^{��v���g�Y��1=�)'��X7mz�5.�c�k�aϱ���u�7���R=~���f[�m&t����!7�]c�6��x�5e''hb�֥�\n�r��<�s��ֻ��3~��|kjslf��! �וC}}Ғ���^��oCL��T�3�]����=���zm�֣�3��u�Tk޼�0U����60���Qp���.�`        �L�7SI�L�d>�L
w�R�	��	���ڽ��	�c��&�  �xZ�����~��)r�k��.ٱOk�lp=�~��'_�s�<O=R��7α�Pb��b*`�/M���+&���,PQ]��}���xl��ݶ��n@]%�G�            ����f����[������o��p=���X�oO9Vg�`M��)���Z���Uu��J��           @D�꡾q}����V[�O?{�#��sP��-U'�~)�e�kFNm؟���T�j")D�.�#�           ���꡾czv������hk�/,���4{��'��/>�
�U9�ؒ5Z��7��J��q}�u��4 3U��?]����UO����R	��           @Xu�P���Wn�@	q��>]��{�f�7e`/=p�9�6.-���Ws��cB~�.\�'�>K3G����y���:�.�#�           ���꡾A����(+)�Z~�������nA��;Κb�����[|T�ϫܳ���;Z��k��맍�CVXU�������            ,�z��_F�g�/P��Dk���t���ՂT_bl���˷��_6�~Ay��߸C��Q�á�C���th�8�G�            !��C}�R�4���'-�Z~u���^����<2�}��L0����{�J|��0!��u�p�>            �TW��P�k7^�����k���g���j���N߼�&%�ƨ�����d&���+�^�P:a��`            B���������hp�4ky޺m��S��iy���/�P�g�H��Mܧ�v���~�卹�:�N�#�           ����>�{�������;�������V��r�����t�pk�3���WY����r�d�LM���i�}�t���6lXP�NHHPee�"Iff�GP�NLLPEEdmoPt�p�>            ]W�_v�F�̴�M0�`I��0�f�z�A=�h�Q��?�s]0v�U��4���u�;��M;���������N�Yc�����y�Z]!0�JJJ�`������P�������JKK��`)**�lo�:�N�#�           ��"�W+�H�\�n��#����ښ��6���9��KO��}�{d��_?ۺ���FqQGW�ۂ��g_(��P_UUU�'%%U6�ϡ� �a7��N�S����b]���       ��둒���i`f�l6  ��q���P��,۠å�-����za�F��wH?<u��5X�G�|�C}���*���~�"Y�B}^�ɵa�p��B����:�}         �&�練�;_)q1  @�sی�:�ї�žCͮK���3z1(��wX�zz��ٳ���'{^oǪ��i�0M+���
E�P�ܼ�����p���Zwz8�G�        �������O'�  ЁuK�׃�OՌ��iv�W	���i��|W�5u4�
�y�p���Jv�����T�p_�"�        B&';C���	   ���ݭj|��eM�7 #���	��(--k��+Tmj���"���            ���0����JE�`��"%��e�}��za!�HC�        �̦y�z���}   �i��\���|���	�uq�r���-R*֗��j�!�:P��`        �aэϽ���;_)q1  @�s��\7��~��ٕ_,t]N�Ӛ"U\\���K��n&���>�����noD� �>�}         ���ا�|J�����4��   "_��mU_��l���h�.";��mo�� �>�}         ����.     a��>�}             ��'��}�              ]S����             ����             tm�#�             @���             `DH��`              ^�#�             ��0���             P_�}�              hH��}�              hL�}�              hJ��}�              hN�}�              h����             �R!��             �5��#�             ]����fZ)��>�}             B*&&F��媪�R$2A���������r�(11Ih� ���            �>}�h���v3������L5�H�^�+--%��A��            �vs�\*--	�������>@��}�             �M��݂���%�p��            V���*����%�4
��            v�
��:����%�T��            BvW�ϫ�mo���p�>             #Ta7�;2Bn��^B}aЎp�>             ń�6mڤ������JE�޽{k˖-*++��111������R��#�             �i���A;''GQQE
�ͦ��+�Æ��ሜ��r��#�             @0�2�G�            ��(�2����*���kbl��''Z�(NkW Ђq.D�V���            !2{�0���]c�dkx��'�չ���R���㟮��M;[<n\t�n:i�.�0BC��|�WT鍵[��˴!7O@�ƹ�{��Ա��it�l�ꙩ���U{��+�Z�#�            ��#��!�����i�:w�`kzq�F�4�=UV�49��T���y�=�ے�bt���56G��4_�}�^@$��eg�aܹ��5����p4x{i�S��>�}            @�m>���{Z�r�dڐ�MOִ�}�?#�Z�qìෟ���8��z��_SNv��|��\�/Z�M�yJK��Ecs4uPo�y�p���_T�ZQ	�-�jz=�A�߹p��5�U�%���FC}��p�>             D��m-ܺ�
�5�T0��)u�YS�e����U�l��׿m�D_�o��B�������w�c���]gOխ����v��)��ǧUU�t@ �̹�ɗM���<Awz�_Ü����9�yEV`v��Z���U���sNP�j"�G�            ��Vlj���[���T��f�Q����>fP��>Ӫ��ic|˷��~�P�ׯ�Z�������ݪ�vŤzr�Z��ߕ͟���\��u���g{.�����*wV׹.=!N��p�>             ¼�n�/��+-��uN�_�ѵ�{�-�\��v둏W�W�i-��g��Q���6_��WjR����u(���            ����?TR��:���7A����~���l�:��R�cUX^) �U��υ2uZ��}�            �s�����{6������e;�79�	�m:����3��4�s����
�t��XW�=�N�/�G�            ���ލ����19��μ"��j�Q�yVӐ�4���Å͎��3�	�#zd�CD3���'��ZG���������p�� �            ���#�gj�5oZ��IK��!}4�H���.}l�ʝ�G�71&F	1Ѿ彅%�>�>�u�''
��υ�iI:iH_߹`����s��"�            ��w���IC�u���r���E��lC�A�Ę�����ʪ�����h��FϹpr#��o�-��o�R�>�`            A2�u�9'�GJ��}��5��։���W�r7�N}�5�yS��t���4��dc�BgE�            �+�|CQv�5o�z2Rt�ȁ���c�v�?=�8���M_���r��u�[��sxư�lG�S_����)�|�u��Y�\H���΅c=������>             J*�|���WX�E����Ek4��4 3U���O�G��s_���Fl���V�q�_E�J*�D��ʯ�g�s�OW��\h��sa�=��Ju�            ��3�Hߝ����E���'�?*�WR�T�˥�#Uβ���5%+)�7�WV! ���/�s.|�s.<�p��B�>�}            @����=�_T�)�Ꝗ�>�iwA��v��~�HC�Ҭes{s�>3�צy:�s�Wj�u���_gG�            �@�K˭0��#Խ݄���ѽ�� TcLe�czf����;,���s.��z�K�            @�9�6�:�����Y�y��>f�5Ґ>z�㕍�7�%�D[�������Q�Bi���}            @��9r���yӂ�@I�Q��ŗ�����l:m� ���iYڐ�'��Ϳ�j�����\��9r�K��            Bࢱ9zo��W6��������3|��.]/����v���U��q�v�q�I��So��tلּy�~�ZAzz�����UYY�H�����M�lo�"E�υ�74x.tF�            ��~�=8�T��~�>ٺG��TTQ%�SꙒhUܛ>���9Ъ�gl���,kt�߼�H����X}m�=y����ۋ��@��cct�a���Ӭv����)�,r^�)..��}f
���B*���}{Ͷ�m��5p.W:�r�=6����?ot�ѽ���)�ֹnHV�o~�g�?$h�
���3E"�}          ���w����q��}�֖�R��\��������6�M5.��j\���P�ʣ���ƭY�U��) �b�u����Ԝ�w�וO������m;\����M=��s���=Ě�=�S���:�J}�Z�	�9���e���j]�;�gB�������퍔p_k΅e;su��5y.��H�5Ǐj�v�����	�          '.Jr����Y��8��F����
�����<�K��ױɽ����3���T���E{V��m��꟟��*��0���%5�;w��\=�x��Y�N5����6�҉�=�ߝ?ݪ�g������*��]�9�6(ҙP_UU�B%��P���"%��υ���9�z΅�f΅/�BO/��E�BgB�          :�g����B{q���h5�Qx�#F���7.�n�/LZZY :��Vl�&�+w@F��''(3)A	q*����N��Vaye��6�K�k���핥�Dk�y�Z��:�P���L���;XPP��Ue��"!��ߕ��)���kk�*�UgA�          :��+4 ���{X��j�Tcs�e��e�R\T�2<�91 ���1��f
��%嚿i�:�p�����S��P��½�&�gBu�nC�s��#�          �T�#ں4��L;hw�����Jng��cR#2��r� �u�;��e�}&hVX�p_�lo���i�  @��yEm�	}Yj��&ב?4      2��wp�d������t%%g�f���i�6���| ��H	�y���V�V�/�p_�"�  :���B�[:W�\\Q1�r�eBx͈�L���rٴ�̡�8�b[�n{u�l�w�C���Vay�2�\J�ru{eu�>�]��j     t96�M��r��U�,Ue�>��WbR�RR���UE����.*�@WPZZQ!7/o�/��nwą��L��T*Dd!�   �rӄ4�K���mvG����R�|�C�%r��wg����^��7�-a��d��~����*)���z�ڴ�/�    �.*:.]�1�2���U%�*?���\�lJN�
���SuU�  ��	�9��ۡ+..�
�J�oo|||@��G�   @�\5��T��ڪwnվ�3��l���0]���$tW���      �d��X�=�=ZG�ui7�g�\��޿�ج��sH%E����U\Bx��	 ��Z��Mp���l   �z�$j�ȁA���R/��l͟1b�z�&�n[�c���;��1��5��k��}ڰ���E���J����U9�2����<�f��zŦiHB��b    @�x�n�6z�Gnrɶ��r�ɮ"��^쮩v�mQ��(w��J����-�p��96���}�@��'�Vb��V�'6���n�J�v�=X����   ��  �����.���7����}��j��_u�yE�z�3*�ly��I�{�kΕ�^;���R���*�J�-J��q�n��mw(����4E�    ᖶ{�5����ƩJ������������\�Sl�͐�}��v� E\B��š��ved��-   ��>    >޲[�/Z�oO=�Z�;Ϛ�����E���r��٧�B}��/����J�R����n�\ժ��Va�~%��� [��a䪩     4�nw���\���)����K���+�ӭ=fzD7�%6-Fgx���<�C����>r�����-JJ��9��б1�;��   Xx�  �.��Y���]�a��oz�o��ʩ�e��ooaI����D��~)��u'���5[���=͎�˙S4�{�o�٥����(6��]%*��R5.��UbR���3jo���<���     �Lu>��T������fE���>xKe���g>�#�]s��I�h�)Y �|q3!e�l�]*+ީ��2���[�%$�QTt�o�������'  @GG�   ]��;�k�=�nv���	�x׵����v�'�h��TV�{/���7\h��{���7ے״����q�eӂ��s?R84�����V���Y*ge�*J���䐲����jΪ"����ܮ    ��K��uwai�s��N�Aٟo���Iʭ��Ar���6�lI�nV�/��b�2��"�ۥ��ed���m6�����4;  �� �   ��i����5�֔��䍔�ͱۣe�L��DEǤX�u'�QuU�ʊw+��6ef���]5�r��    �Sn�=���y��?*U(���<��]�?z��Ꚛ�{ވ^- ����~����[�mPUe��zSll�   X�   ���kuJN?�L���j�{�Yu[�>�t]X[��^BRo+�gwx&{�5�P`�\���x�oQA�.�g�    ��s����5����BE���y����)���Y����-*oH� ��>�Ȝ[�)���_H  @��   B��ʩ��~�-yM�O�ۂ�s?V8�of�&d��>vG����(o��
r���]    ����[,���zqv�"\����K�ɣ�k�+��H Ħ��D�\%*-)Rjz�   X�   �0h�%oC-xM0�Z����*�ۮ�"��SZ    D ���l�����|u ������/I���J�{$�C �-%}��K��h���c�$   �>    L�j��P�w�oWGf�����UQ�.,/����Q��$!)C���_�%��.    @dp����r�,���M�l��{�������ٞ�I��.Q�	JN�jg��mQbJ_%&e   �A�   ��Z����ׂ7P�cS���Pi�N�]�;j+��t��|^��     r��Z宙�w����+��ֹi��?��͵�l��N6�e�\nTq�U;+���S   h?�}   @5Ԓ��k��iZ�6Īܗ1B%�U]]�ظT��&���P�iY�����r�    /�[+�q'�Y�l;��{o�(�����{�M�h1�7��$���w�J�����H�=rd��  ��#�   �Y���Q~��:Cކ�?��%f)**N���:��^��"E9����    D �{k�=ꬢN��*���e����gv��]j� �HS_�LLh}���`�vo_�n݇(>�   mE�   3Ӓ�֗��.�s��������mHBR�7�m�*�j�'    @p����:�쾛���*���Sn���mn='���n�	Y��IRl�n��(�#�
�EG�7��F��������ҳ\-��:��v�,�'   �   "��nG{��ͻT؉Z�6%.!S.�Sy���go��    a�)�uU��}�N���[^H���ђ���x%�Ul|�J��(w�j��JM뭄�4UW���h�l6�6�l�_:��Zw�K�   �>    ��e����N;��K'�>�B���Ug���K1��:|p���٠n�    n��{oy_]DaR��)��Sl6����tEǦ)1�Pe�*.ت�<�l�(�8Ke�K	��)�	  ��}   @�N��>MI�1ֲ���H{Zs���i�=�
g�:3�ͮ��d��P��mV�/�G��U/     D������~����]Q����[�J�R7󷝘�4kJJ����HUy��v5���e��   �   �����1�>��o���TfR�.�0�Z�����q��z�u�ٞ��Tph���Z��G��     ��R���������������[�' (�X�&d����-�g��  �n��K �j���   ��)�󬩾�yE��;�e�[a�^�I��7�4^��ޢ�rՙ8���wD�*%c�J
�k��U������g�>��(ϵ�߳U}e�]r����fll����	)�BBL�!'��IrR �G	�w0����p��r�-���J��팬�E��J��Ǡ�ݙww�^����y�    hc���»oި.��/7�+m��S�͸�<�dE�!��*�V�8ư� t>�O��媨��YA����V�:߲�2�B!9Q$Qrr���   �`�ٽ���J�WW��^��g�QIEu������S�=�^w�=p�tM��IUT��x����׷E{ש ?A��F��r7�xӌ��2���"    �Ԛ���V�f�.��������=4�����J�s`�T$\�H�Rftq�U�� tYYYھ}���}V�/,n�`�U/;;[�����E"a����s.J   �����jҐ����,���Ŷ�X�IO}�:֒wx��tڱ��[���p��JI"�?_%E�ھ�%$uSf�A���u���w��3�p���)\Y     @�LEf��۝��b(��O���<���%�w�r���b�x<*+�' @��p_M���8-�W���   ���̀~1���vnA�~���#���KҒ��i�iZ�=O]�!b�|	�J,٣��]v���MRJjO%%�ʭ��-ZjڴT��W	    Р�E۲�l�;�{#����7Љ�\.�R���<'�>? @�pJ��*$�}�X����9�>   �Y-x���I>o춟<���G^��UҒ��r鯗M�i��Ve8���0�JL飄�^
��SE�>�oQQ��pU���81�/��q�z    _1d�V�^l��iM`��磫�p8�/Q����S����>d-'�"��s��տ��盘\�9�]VU?S �Υ��}�����>B}�G�   hG�O����ƶ���J��zK��ޒ��=��)�t�{��+2���=�%%R�b�ʂ;j�������	    P��SL|B8DD����"�����s��?�W^5Oa��Cn��rJ��*�q�W!=�a*�S���v�_N� :��
��w��FG���@}i)�>�#�   �������3�j����D�x�������i�{[t+�zw��2+���w�;����    �n����R8D�_n�4p��524\���/��. �Si�p_G��j�w��P_� �   ��������W/�oy�}�5|QZT:�%���ֽ�Nӌ�>�p�k:�py���W�H(�T�W�_�    �0Cƿ�Z�2�~�   �]{��::�W���}����>   ��x�M��+��ܗk5g��FxK����5'��-QWf��MH�u��i�PD�e�T��\    �#�Ҋ�;o�R�U�������>  �b��֮]����6������9�o�p_[����S(Ծ-��2�   �66�W�~:������2���M�𖼳Ι�7Wm֦}�¡\.�<��j�_    �:�zC�S�_n��y�j�!   t���"�[��M���ɑ�㖓j���m2���9r��u���>   �U������.���6��V���M�zt�%����� ��;�Z~�aȉ�����    Nb�{B�L�]"�   ���   ���T��Ӭc�"�6��V{.VK��>����������*���-8�6��#��A�ʪH�{�m���JJR���pDr�Fת    ]��*o���P?CV��:  �!�8@��$%�<���w�4�����{��(-���P��KU^Zs.X�"�Ғ�q�x{��!��   `�����E    �.�����{c�P�J�=�k�F8  h]�O���zilV�읩@����� Ҽ�zd�2��zK����Q�t�Q�5.��R|��*�-�ݣ'��W��s!�3k-#�s!�s��q���_�7�W7��}�쳯�L�ݦ�?^�O6���        �b�\%4�����J�9����  �J�|�\Fݝp�j{g5�^�_�V�=�U��{���x\N�cy�.7���|�1���^�����ௗM���:s�[R����z/39ў/����>^�����"-)	���        t1��5B�2�F�}�   Zٚ��Z�#�n��;�XmC��S4yH�e�}� �{��ߨu�>iɱ���*}�y��n�Ӟ`�x'��ԡ���VE�׮�H3�{N���p
k.,۱W{�K�=jXA��;�i�ν���[V��R5uX?�	�����Ǩ*�/^�'�"�        �嘫�F2�F�E�  ������߸��ƪ�w�4�������yu�]�g��x���|���CG�?qP_=��s�=%ѮX6���t����hW?��\�����9��m{.D�?ٴ�}�+B����������:�����N�Nko_7e���L��ʉ�        t1.�{��8��M���  h�����~���]�.҄��t��!�mg5��`���Ӛ=�����M;������.���*~9=�ف@�#5f.����ѹ�[�]=�����J**�����
�u�+�}��e�9P��DND�        ��1�p��(�a�  ���b����)��zw~�Ʋ���ڵO#{g��c�{�C�x}��X��o E-a�`߈�g�Zc��D�        ��1�"��hf�{E�  ���Ae���hU����`_��' ^D"ͅ`��B������xm�`        @�A�Q\R�) ~Y�Ss��_�Te&'�2���-߹Wo�ޢ`E��c7���}����{������FD�C��${ݪ,���D ��M1 �n��m�A������3��6b`l}َ��7}�W�-o���V�        t1��C	�Ɗ��\|�_������̘��=��ܯ�*�'�����@{����4է{l���W�O���q7�2^W;�^��S��S�V	 P7W��uS���19����"��d]��<�o�^�����g�wp:k.�p�X]4���������ۥ_�u�&�ko/�ݣ���ʩ�        t1�pE��(��F���j���o��Ӈ8������]T�D�W}����{ܺj�h}}�0]��}�a{�����u���k��} 4ϙ#F/W�4�HJPVz���ְ���6�+�e����ʪf?�����I��W��W^#�@{�m.�<4[9=���7a.|}�0��z��D{�i#(;��bU��s젫S�        �b��`_c�J�>�	���Wp����ao[�S�{�
=4o�!m������/gL��@O���5蛏α��6�UEǪzc�� h�2��a����ju~��z���*oA���1&ɲ��*�W�	p�FNO�e.䗖������\hJ���3O�����X���^Y�^�ሜ�`        @c�T�Q��{��q�%��B}V��|�֠^�"d��}m�F={��:~@%x�z�gj�_�Ў�`��eC�@��Q��vv6�� ZSfr�~s�d�MOџ������#�s&��V��j��[P, ^X��~�Yѹ�̅V�?\0U=S����rp�>�}         ]M$�l�qL3��_8܅cst�1Cc��{�����U�҇_ч7]��i����}�s|���}�Yg�d��:g�f���  Mw壯��~����h`����隓�QZ�O?�~�F��Է�9��-C�6��}������>�+7	p�+�#��e�<�>0n��B���ft�4f.�~��rx���jh�t�;z��s�h�5��6EC������r*�}      hS�[�+s�R �c�t����~"9B�. �p��������u�Uy�/����w��}֨�vۺ�{��{ܛ�6�̑u⠾:q`�u�`��b�  McUQ���N�UT�O6��#���^�A��3z��?y��hq�ǵ~7?u�yv@�r���z��%�����:������F������_�-���� >Z��~�\/_{��B�Fo{e�z9�>      �)�L�* �fFZ�Jh*��Z�E_��P�N7&���f��m���M:��U��fw���ʰT~�����9�<�������.��u�D��j�����8b�����ok�u��?�:Nkd��	�{�٫��d�����;u绋ģ#��)�[�Bw��}�����3�Ǜ:�`         ��4��B��n���a��8���}c��hq�&�������'��'�j�16��[�6댑5�w�.?BO.Z% @똿q�]��wZ���S�H�CN�9&������&����>�B�y}��xv�\�HQvt>l�_��zu�U�#�]߯�|n�Bᰜ�`        @c�с�J/�}S�P'��, 7�wl}і]���c�V(��q����7���ȴ�2;h�n�q ���WRf��,i�>��WoV����_��D����%�ūW`��!s!��o~��z�b�� �˰�[�J����`        @�c�#nY��9B=�Ӣ�+N�+5)��qo������֭�5�ɉ�Ql�e;���u�hl��uK��N:F���  -g��J}5����7�g7�|����ߖ��_f�:�#�BI�Z"-���� �U����BND�        �2�*�}9]@�HJ��7���Ï�*�4&�g�������ځ�����>[���  -s֨���{V��=��Z��=]���B�<��ק+tˋ��4t
������wű#�jÖ/sw+���B�        �2d��2S�U`�=�$3G@���Ԩ�4�i�Z��|W��ݰ�@�/\��:q�])��S��wo~" ��.7\o�٢�����7�/�}�i��'��5�7 #M������~?y��N��֭���&c'%%���Y��222��|
9�|/��w�lm�\X]���7�����Wi�����Yg�t�x��T�         ������'���υ#�2�E^ċ����&��5FM��%���~�?���.�0B�^���:N��T��K 8�Փ��=����Vm���۵%�H��J�#���WZ����#�*��ޝ���]T�x�}�X��򪰪���yѩ>�����k�d�`��YK[0MSEEEѥPNP\\ܥ���Ict�Ӛ4�D��,�u���y�~���r�n�iW��Ƴ͊�g�_��h�Yc��v�K�"�   �����a���71�[�VB�!�6��ZU ��S��!e&D��qEUX�U^%    �L�[�/�ja���H�!N\馦bSS�	z\~iӂ}��J���K��S�+���-ӎ�O_|_ �#Y!�3�^�p�.]���U������z�ǭoT���tr��
��Bm���0�kaa�:�ꫬ�T[��3--�^wJ��)sa���\�G�s�H���	#�!�Y�EW=���^�S�   `�~B@cSw�z���׀�W�ӂ��[�و���G�R���?M��@u��[���~�`��Z��~����    ]�a�Wh֬[u��m��i�I�安2�6=Ѐ6�8w�f�d����٬1�e���o�[����Z��IY�x������?�R��9#8  N�м%�YԤ!�ꑒX�>V��/��֣�,��V::x��#�w�갛���V{��jԄ-��®V�yg��1PgQ���u��M����ezi�:9�>    ��+T*R�Y]��T���U��8�z��럘���^��     G3����oJ�1Fĸ�j}�'�n��Ú��R�Ԥ&���>r`l�jK�V���>�B��y��n�~>�D]��� |���k���������;;39Ѯ4V�Ԟ��ܵOE�X���?ԙ�w��FZZu徂����g�o{���p�U1��j䀌4��pK��?,��m�̀zD�V��x��,�:0^i�����Żl   �֋����ջO(�_�[�\�+_�Jʚ�8��d��}b�;
�zk��&�sT��:n@�����b�lx[ٽ�]%'�R�7I!�K�e��Tx���#D_��&�T��/    @�0�Y����o��r�]#
�#�7n��|V8��r�Ǎ���5V��4�>�l��T��뇋u��1v坋����� �HV%���
��:*�W#5��Q{��:�|��gْ_d/�!�\��K�#�   0�_/�}�iM:ƺ(x���zd�2�6.䷳�D�}�	�'�,U��θ�Y��xc%��z�s�O0Y�? ���jK��|u3<
x�ǐ�r���+1!]^B}    _cHZ���E�S���ϣ_\�HEUX�D�3c��=��c��k��6�/�j-�w��;k����`EHw��P����bά�OR^�i� ]OG��jX�>�=��¶�9�|��Ñ�   -0�{�~~扺v�]��;z}����_Z���OO^u��m����˦i��O��m�;Ι�Y��T�6䪭%�j��0eD�W�0�K��|�$�d�SD�q    Nf���f��%�~U������c*r��Ë8��GKtű#5�{�R�>=w�����^ԞZ��򬉚1j��n����-a}�GS�);=U�F��NP1 �v�r���V��K[���v�����`   P�܂b��;����2�-)A9=3�u�����D=���u�c���e�
 Z��.�0���;S?;��1w~��N���N<:�m����܏���?��
�7*�\n��S2�����|C$T����    �khZq�O��ߨ�2�5���5�[@�*�]���������qkd�L}x�������u���`s�������:w���m�}���_����������T�]:�޶  ��i!�V����������}.E���`   P+�w���z_�ףK��[�tOI�o�*��s���h}�
�*�����a�b-yo8e��D����V�{/����>=mU
,��T{h�
_rjo;�WUY�ʊ��lWIp�z�� l��E*CEڱi��H�*!   @�f�~r��w��p9�N(p�=ߋ~NǬ�+���z��s�#%�������L���S�ٖ]�S\"�ǭ�=3tt���zw��x���6֓�V�S&(�g7 P+�VY�>�o4�ߟ`��Z����ߪ狖#�   4Cye��l�>޸]��x�����V5��8Z�����1�Ӓ��Z�6���ʈ.no���4�2d�d�*T���\��mRf�!�ޞ7���    �a�+�D��zX�<3]�^ڥ>!�q���p��Z�3�l�NM��I�v�	��q#�9��>b@���ٝ�Y�}�7Vnj������7��>[  ԥ��L�sh�}   @l�[�{��\�:���[$mL��Ҕ�������ڞ��^RJ��s����g��سn��J�$�x�z�oS���    8�!�Դ~;~Q$ݮ�b�,OUPOF�c3t;����w���|�3F����7=E�ɉ��
+/X�e;��֪͚�a��"5ƿ?[�^�O싎ѐW������DI>o�U;�	   #�   ��ܕ�	��Ѥ�Ӓ������-���ȟԳIǸ�>�t����**ح��^    8�!�W�[�����7��. -������:�܂b=�`����>Zܤ���aY�B   4�>   ����/:d;39��5��zcZ�:�oc��	JM����*.2��ִp     �r)y<��wO.��O֩K���+E~J^    NC�   h�ϡ/��F��j�ג���Z�n�/ү�o��`U�KK梨�m�+���Rnw��.)%C~�W�F��.�K    �b=���f�O�Tz��;�	f�s���b��   �9�   -4�w�!ۛ�����}o�V�wX�=��J*ڷok��
d�UR�U�H�\������a���    ���1��r��xש��o*P'�6���LE^6d�    D�   h�o�p�!���֬qjk����/��ֈ����+�e�Tp�UU�ɟ�ߟ���B�{�0\�۫�D    �X�����5/���3��xc|_��y�)����H    8�>   ��>�]2nxl�2���/m�x���=8Էy_�f�-xkc��{��I�?����^�ʊ"y�RJZ/    �Ð��
�ԟ�5��O7�Q�r������   ���   ꐖ������'��::���q�HM�}�}w��Hk��o��Z-yO�鯞�I��"���yG���l�[����v��b�!E�U��x_    �(z�6Ј���2�ʢ?����ͬY�����ѓq	    �`   P�+�e/�a��}�?��i�739A�	�Cn�Y��-;�Y%$e*�T����    �����F���-&ޢ����O���xvw��O:K    '�   -��ڭ�����r۞��v��eӕ�=��zVz�f�~�~��'ꌒR���h_�*�ھZ�{    ��C�nHK)�����a�,���7=}�}    q�`   �B��di��~��n�8�0������jo:�X��l���ث��0\��S�6P�6���sb�z    ��^;٭����w?�+��O���� ����u�)]"    �C�   �:<��b���m��^��d�Х��	#��q��v���L�xw���ُ7�W��g����ʝ�t�_�˧��^�K�l�N����"uF��=��6T�w�vn[�^Y#�v{    p"�kU�H��Z�����0������PG>���������º��^f
    ��>   ���S;
�����z��ez����\�>�/Κ�/s�حy���r��˦�AA�ܻ����Ŷ�:g�`�;��5혬����	��;�*++k���(-c�����c�e����t    ��0�2��҂��̻�������ۯ-m�����?�ޙ2C�D�P��   �;�}   @3-ۑ��{]/_{����Vž�/��	���JC�j�N�	�{Ŷ����v��r�����Y�HJ��o�~��,ߠ5���Yy����׷E{ש ?A��F��r7�xӌ��2���"    �G�Ҹ_�������9{Nt����}���K�m���(.</zQ�툩����A�   @�@�   h������W��cG��})vH�o}��1����qBl{}^�~��{�Ku����+g��~��n�{�}��U;+�˫��!���UR���[�PBR7e��E"a���f�L3\�D���"rR��@    ��u��%�+�K�����ͳ�c��>���}���l�n�o�i�O�H�*Xx�#��A   �3!�   ��/���YGV �oo[����_��`Y��Z-x�v���Ӵ[�WV��s_��c��Z�ۿ��?i��h�:7C��L�ҕX�G%Ż쀟Ǜ��ԞJJN�[�����y砢~F�J    ��cFv��UѯWUE"J�9{s��m�Ls�)cu�����"��(0�U�n���e&+�gf2D�ˉ���=*b�� 9>    ��>   ��� ���-�[�Z�|^]?u�f��q���<�X����~(:�'�j/^����	��GJ�����Oқ�6k���_��0�JL飄�^
��SE�>�oQQ��pU��{W�I~y<�k�    ��4P�bgV��L��mʈ��U����{�o    �*�   ����wݔ�J����k&��>��ު}��v��i�Ŷ���7o,�s��ѱn{��XK�D�G�\r��{�+��%�K����)T�_e�ڃ�.�G.�O        ��"����0{iM]�|�2�   �V���\�~�ܮ�gi�j�Ղ��K��箮0g�n|�]�TT��8VK����joO���N<Z�,X���
���������        ��������^��4M%%%��x>�O���=�H$����9�   �������'�o������Ym{n�k��[��Q�s��i��XK��ϙ��VmVnA����Qbr���f(�T�W�_�        8�U.++K۷ow\��
��ŭ�s��Z�KJJ�9�>   ���..տ���}������C7�vll{WQ�~=���~�9�%oj�O�]6M_��.Ӓ��՚7!���[܆"*/ۥ���        �䴰�iF�l|�|sss
��ա��;_4�>   �������	G�Z�^���q���ϐ��s��並�i����=eX?]>a��\�J�\.�<�B~        gsJ���C}5����#��l�   �V���X�~�FW7��>�j���8A��d��j�*��bc����w�T��n�v�����K�;������        @�::��^���#��|�   ��_��^Z�GO�m/��c�|{iVK�a��j-�B>y#�ߧү���Cn�{<r����G�K8�mV�*9mH�������֑        ���}���Q�p8������   ������"        �c���3��Q����#�?�            p��
�ut��F{�/���B�            ��Xa��kת���M���}���>V����׫���M���|
��s�h�>             �STT�u�ֵ��999�x�r
�0TPP`������9r��s�h�>              �`            �A<nuOIR�ϣ��v��4t9̅C�            ��eFh\vO��.#{g*��?��²
�ې�G,�;k���~0y�.?vdl�����L�<FD�Bz��?�}�d�5��oy�}-ںKNE�            h'\>].è�~+�w��!���⵺����*������M�>w�]���{8���M���zsaD��.�������            ���=��t{���UT�D�GY�)�<$[�2�>�͑{���h��Vp�KN?$�8պ��Z�ۺsa��=��-.���            ���������� Sm�Pލ�NЬ�O��/����-�'�w6�1N:F'�k���r�.?\��\�D�s�S����L�����R}�iG�cO��Y��M�t�$�            �v�����1M���"M��K�b�v�Q����-U�:{����Z�i�>8Rc����}��u���s�lk.4"���            ���b����)�>NS�ߧ�ť�ū�c ����c�����υxg����|�8V��O~wD]QU��+�+          @�����W\ڨc.?v���`�����*(��"���B�qs�3��}%%%�p��е��
v�`_8�*�}          йL?г,۱���{�&�w�l��Y�A//]/�3�6b`l}َ�F�2�'�U^Vi�R�V�            �CXa�릌Ӆcr���Eziɺ���S����²
�����5~8e�.��\xqq�s�����k�����vIE�>ݲS�,]�����~NG�            � g��>�{�
�e��jʰl��;mK~�.��+*���w�sF�c��뿜3O��Jē����C��ӳis���a��N�{uZN{�y�q�޿��g[v���            ���wx ɲ��Lw�]�g�X�`�)���_.<�^�p}��l��x���\8����_Z������3Mi��<m�+��Ve�>i�vH���`�n�z�����-��T�             �LN�oΛ���)��۟�2�s��F�띖l��~�ܻv�	�,��}�9w���Ssᡏ�荕��������.C�8v���)v���[�r����c�ph[^�}            @�����q�z�ף���%��'���~6�x�o�s�"�$��j�<�({��o~��{ģ+�#��e�>R�s�Vk.��oF�L������/�s�pĴ�Yn�/�K����럑�KǏpl�K�}            @V���(��[�~�i�Y�L���B���C���c��G�96����O�aH�s����W%�_m�1�>j���΅>j���G�s���u��#����            аm���������.��<u�����kW5�Z�^��۪��ݢ�WG̅S���y�[�r��eb��Q}�˩�            3�v�jY�de��*;�����=���2���Eu��s�b뗌�s�b�o�_���|R��<�R�`����y��� �"�            8о�2;�dIK�IG��vJO�7j<��m/�²�8�!s!���m~�/�獭��*�T�             ��{V����e�ܿp�.��F����e�o�/җ�v��y��8�s��e?�'�[�V���`[#�         �aL��3��-��Z���w1͖�rE��P)
 �s֨��J|V��=��C���/u#ƹ�QYu��������ē�����f�������cb���&�"�         �q�p�	-��)��5s�Z�_�>V�I-�,l��
 ��K��VoVAYE��M��Kw_|Zl����Z%Wo�u��Ç��؉�	
�Br����6<����V�).���Woi�\xr��Z�cs�Κ-*�g��)�z�g�O ��.�
�_���S�         �0����V�y�;��Z<�����i-���YA
 h/WO:F�/9Mo�ڬ�vحq��
G"�HQ��dM��3F�˨n��fw��zw���`0h���-�������R('(..�R�{��1���[m.|w�h������}h�g�w��X��d���#�v���߼>߮ �T�            �v����1��!��ҕ��QYe��+������P ��+,�ذ�ꫬ�l�ǰ�7-�:��p_S�¢�ѹ��9*��}J�{u����R��HD��֧��_���            ��yK��0�IC��#%���>ߺ[�~�\O,Z�p�k��m�P�����׎
�Y��֡�5aFKG������s�m�s���υ9�7*#)Q9����rպOye��߽��%�����`���Z]��

���ϋ�� ]�ɪ���KG�r��޴��-�\�;M["auE�#-oC           h{�/^k/V���NMRfJ���
V����T�v�SaYE�=����x�ޡ�V��
����v��:!��BtX�e`f��-����[iꞒh/)~�=����V�ګ�pD���]���_f	h�3�`*�`�w�(�kt��О=�:�D��S�&��           ��)m�Wh/��Q!���i�����	�u��R��Қs!k]�~{�w��  q)��Ɠ�!t.��V)y         t|ȭFZZuq���9�|�p�U���h�}   >E_`Fܼ�         �SBn5�p��*����:�|�6��_᮳��p             ���Q!�V[��f���B}5RSS��g!�            �]Y���J9���o��su��&$$�s�}             �]W
�����D�              p�}              8�>              �`              B�              !�        �
Ҋ�h��E2d
�����Q����    t�         Z(P�G��},Chon�tԲ��b�4Uy    ��>        ��C}k	�u$W�RG-�p   �N�`        @3�s�}   }q1��*"n�"U��*LW��o���        4�>�!�׹�����_ZO��Hy���S\a L�ߢ ��D��̰�
#�r��A�        ���9��#bF��|��Sh=���3���8-  �3#�        �����p_�`����h�f0[[��j��..�}   �!�        �H���ᾎuͰLe��+��J�<Ʈ��C���nuK�6y��^�q�D���U�7i�*CUG�����7��=n��������n{g�   :#�}         �@�/���8~�2=a{�G�W�IB��=�g/���v����V�  �Y�        h ���e��F-[+	�   �#�         �A�/��	�   �3�         �@��� �    ��        �Ejq��N�&ܷ|��x|   �b����\t���         j�=o��N�
���� �[   �8>�Oeee
�Br"ӌ())���s��F"a�|	�9�>             �.;;[۷oWEE���
�����j��b�onn���}�pX����h�}@2M           tYYYY�
�Մ�ڊ��}��Z�>8�>��h�            �8���j*׵5���"�H���2���+�           @W����
����6�ա���\���bz�$A       ��!gh_�|�Py�-��~�>���r9Yΐt�|� y}���n�.��Q�   йuT��
�uD;ڎ<_B}�G�� �a���       �"�}*--V�>�� ܷ~S��*��t)���U�wz��>_��Y�!7z��A  ��h�[G�ܺ��������ria$U���       �ZUj�΂f���o.�޼]с�#�a���=���6lܦ��J  �����nN	�u��E���Q�7As�	�jy�       @|��}�
շw�Imy�Pߞ]�75ι}2��y}����K�  ����nk׮Uiiۼ&LH�{��t��E���S{co��\/bJ��d�(si_�@       @2̐vX��z���n�oǛ��g����۱so�|3��4��Ԧ�;��   iݺum2vNNN���[NRXX���׷��N<_ԏ`:���a9�       ��*�mڲOUU%�[RQ�3�6mޥ�F�JI��:B    �U�            :���V��$%z�
VTjWQ��hÐzF�M���3:fi�R����\�W�            �vrل��Sc�ˈ^ꖔp���e��!W�,X�w�li��V��k�����85����Qw�νzw�V=��+B:�5�F���V��}�	�1jP��CyUX3�{VND�            h'\>].+�W�@�_�b/�}�V?z�?��
78n�@���M�]����qO�e/��ؤ;�
�H�_6]nW�̅~�R�`S��ɩ�            �l��Z�=Oy�R�).���e��j�,���\<.Ǯ����Q�XV�o�/�����vU$�y�kі]*�)39����wZ� 'Y�W=�yP�\�2�߭c.l�_�Ź{�x�<IK���/-]'�"�            ���S�7n׮��Z�*��x�����������[�O6�s�����X�o��]�������Y�OԷ����5O�?���O��Y�ѹ���K�ɦG����>�����n���wcۏ/\)�"�            ������p�ԝ�.҄�������\g����c5�_u�e;�t��^R�"T�Ӵ�T�44��׻̅s̅���PK����=خ`i��Q��qU�:�>            �a^_�)�뛞R�>V��Og�����gީ3�ī�Wl�����-��G�����s��Y�            S�����j������@���;�8׹�ǀ檊<J�=Nvz�N��o���a=��9�>        �R����lp?ӌ�P��U������o�[   ]���c�K��պ��C�c�sWl<�>�ۥ�OE�v{_ ^M10��tG�����F�eT_Y��bS��Y� �        �
���U��obB�z�H�ˈ(^kŚ���7��V���%�  �+x��)cu�{{k~�^Z���}���[_�e�����x��s�Qʉ���Z�Z-z�����g�>�#+{�����ٮ-,K3u���t�.q��q��\'�'�&!�7	��8v�q��`���bvav�e�����F]i��y��[�U�9#�������>B+>��y~��>}w�6��E�0�/\�V��qx.�u�艭{5Ƽ�������&ko�k �        H0#�۾sbQ�!8Ы�V�l�gD}�w����a5��� �9G����{U���uK+TY�c����[��S
���񢼬��p$�W�r�V��s�G�VZ`�>�4}������-{a-Gυl�'62bs�\ˋrͷ�7�sɲ
���i�7u��=��:�>        ��l�wlܧ�1٨/n$�+ȓ-��  0_\������o�٠G��}Ґ)��9�ΝWiYA����rk�ޮmV$՚��~�r�\N�f��W�ެK��sU�X�bs��1��}�n�#o�r�g����W�{x�.G��S�}         	2ը/.��+L5�3���v�g	  `>�K��]���4��K��X�x�/?�{�#ύ���@7����z����������oVEN��ڿ�v�n���Θs�E�j~���[�΅�����a���ؚ��MS�o�D"�        H��Cut��nϙ�}CRu��WW�9ԭ��������FU]�)  ����F�#�1{]N-��2�$��k��u�Ϯ��N+������ь�C��܎�����֟��u�3?}N����fh�xzY![��2����r����hs��W���%y�΅��q�ry���ɛ5���ڡT@�        � ���/���!   �D��[q�A5u�i��=�a����-���W/�=��w_�v�����?,��=�eϘ뭚F�q�^.)3�_�ba,��Zq��p����������?p���O�ڡTA�            XH]G�����o5��ѥg��u������J}�mS�~����oEq� �;~.|96���VMtѾ��:�$�<7��'��U� �            ,�X]�X��83Me�*��:�]����\������=}#�9>��Tp�\(�J7�B�WC�������w��2���            ��1�!��:�}}wS@׬\h�{]�q��s�F΃C�R�1s�����a����mk��<�I
m�k �            ,�a��+��z�'\���}岳��9���Ԓ����W��ꄹ��D�x�2ez�����Nm�nP*!�            ,�U�����F�����5֫��_E~-/���\�in�~��>�z�����;$ ?��R�d>~Ϊ�󟽵SѨR
a            � ���ԋ�k�<�ugV�[�]>���M�F������M���.��&�������c�3^�f�xU���sT��rrr�bŊY���������$77wތw�s��ͻ'�-������sc�<��n��>        �Q����c�p��  @2|�����ۯ���Ɓ�vt�{ �H4���4ǎuK�uͪE�5^����/o�nخ;�Z����tY��썺���r�ټ�%���+�Շ�,5�7��?}��?����1�>�-��]������Ϋ�~v����>w����^��UcW�Ra        �(�*���ߩ�ހ0w�W�7m�~X
  0�ۥ�N_f��\ۤ�~�C�c^czw>��~��۴� [�,�0#�2��>r�p$��?����yPVfD}CCC��q23�d����٩d2��P(4����*q�d��۵���~����_���G�^9���o�P*"�        C��uZ��5�������Re�
   Y��65u����e�O��y�1������M;�mD���ӯu�?����<}�U斻�*g�Ό{���V��F�S�,+KT����i�b�Օ��/QQ_�Ub�^ߦ��\0��-8�\0�^�q�s�p���@_P��v�:�>        ��ػ��g�����  X�c[������f�(ï�t�����@oWS@]��I��X��ϟZ����涼%Y�r;�j��s�uNញ��/.33�|Ltܗ��1�!�q��[��Øbs�x炱"e�׾�TG�        0��E�  ��X!�`��<fZ(֛ՍJ5��uɈ���%+�K�J�qƟ�:6����J�         &��/��  ��DoG;�D�}Ɏ�⒵R!&��        `���R��o��V	H�H$���A�����^]��njVOc�zm�j8������b�x����x��z����QP���2e�>rO9E.�O  �%V������v���M�ʄ�#�.�>        �I �>�>$K4U0TOw�Z��Ss�v�Vہ2�6#�k6��v�ܱ���%��)�ࠢ�슪?vq�����c��.����5�˖���T;JV����  ��jQ_��M�l��x�q���        `�������000���.5TU�i��oޤ���p��i�)�i����&3���z��+�<?��k�F���H�#�C�ӎ�U�߽[�G�/-MK����_~�JO[��M  �
c�:+�\w<��3����x�^��K
��>        �) �3�+Y��ҕf���nGG����԰y����Nݍ�
G��8��s�͕��6��9��|�o��q��h���+�y��`hHU��������B�v�u:���خ ��[D%��$�        Lq�u�!Q�A_kS���nվ�Wo칱2_��%��a�����|�an�{d%>��x��E�u�o�ޮ?��6?��V_w���r�<��  @j"�        ���q�������`�s���jkmU�;��7O����\����6;w��i�~�7��F��t�̯��H����؟ahxX۞xB۟}F�������ew8  ��B�        0M{W�#�K�>$B�����YHUO>��}�d��T�����������.9�U�B�����6��G���Zw��U~��  @� �        �Fܗ�^/�"B����I�0�mw�������W����56���r:��G�ɵ���s�m9�.�4���+���J]������   �G�        0C:s�@z�`�������-��5�333����T
�t��!�ڴ��G�TU%�áB�׌�\
��g~�؟q85Ͻv�����w����'�]�@��a|�].�|w[���y�y�  �\E�        0
Z��n��
�q8�wť
z3��9�+h��^�W������z���J����o�˩��\�ϺI߱�큍(n0������F����u�ޫ�K/S*��>�`8��;  0��        LS~���n���/�j���e	��@ ����n٢��B�HD��Ҝ�^�o,Ɵ�X�ψ����b�y���V{m����'   k"�        �#� �K*[4��]��aZ�Ѩ�����ޮ�ohׯ-cm�R�G>�Cv�6#����1+;���WOjh ��>�9��>:  ����        `�������aD}��5��������v��������x�|��ph 6��ؠ�?�[���ʯ�1q  ���        LQ��q߲]�h��ˈ�0)MMM���V��^3�>�ݦB����v�1"E#V�H�g�7h����u_��   `�}         �D�g]�h�����Ң��N�nݪ�瞓�X����>�W�3�E#�Ǝ�^�?'[g��Q  ��         &!�e�*�������ѡ@ �Ϊ*�x��4?��8c�F�g���_�Bi�yZy��  @��        LQ_���V\�~����A577+�ե����ш�=>��I�g��g�=��Л�@K�(�   ��         &��/�q_���T���>#����A�pX;����U�v��_Q_��aW0UzTz��ԭ�z��~�   �<�}         � �K]�h��'0��P(���W��Z�N�2\.�4?��:���ޮ���;��M   H�>        �� �K}�}8Zww�zzz��Р�����nS�ۥ��V�����v��#j޸A�o����+   $a        �����>�-x����=V��q�#a��|r���Z}�r�>n�Mv�Co<��*[�F.�W   H<�>        �Q�jTN�7��㾝��R��柶�6�i�&u��+���>���;�;������Җ�׹w�%  f��[��f3��4�Ƌ�!�        EfW�����c�}�`7a�<
���ޮ���<�����r1Ϗc|>��q�X��_i�UW)��P  �4�ۭ���˃����H$�����_*���O#��>          s��Z_4U�
��v����ːlJ�E�嗿Ժ{�  ����L�����݌ȭ��oF�>���k�}��>          s��А����=֮_/�ͮ�C��n�@$��W_V��+-/O  ���n��m��=t萹����x1u�}          �@ px��M�4�ק|�KvV�;)��ci��۶�~���� `�X%v�����ȭ����%�6�>          sV$QWW���n���۔��Ǥ��4�������]rz< `�$;vKT�7�Ƌ��;V        ��\Z���[$�k���=�K�m��-_V�>�H�y2^XWOO��u��h��K�N���7!�W5��������� �lJV얬�m���C�        � i>��}��*Ζ�=��h��.���eu~�K��fOs�{c��CGL��Z_L��-
�3�ӏM���&GԦ=/�H� H�D�nɎ���x1q�}         	bӐ��:U<��͈��M�y�
�;�}���?15CCC���S$R�֭��mr����9m6�w�Tg���� `�%*v3V��B䖨����>        ��j�6�����׈��Rp�����^󱫶ƌ��\.�	���c��t�M��7kŕW
 �D0b���*����j��G�Р����L{��7����         ̌ݚ;UX�-�s���jj;hK��m�㭮�P{�Y�t�0�u��"Ѩ�نwJ�U�"��\��6�> @Buww���l�����B��b�vuui߾}�r���#�        H[tH5u��V__D�nr��	�6���={��就^�T��p$��w�U45�   �.�>          s�����ᰆ����ب4��mx���\v�RNy�  3��t(?�/�ˡ��!5u���'��T���4�K��߅ͱ����������|��9����gH���         ��c�}�����X�&�4�f���k��e�^�> ��;�\��E:��P+�r����zWpP��҃ol��U���N[�O��Z�-,U��5��p$�]M=�e��'v�T��0w��\�z�B�{��`q��Gm?\�ޭǷV�ۯ���ؽ���         ��
������G���o:�6��v54
 0=���ձ����l�ϣV/1�ǶT�yA�'Yq��v����յ���������|��܅k��<�w�[$��y���9����˩���Jݶ�r���f�/?[;{�>��g�������         �s��lm�-��N�7F��};j� �{[;������<�mC˳3tђ2-��2�1%���O��>�����D}��2W7���6W@;��@����܎�,v�'�I������7(�
��vj[}�Zc��$s�h ?=�\0���y�n>}��<�m�~�c���y���wq�>w��J��U���G>�a]�iwS@VE�         `Ή�����"��.�0���X����  �s�C��������7���
f_��,���/0��zF�x}ۨ���}J��o�ן|Mߋ]{��ߪ'�����|�r������ɘ�?0�\0~��+����{d.�����w��`�	�޴f�H�7��?~F��8p�5���-��ǯ���.6W����t�>&�"�         0�����6�ld}3��,vv 0=Ɩ�'�D��/o�Y�郫G{ם�x԰��F�7�4���Uɾ��z}��k��W�ޏ����֓�c����̅��#�-���K֎�w���>����==�Mz�J��u��R]Vy�^����         �S"�����k1C��|l�;#l6��CC��>�6>� 0��yp$�+�N�������-��Oz���Ս�g�H��88�������̊���n�>�zC������לg>7��%�         ��G}�cxpP6�L��>��`P��4 f�p82r��������ng�ڣ_7�& UG���'��0/k�뻽@]'���+�]�j��w=���        $�@(���~�d�2M�9ށ�3b,6N�t����'����rv�C�>c^?4"����j��w�[G���b7nui�I�gl;�Ɓ��G��m8q.dx�#����q�g�qyi>�fe���GVC�        �]���]�&t���WI��
E�~��ϛ�����x#�"�b_�H�gg��al�k�ICA f�Qa����J�ym{��ܶw�k��q@�o���I�[X���D�޾���
3����_`��#���o�:c%�/\�V��qx.�u�艭'΅�����t�[���y�y��(��         �#��;'���آ���&;��@��[E܇)�ي�v$��Xr&���o ��# �̸f�B�d���9~�ʲӵni�*s̷մw�#�J���Q��x�]?|Z���T����|�z~W�^�ScFP�=�h�c�4W&���V�5�	����B�����P�屯_�����G�������}�\h���c�YQt��L����         �&���)eLu�G�}4Y���
}v�K�Y�hT.�W ����ukuɲ����g7葷w���m�k����33���������hÑ�~��{���ێپ��/��¥S�-=���ڡe��؏��R���y�k]�>�S�y[�V�K�>        ��j�����
�;^#�kl���0_�d�l�k���v�ugN$*���\� �cu����"s�yi��}��,��ҥ�N�)�������xy��nj�ޖv�#��
4��\0V����s.����/v��kW��W�j��P�1��0�w�x$ ���� �}         	p��M��ɖ=�����]�����
�w��x�v����/���):l��B�7]v��������� 0S���o�<�������L]�j���^�׭?��:�4_��3檩��������.3��А���v����܊4#v�����y��0/K�p�:]Vy��}�P8,�*�-�]G��m.|��s��$o̹��7��sV�[O�y\z�o�w�o5���iIA�� 6��Cgp������+�;.        ����5��b����t:5<<,_N���n�A(L�=�9udd 0sz��b8���z��`�ܰ]O}�f3����%���5����Nx����[�].��fnYz�wמ��c�1"������N׮Zdn���?_���XE���q��s��o��_�{��s���`�xF���<�G?�a--Ȗ���W/?�<��ﯾ�U%y�b����gE�}          ���c�}��"u�es8ee�i��lJ+- `�նw닏��g�x����.=s԰�/�;ߌ��������а�}�ym��O)��1��xm���`eu=�̅/����^ߪ��<�֩������K�4W�,���z}g��酷�m{���w����E!��         ���v����'a����#{f���05���s(R�) H�7ԛ�]qf�ʲ3T;u���nl7����#ϟ�q��3V%{iO�n9�Rn�C떖��w�����BiV�9��o4=!��o7��ߨe9��n�Ü;����m|���*�r��Ñ��j��         �s������WxxXQ�K �*�ק��N���	 �8���F�d����n�|���4��j}��e�=㯾w��d�������������s����<�w�29�v�����c�Ķ�>          s���5}�����.�0U�K�pDy
 �F�g���=6P�9�٤�[�'��Ҽ#�=����0��������󟽵KVE�         `�1�>��.ON�<�����'L��aW�nS��e $�u�+��1ύmD[z��y��@�#�8ֻhI�I��5�߽���{�;����B}l.Lduʱ\��B7�^b�s��o�         @�Q���S__��Pw�ex�&�X�/<4���r8�3 L�mk+���uOzݙE��m��<h�.skѣEboxaW�>r�
��7�=O��ShH�����$+�<o��צ�FY]nn��/_>+�NK�k�B�Dc�<��xo=�R/�Q�d����'̅8c�ަ�uK���O\o�pi�Ư׏��e2�]        �(��es�ͦAO�0?��~3��Y�XM[ޑ��D �,of��:;Tv�U L��.<]߾�
�vW��8P���3,2"���43L2�kV-��H}���]�z��Q�w�˛u�����N-���_�C����z��ּ��a���"}q�����W]���6h(�����*;;�<fKOO�:;;e��,99�1[������%+��E����Bϛs�A���΅���k~,�����7���{�z��u9�(?K׮Z��W,��~�y��l����}         �h*])�PP9�ղ����Ws�Z3���������Ve-^�h8�a�K�<�ߧ��FU�]+ ����.�|�2����&�����\�ows���ȋ���\i�}+����O\o�60���8�}��-��;deF�
��Jj���o]]ɍ�5���,�m�3s�No��\x��Y���ǜqk�
�c,�?�lܮ?y��1W��
�>        �1�,8�|$��������؊����˖���S~�B����8c���PH��B�-\( ��<��m�V�..S~�o��ީk�7���mکp���ѣ���{�m���胫��s$�;>��x��\��X-����eff��Ɋ�=^�Č��Mͱ�pAl.�3~�q�~�iǸs����+��UQ���׆#���^��ŷ���c* �        8	3�J9m�}���o�2~Xo��W|�Y���c*����&̗����v-��f ��-U�a|[�07�������{�32C��Mu'uߝ�}��ϙ1ߪ�|U�d(��Q_hH���ޭoUG����Ot����o���h�o�2����=��<�m|�f�4;C������+v�T�G#�        G��#+���$���-++��r��P46�vٝNE�����9ry�����%_, ��1VL;�2��dl�k�pf�&Y�[����'j�Z+�א��fc.�b�ԨTF�        0�}���.�Kiii2~�[r��jݽKr��ߒz�C���檿�G9kNWZ^�  �-===J��ܦ�0�q_���8��}a        ����>���端�Oe]�����Pq���"�0:��._V�����e_��  �-V���f;�J���
1q�}         �@ܗ��p4��o��k�T]����mfվ��s���١��J-_!  f�բ��x�7���x1=�}         �D�gmD}��j_mm�*.�T��ܯPQ��^���c9���r�g�.]rϽ `6��Y1r�s�=3z��6^La        �����i�!��>�%--�<�眣ƽ����H=�5±2KJ��P�U*9�T 0[�Ѩ��6^La        ��,<�|$��>����X�«�Ѧ��Sw$*_v�:;�ü��rx����֍��   9�         ������0n�[���
Zr�u���ߨr�29�Aj��;��,-U}M�N��6e	   �A�        0M�}�Eԇ����WOO�
�X��͛��PyY�����D4o��ݕSQ���}>�~�M  @��        � #�k,]%E�q��K�������*//Wuu�V~�N�����t������ؠ�*��P��|:p࠮������   ���         ����xTPP��HD+���v���/�TZ^��m�o|YY�ث��t�g>��E�  ��"�        ���QN[5[�&A͢�Ԟ{������U0��.Uم�Ж-Z�p�|�C
vui��dd(��\��)�̳��+  ��#�        �&���Zp�m��URR���a-��J���u��N���*�h��Gs���WvE�Z[[���%_��   `�}         �@�gf���=�������Puu���x�v��'�ki�)ee�76���<��f���ѩ���������   ���        `����eA�;�#q&#����h�G?�w����j~v�S}���_v��J���ݭ�`P����'-M   ��>        �) �&�>L����U[[�5���v=���[URX���k=��R4�� ��P��jkoW��n������   ���        `������S�t:͸���N��[{Lu*-)U�߯�C��������+�NOWCK�B���Ͽ!wll   ��>        �I0�1�>�#��Tķ�mhh��;>���U�Ν*,-U���ml�@w�R�'=]Yee�é}�5�\V����9\.  ���         &Ȍ�Z��Rq��������.��T`�"��i���L��u76(<4$��;��(*�/;G���:x`�N��6�vÇ   k#�        � ���Dܗ�2_��y^Z����l�܈�REnn��~�\.�ҊK���G4��{{�r�-UK��mR4*ˉ�{*-��O/,T�fW}[@]A]���P�eJ5�pX�`�<_���sw_j����KϾ-  ����        `D}���/����G>Wl�8���cI�׫E��5=]�{>��M�T����+,Tn^�
cGG��E�a%]��Q��,���r�s0�C�Zx��ꮻ������GJ�ît��-�3<l%  ���         A����>L���`QQ���������b�>��j��]X�̜\��?P��3)[�[�������]����ɗ����ꯕSQ!   ��>        �1��-�}��ǣ(''G��jۻWu�����VeŞg��)��HC��f�7��3����y32��ʖ;-MQ��;RC]�\YY:�>���+   �&�>        �Q7�"ꛃ�nQ0=WAo������4���._����{����)=7Wi~��KJ�YZ�ၠB}}���~E#�)\��nn�kD|�����ͭw"a5����-���b���{Uq�  D��w�l3�;`��[`���C�        0
�@?ؚ��Qy��0m�QRR��իh�W��ղ�B!����u��-r3���]�ᐆcG��p�F�#�/ˈ��)��v�v��9b��4�[v�;�Q��]6�=Tgg����)?����{��h�  H���q�EbO������Ra�~�d!�}          0E������
~K����պo��v������������������n����m��ُ��X�'j�D�
��B���HD����ѫ��~���py�N=�,����\� �TTVV���z��n�pX��}3��:^#����3�>Xa          L���Mzz�yk�y穿�_�]]�ؿ_���iiQo{�B��2�>#ȳ��
}�j}F�g��g�p�ض7�*-/W���/����t�jy3Xq 0wX-v�G}��j�G}��>          �aN�S����QZQ{˥�F�V$�P_�B��B�}
���t���ʝ�.��k|�� ����v�g��СC
�BJ&�{�>�"�         �0V�s�\湱�/  x_��DE}q���I��G}��u�        $�������r�Ӿמ}mz��2c��b�u��x��+   �mɊ���%+�#�K�}         	�����ݭ��yܶ)�g��.X�,c�]30�}����#  �|��mj���%:�#�K�}         	bװ�:��Q_��)v�[xNw�F�זB�  ��HT��/n��C�        �@F���ԩ�ly\����D}�e��}?�  �|d�nUUU���{�^�*f{��G�Pb�8���        $�MCjj�TAa��N�����u�d�7��V�v���Y   �ߺ���w��Y�weee�{S�����K��훕{[q�89�>        �$0b�ں�����
��/�T7��    �a            0��y\*�HS�`H-=���+��E�            X�-gT�˗�9�|SM���W'��^�S_�d��<k��d���g �߼�_�z�m�nn�
n>}��r�Y#�7�6�k�|u��s9�ZQ����򵦬P�K��q��m�o�W~�Ra            �d�>��-�*��y[{����wa^��􇴼(���2�n�y�J�tF�����zx�.V�yi���uL`.��S�U+��p��z���R	a            �d�t�%�D}������|X��9���ޠܰ]U����{t���`q��N����+��ݧW�jX�?����Q�D--�3�KE�}            @]�bs^�/����k�O�}���G����.}�;����w��￱]������uN�]��z����O
�X�u��p�炡��[�ַƎmoh3W���^�TD�            $I�׭��2��XI�M�&3e�<���G��/�����]��BgV���~윕����X�9n��<uo�~���I�}�~��
�)��i�}            @�����T����А��c/kq~������s��kh�����H4��ߪ���5�scE4�>X�1J���8﫱�� 7sR�|ԗ��            �$X��\�8w�y���m4��\طp��ٝOz�owU����f��˔��+8(�
.Z��\0V�4���l�7��        $�`(���.�jN0����/  ��+����W�f�6�6�{�o��=V獜����_UK�V��a�ie�}7l�l�\��헛s����)ͅ���         	�{��vM�Z�7]E���&�Y�d�����8?��  0����|-��R(֗���v�A--xu��@׸�c�h�}��Ź�}��o\{��R�p$bnG=ٹ0W�        $XW��}��"7Cp�W�-�f�nK�rMv��^5�*�cF  ���uJ���������������v��v�<o0��G�Q�e�	H�3+��ך����fmoh#�        H��Fnq���jlё�O)c��5b�x�gK��  ���p�?��������6M�>i�c������z��t�K@29�v}��͹��u�sa�"�        H��ި���=����}Ņ�J�o|�¢/  �D��gkeq�"Ѩ��ȋO�>��V�3�.5�1��a����L_���)+0��=�Ҕ��\E�        � յ�
�{$[���3��v��fr�S`�   QY���^~�y�߿Wo�4N�^��"(c�3��fR'��G���_��-�\�_G������`�p,�>        ����5��b��  `<F|��;����P]G��{��iݯ?4t�s�G��7���T�wpH@2��R����Nc.lND�            ̲O~`��>��<���/�o�a����:���W��Wm{�Iߧ �7r��?  >yީ:oa�y���^�}-���            �lI~��h��?w];�uGo�{�rU��y�|(Ѳ�z`�5#�tki����gg���Ů��ji�Gυ&8.:j.���ң��\E�            $��&e�<��小\k�}�3�xط��@o��^��~���<���LS�F�:�            �l{c��ܶw��
3��`q�y���?녍�͎���:]�b���������c�����]������z$�{���sa            0�~�y�y���S��=�c������<;���8��q��6��\�Přij���ڏ��j�|"Q0[&:.]V�'?�y�c��0�            )���GOl۫[Ϩ4�*��M��?yF�/hv��R�y�J�+8�~��RANN��/_>+�NK�k``@V2����}Ra        �(�3��Q/�-Q�M��  ���]�|��|}x�R�������QU-���u�����_����[+hMOO���l���VWW�����W����1[���bc��\���@�>��c޶� {�|I��[�]~���
������"�>        �Q�����v�07Q��ʋ�	  `�8��'~�����w�t㚥�1��i�s��R_*��gD}CCC��q233�Q��ɍ���/
�����ʊ��f��q�-��ԧ�[=���V�ǿ��)@�        �jZ���}�/����	  `�ymo�.�ׇ��7�3W�3V�;:���֩o��y{��.QQ_\FF�����/QQ_�3ƾ;6W�        �q_���Z�N�i���  �Ly��V�_����ψ�>���T���i�*�LSWpP5�]��P*Ht�g�}Ѩ��]�ƛ�yx�d�T8�W��Mj.�z��)��"�        q_�2����ߟ-  ����7���j�j�����^�.qq_����dŌ�8�>        �	 �K=D}   �!��юň�l��ߖ7�Q_\�cFLa        ����>  ��`��/�X��0[q_�W&<q�u�        L��E�QUԽ+XQ  @j�Z���f�U�_��B�        0Im�K�G�>�!�  HF�f����v{f�~�m��>�>        �) �ͦ�D}   )�X	{>�o����        Lq�u�Q������    �:�>        �i �K>�>    sa        �4q�-QY�Nc-!q���*�)H�   `!�        ��E����p:���P(��v�]6�M�����9����y   FG�         �r����Pn��x���E���������#g,�����<3���H$���&  `t�}          f�{��Y�no�l��I���O^�L�{��������N%�5�+t�ى���w�58��U���,�eM���}Ca}��w&�~v�M�?{wW��}�N�h���]��+u�EZl�XX��wم?�-���,�Z�-5���K�j���)�62!�ə���:Wf&Ϝ3g�<gR�7���u=����j�   �D�         @����1p��ڭ�P����vᚸB�����v��K\��Z�T�.5-M�F�	   �F�              !�             ���             �B�             `!�              ��}              X�>              ,�`              B�              !�             ���            �r���bUf)H�m�?�             ��������KBB�XQjj��,X`���������D�"��}             \�Z�jr��9˅�4�S��>U�zu9{����}ꋉ�6�>X�>             �B�}V
��C}�b�p�=��!�            ��X%���P�]q�_�1�             ����:�V�����"������`            �BWXa�ª\WX�K��=�         `9~>>�����������c�O�n/�׷@��7U  Ȓ��n�r+n���            `�
����Z"���%��^�         ���a�$�7���.DŊ�\������JHp����%&1)��)�u  �6�9rD��✲~ILL��V��=z���/rG�         ���5�Wq7?�9n��l��5 ��DFF���34l�PJ�����𐈈			q�������>              ,�`            Pxx�T�`?�ML�KQ���"@q��]B*����(m����            ,`t���x�6�׷�� ��^��}j�+%��֑A��J��%��'�wI)����E���L�z����(�\x"�\�v��<=kU��}Kxɸ6���m�ҨR	���4�JL��<rF�\�[6��#�            ��A�֨^R6�/�����9����eL������S�תl������~X$�®
`e��7̅k�̅2�����r%��|� �g�w�?箑Դ4�*�}            @!�ψ���L��\2�r\R�l9*{�]��ѱ�i��դg��Eo���dᣣe�G?��K���?2�4�w ���,�m� ,*�T�U&Hz6�!UJ��0�[KINI����"�            �!���Ȗ�埶���6v��G.^�/��JT|�M��\���p�)�o*��?���d� V4�Y]ӆW�e.D%$��oʆ�粭����%/�*���2���Z�ܰWN^�+"�            �R�����^��#�eZ�L��R_�*9u�x����/�ˣ��u��װb�D��;�{��+msa궃υ��$Y��X�cSR���H�ZU�m�J���!�Ԗ���+"�            �W�u���%%61I��y��+_���
���8�bv��iR���ުzE�}��W�f�uʕ*�mhv��&ا��
�"�            ��jȄ����Wm��W#��ˋs�����@_��G��rw��s��ś�m.8#اRR/qy1:V��`            �b>����>��!����|�sہ�)�{H*,ʺa&?��%���}���g�v9u{���N����e�*�}            ��=?���.WJSR����3U+h�jVN����&[N��*���T�ӹ����o/OyaP�\������EYrV��`            �B��ح�����mr���mK���4�k��y{B�Rt� Vжf%�����p �`��Ȗ�����\!�_���~�kIu�O�����f�	�Z�>            �E|����q}���C]�b�L��h��ҵ^5s9<.A���N +й�Ѹ~��B�UywE�ͅ�$+����s�Q��2oo�$�����            \䩾�I�r�R��3�����ҿq-yyH7sY�M��TΆG	`��ӗKB��悝V�{cDO� ���%.�G�            p��Uʙ0��l�n�z�ӶթNU�����z~�ZY|�� V��>�\�|��r*�@�������������-�+�����ɽ���ּ��!�l�==k�X�>            ��<=<�1}L��3ע�����������K������/���;��j;j�\xeц�FT|b�emA-kC��w���܉�L���.-d��y{BĊ�            Nv��&p���y��$$9e;mkV������C}o/�*��&�U�۱���Y�\��L�ͅ��"���Z�?�\�g�}            @qU�\i�3-M�	����~�{��r��rRJ�4x��ѢZ���	��1�?Z�C^Y�ʀ�Q�|)�S�=`���s�[���l��s�9�����O�^�ҦF%S901%E��`            �""��}��#�X"�a�2������n�<?� V�G�Brj��GBr�D'$J� ?�X�[&��            �����e��� ]�V3�/F�ʆ����-o��-xd����j�^�n��}�W�6��#�2f#�Ċ�            N6m�A��wÚ2���a�}����8�n��2oҨ�P���٫$��'�i��Ԑ9G�������]��r�6;φI�E'�>            �U/$s!��K��S��ǧ/�lP)�ʔ)#�5rʺK����x��4�kV�l�b����Md���ML�q\�Ƶ�_���_��@����            �Д��JͲ��r|r�$���;�{�z�5!ge֮#be���&ا��DFFHDD�XALLL��߂������zȢ'd�P9s-J��D�U+h¯�ז����g������bU�             7T��_�e�^rw�f�OC�V�i�/11���	.%.�ɕ�+�!����R��W�h��,�Yv����"II�nuK�}             ,�U!7����+�������E-����rk��ҹn5)����m<qN�ܰW��>*VG�            ���GNK�?phl�W�����!7��
����K�o��3υo6�3�����)WJ*H�����#Q�r!2F\�"��I�.�            (TQQQ��Tx�+����.�VX�>;�]oC|M��Tۋx�r�Y��>             ���C}v��dg��

2?�Z��� �            �PX%�f��p����p�u�            �rڎ�J!7;{���Yu5ܗ�}�a)�             ��ܬr����+а[q�_��>             .U�Bdi��G�              ��}              X�>              ,�`              B�              !�             ���             �B�             `!�              ��}              X�>              ,�`              B�              !�      �J�-)q�*	  {��>     `G�      NU��Y        �!�             ���             �B�            @iii���!�Eq�_w@�@�Wc�\	�L�O\R���<F           �/������D����T	(Y`��������%�g� y1�O��2���'�c���$2,L           ((իW��g�Z.즡�����)��oJJ������"�(.^�(+V$��h�/,,LRSS       �?��-�Z5th�C'��K��=����ڛ۞��V&o=p�ؒ�޲�����w		������,   ��ja7{��Y����P��`�b�p_��      ��u��UYu�t�ۆ4�'I))����L��;������������&wwh�e�oD�R9����#   ��*a7mG����U��P���P��s�>       (x���m��μ:I����}?,��뎝����K�r��ĕ�L���ߎ3aR�|i  pG�vsuȭ��/�`�b�p_��      ����uD:Ԫ,��m,o,ݜ~���:֮*O�^)/�"   �n�r+n���!��X�p_�r����Cp�+W�HZZ�        �#2>Q8a�}�Y�Y��w|�����"3w!�  ܞ��n�r+n���Pl%''�����f��       ���m?$#Z6����擡���!��i$���  (
\v�Jȭ��/C�         p�:%�bM�>��mTS����[�  @Q�a�#G�Hll�S����'		�b��____IL� �`         �&�SSe��rG���kd|��r>"Zք�  ��&22R�=�u7l�PJ��+��������ۊ����         ��O�ʤn-��vMdP�����풒�&    ��}  ��\�O����O��[����       @Q���E9vU^����xyɔm   @�B� �0?O�,?O�?@     �"�rpI�]6Xj�	�r��R��.~R6�OJxyJ���xzx���rBr��OLB�$��J�����X	�������Q��������"(l���*[JV,#��Z�@�`�YU�c�ϻ����2��v�]$">A�c�ψ��O]��c���m9s-ʴ�-ʦo?$/�"뎝��W"  �[5��{�I����yf��?�>��{G�&���?.�Y�E �e�Od��N_��g���>��3���`������Z�>        ��JAҪzEiV��4�Z^�V.'�˗N[$c��)�î��K���e�t�	j��i��i��ҾVes,�b;��g��O�oKã���H?�b[v�	���d)*>\�C�޸ׄd�?%}��OÚR�t�\����OIx\B�c==E���\z֯)�)�2s�QYr�D��֊�=T�zʘu�>zFB#����AK�R�cKd|b��5`ݫA)�gB�������JK׺����K���$�O�JjZ�m��լ,�kT4��7�8//\�vl	ۓӽ~uiT��D&$ʚ�g�lx���<�|��_�����+�����t�r��[���SB��^���帯-�U4�4�z���';Z�V��y?�IL�5!g�cʎ����,,Wc�l�zZ��~f�����ۨ�m����o�m_c��_�L���_C�lϩV�\w�\��f=�v�]E�<=d��0�a;?洯�tlf��D۹u֮#�8�c^���z��ڶ�_���ٙ�s 3���F�4�<����x}l�?/����}����ӹ��s�s�q���ȶ8��)H�        @&<�ݠ�t�SE:֩j�����蒑a6�5!�UG�ȡ�%�=�z֯!=\_*d�`Ι�ҟ�8Ҽ��MC.{�]�-�BeM�YYq��[�4��S
�j;>���|xl��(��_'�nڗi���f?<R}��oצ�	���'Sy���_���j��n��.�-�tS�lL���Q����o�mZ��ٹkd��5(���婾�Lx����Hyx�s��H�e���}g�&�v��^��X$'n���ᬯl��k�j�n��'D�<�כ-�U��&4;�s���%/.�pS�,/ϻ�j=����݅�yd�2��ȷ��	�h�3��j�E���k��k`����]FK��IS�������I�*��o��R����������ג���3ϩ��{^Y�ф�n�`��Ґ�&�hw):N����T��H�3_�M��҄���]�?��X��f[����nV7��zN|h�b	���i;�'�0x�Ƶid��>�n^��^���<ҽ���j�p��2c�a�8u�䐫����)Ȕz�p\_�|p��F���\�}�b��=Q9|��
�       P�i�K�j2�I�ߤ�i�j5Z�jd�fQ�zt����x�q�p�<�{-D�tcZ72�U^�e8�`��.��4����e��7T\i�c�C5.��5g�Q9�{�ʅ�����}��߻���Vg�N��)\�aSmז1�4��ޘ>&|���C�6e�����VK[��]��/�o�y0�7U���?ݯ�	�i��n��ܫ᲌A4�A�On�oBo��K���~��[;��X4L;Ӷ]�qc�a.��3#��:o�(��Δ������<<BW.w���Z�7�i���?(���;q��2��ι?�lc{~=�sפߞ��]iɗ�v���k2�O�d��3d癋鷿o[GƖ�vZqvޤ���ݩ����c���y�F��^���ͬ_+*�`;��|�ό�u�@��
��<�vwN�h�����ۺK�m�~�ao����75��i(��{�m��6��^�C����z��}�����
�������ߨG���Ǎ����/���=G7����u�c��혷T��|�G���ꫬa��1�י+o���.�ʗ6aQ��qI��P|lZ'�\�����6�����ЩNUs����	��@炶�U���?����N$�       @1�ّ���ʨVdx�7��N[�i�C�h5{�Q�������Ӏ���eL�FYd�H��h�J�wF]�\6c�a���Pz��U&M[���5Е1ԕ�GZ&��m�k�{H�A3?�ӯ�BQ��vS�,#���y���QV�>�
�s�V��`�s�:�����>mM�7{���ۺ��ӛ�=��,�w̄3�z�S}�g�n������2�ۅ�z�ZU���i0����߂��th�e��N�y��M����C}=ܵ�|�n�yT^�� oyn`�l�j��!��Og��Z90�P���ğ��V^X��\�rN�,�n��v^8l���w��/'�o&�[�K�^�*���|����� .2��ޥ-�u��ώ�:_��2�5<�@�[�����'�u=L7�y�,C}v���}�f������e��N��'m��;+����L��Iuo����/�{����wܚ���p�K���v��`�{ƻ�{��ZE3��>��ߠ����[�v���t.��a.L+���;#�       @1��k+�{;5��2ѝi���:57��X����� �Ɩ�(xZF�����	��+N٫��8��,9pR~ܲ_~=|*�R܃�>��֛n�0�GȀg��l�L,'�~��L���U%�m�l� =�ׯQ��j�K��i`L[��v>�J|�*�5U��֭�k[ž���q�A�>�jJn��ڃ}}ג��������2^C|��V��y}�;֮�c@R��û�	��m��c�}���9����N��~}�u���P��#s��_jU6����[��65*���+1q����f������rv�������>7#Z60��ֶ���1��U+0iX�Z� Y���ڳk���Q����~���'����	k�Jm�]����ZU+������_+C����:��T�m.��6���`        �@�*���mLK#�\>|wg�yap����睇��;���+���ǏG������ܣ:_^h�J���h5�)��������uiհ�n���5�φ}:K�|s���*˩�]I��c5k�����|��@����ݔ_��1k[�`���>Ƒ�C�C�����L�x,��6���<�k^�������d{L��2��}p�������q��+���1�T�1���U;�瀎7��2��A]L�&{{h���^�����^Z��T8�O�O��c�>=k%s	n�[��rw����/�m.�        E����k�v�����"C�g��7���5��O�����ڐ��?N�S���Ǔ��-t?����{�6U��[�]�]m-جJ9S�e��0�MLJ��V3��K[���� ݹ�(���?.�jwG.^3�/��JM��?X�t-�~zY[����ū���k�����cxP+Gڏ���SNN]�0�>u�R��fX�^�K��L�m���>'�������������;<�H�1�:�ڤ���^
7�r�u�'�b�s��Ǉ8pn�NH���ѿ=���>����k*E���o����8b�����fus��Am�<wOH�۵m�V,<s-ʄ��@χ��k�N�v��|�aO�֧sD[���N����p:>�a.�/�ʭ�/��+񶿋2���.�       P5�R^���޴�+�L[�Ƶ̲�d������y����6����L;��HWZ=DâK���~�"�O�	\G[�j�ap�@�~8�֯[录�LL?�͍��ݳ�Q2u�A�S�[����I9�[�����-���Xm����ӯ�i�m|���]��ǯ����e��#rG�&َ��7$=ȴ��S��I�rَ�fӾ��sv�ȋ�����َ߸7�������=�0�~0�ϝ��kN���W#e��S��������T�tȡ�w��Ij������Wc��`Kv2��[��n�Lտ�$�����v���B9;�be�o-�5����W�l�o8~.=Lg��#�M���L�zЄ@ղC���T5��a��@����i�m�T�C}.�>Y�K���V�^|�}�Χ�ån��َ� �V۱�s����2�%�T���5���R�B�c���Jd�����l���������ܑo��ΟH�{�_g��]<?������;Ԍo��u�����$$�f������4��b�o_��2�}        !ڪH�t��~�������Y�����h�
�*Ȟ?�[5��cX�8�@���u��������u&��
����F�d���5��	���p�iז�@7,*�\���>mkVʲ�������ӯ�o�Nޢ�tʦ�ݧkv�����~�~�	�eU�L[">4e�	���c�ZiU��4�"�r)\���*������D�M�e�MO�ޙ~]��M��T��gp�����v����V�yu�F6��~����+2��~�r�TW��ō4�������<�j��e�s��,+�j0�e[2m��)Ke�}C�/���_oܛ�z����F^���L}����&S�Y��H/۾�ӱ�M��J���z�ٽ�d�t����r#m��ȴe�n{|�rY��S��F;΄�ˋ6�_�����X~~pxzK܌���O�`jkϧf������)Ȩ�H�C{�]J��S�q1�E�l�y=�w���~}��se�3�|��X��<��4�Z�2�֊'._��ڢt�C�3�\<�Imi��8���O�J��jW��	�w�o�C�H~��'�/�<g{_an�]�����>��o.���'����u�[���}T�@`e�        (�u�_z��'���^��ipch�z��V����L�5�PF��Sz�P9���c�����ƽ�RǑ�L��2��t��lc��i +��nӶ����:}�}<Ӝ;ǵi$5�˅�h������l�	�e4��奡]M�� _S��rT���p}�
vJp�[(ui!�vj.�msJ}�:)�/�l��e�����y�o;�Ӗ�ڶvΞ��[L奌��^��N���Ѵ��v��.]�������Tڎ�����[;H��5���>���%�d�.V���˷���s���t�کV��|2���{h�Yw�yn�qtB�m_O��}�1����]���ݩ���w�!��JT✲������T�~]�^�ڞ�i�L���e�n7���|i�����}�ʒf�����AV-����r�\؏K��<rZ�c������Β�l���H�r����}�m��Y.Egn'��y����3�;�m�ԓJA%M[��;�{+��0_F�8t��m�ڷQMX8t�|�a��`�i7;����}�_{�T��	�i��wWn3�׍��qpy�k�ߏy�c��?n=�i�I��l�ڷ��=��}��R���7�B/�}?,���/��dG�Ǻc�L���1}��2�aϗmsR�?���q�Ѹ�A[}�zwŶ|�/��G���\���[���υ~f.��h~���?}�����1�2_�{����n5D?�Q2�3MEY�"�       ���𕶨̪���a��:57�M���V~�yD ��c*�=Ե�i���y{yʤn-MU���;��A�i7'�A�V��p�ylگ��1��x�iu��~Y��6m�U�tqĿ�7�#4Ԥ�1]��(/���,��؟��*��{����v���<iGh���∼>�aQ��Y+��}����qԪ�g����L�1̙hHPGh��g�6�#�^�&N^,��0��/�:<�E�����Ǥ�N�>�9�qR�Өf�!\/>��2ӊ�u���V�f;?h(�ޢp���Ti����syB>[��v[�R*�̡'f�����RC����<�sA+�.>p���t#���vMM�y���?Pڿ�C���,�        pSZ���a����h��i��/�4��3��6�ŕV	{mx� �=�>�k��۱�L��4S�R�_V!�U�~�j�I+�i�a��3�z5(5m�!yc�f*+o*�6U�&thjZJkv������&��*�.��X&�ׄ
wѴJ9�k����g�v˦��k�U�Ʒoj.�{ɦ�*�V��>�����)���_m؛����F+�j��9�4A��e�e\���v+"�       �j[���.P�\)A��lPC6=3A^�e�|�nW��rR��W��Sno�X�?]�U�oZ<�ɱ�e�NÑ��T5�S��^�}�/��N�r�*���3�rφG�ĩKm��*��� ��6��Z�^^�e��𗘄DS�0�Ј�\ף!�k�	��5����������:$`%Z5���ZL�^]�1_���.a*w�|4��5�pz��p\�����"Ǫ���!geƎCrG�&�����	�       ����&vk%��f>�F��F�-S�F�L{��1R��k\K>�״nC�� �~`߫A��̕r-6^�==��l;����yݱ���r>"Z~�q�T#ʎw����w�� k� �V��ʞs����p��C;�y{���ὧc3�N^��JC�m�//.\o����߹yz�'^!1	��>ݯ��)WJ�RR�i�$95U w����լl.�uf��B^���=�״Jy�*�}        �	���mc�7�%p��{�.yx�Yq�E��>����m��#Z6�v�*˟~X\ mŊ�wF���8�V���d�i�;u�Aڼ�lZ�q
zf�j�pEP�m�?1c��~x���t#࿰`�����v��{m�;�[KiV����l�'XB�r׃����Մ�َ��v�n{O<��DsY|^�����|�J����|2|!hl�F2��z��k������Z���+��\��f'�\�a.$��B�s!��³]� ?�*�}        ���n��C�Q���+�/3!��./�������������KNW�t�	��e�r���� ��*Ȅ�هK�J�#�[ɛ˶���-��������4�Si5��m�_� E��c�d�'��͑=�U���6}O^z�<=k�	�i��go��:4rwǦ��FZ��:�
wi_��ju[�X�eEۚ:�>�^fQq��p�?:��.��~��m�	�       `q��������}p�����m�Y��2q��ZZ�j��wG�6m�������U�/-o,�$E(#�o��6�,�1uL�O�������R1��i�I�c�xЪ�Z��Z� ��/��Ff���n����wVF�lH���7����}4�q��K�j��ŨX�p����r�[O]�\�J��e��M�J�Ρ�g���K�q�}�W
t.�U��U�/��P��j�W        6�E}����U5�z��x�w��_͓CaW��َ�7F���:5�����޿�ԯPZ��L�SZ�%��ge2�SR�$4"Z ?�£�r�*�s�o�ҹ�\aڶ�f�M�5e����L�B/�}?,�r�'kv�'lw|���������!g����09:z5�!s&�4���0�"��Ǵj�[u�X�>        ,������Q���Ñ:p�Ze�eɟ�ʽ��"��Z����h��)����*

��VM{�1_Ε��D)�_	�u̱� 9q$�{>�@0�ʖ-+�5rʺK���xkU .n�[�F���^~��D�%d;�|��|=aPz(\�p����bU�        ��{;6�wF�2}֡��~h��}�j�j�^qͫ����&UKQ��*���L�q4��}s���KC���)��a�u?h`���wɱ��G������ҥK��yۈ���ܿl�
���R�L�8Kdd�DD�/N��ss�pl_Y���l>y^�\���$IKK���%�k�j2�Mc	���o�Wm����        �z��-�ߑ�	�Y����b��@���beC�ד/�U|��ҡV�����脢��\���۩�iE���z�|�q�\���ǧ/�/��2�3y���'D  ''�D��n��v���돝�60�5�1�Y]S��Zl�,9xRN_� ֣����$�o'((X��D""
7ܧ���D��]\���L˄ZI_oצ�Yr���j�;>^�S��`        2�u#ykd/�����IXd���%g�EJLB���%HrJ�	0%$�H�m\� ?)[�Oj�	�:�J��}Kx��x�_{���^e��j&uo%������8k��aW���p	��5�=~�8�IL�X�e;�*�6ZU�K�V�u˗�z�KI�RAn3w2V�+��go�h��z5�!�uj.�?�-�w5m4�9��t�[M�<=��k�5��M�Q@�{�׭r1*N��I*�ۮ�W�'�Z��84��Ѹ�R���m���Ty�vyu�F���9Pl�*�gl~V��U�>;3���[����h�ҰR�l���'%�q��!��]�#�       �E�k\K>���ۄ��GD��3a���E�S+���Ĕ�<�K�<�*��V�+J���{��Ұ��ZP����]B�񫤤Z#�ǎC���tm8q^6�����.\��s�:n�Z�G�hP�F� �*�M`���|�	�5��ս)�g�����0P~<C6���>�e�ޞ�&� y���}����ҠbY�����x��U'���ۻ��W标?�ַ��ΊmX��#�������
�.��ա>��
��:�gg�J��Yu��s�ӵ�����e�8�_�%��G"�̿U��I)��.�       `B����7}�l%���d���mݖ��r!2��֭a��W�2e�As[���ҿqmzK=�٠��Y���]훘0ك��D��x\?��]�*��P+c,�\~�B���T���`Ʀ��b�!{ԯ!�֖>k����>�R���?��L��T���{����l�X��	�)=������y�Ѕ+7ݮmzs����{L�X ���B}v����u���V����Y�_. �­U%-%Y����      �ڴe����H���X����2k�QY|���8�Ҷ��a�~�h���-����J�:U�J�qyy���_dZ��}r{��mc��CaW��-l��S�ѕ���.Z�I�حMj���e@�:ٶ�r�;l��a�s�n�ղZ�\�h��� g��M�ΉV�ժ~�� ���Cnv�
����C�@��,��q'�`      �L��hk�j���.T[���{���;+i�2����BL[�N���T��H�����ɗ�����-���0P��RO�D_�;���l��b��I2g�Q�hEȻ�5��;�b�v�/�"'�D�l�c+*�b���>�� �'_o/�ύ�`V	��i���v�wN�͊���Y�5�� p���?X�=S$҃     ���:�{�Ud\%,*V>\�C�l= Wc�Ū�\�&��R^]�Q��B��ZJ���Ò-HTB�<1c��ڞ��{�Ȁ&��*�e�W��g�v�5GZ�����;dt���d�Ҹr�B{<���Ƿ���K�ޢ��l<q^6����� 8���=��(f����Y-�f��Zu��>X�> ���<�(�e��     �������][�Ð�Q�������ƽ��,�BCco.�bd�ӥ�o�V۹�C3�IH�g�q�������L����H�����'�ϗp��ܴ�d���2�uCyap�^H4�Z��w��Lu�������U�6�e*�fE���
_n�+���߳����� ��7+���||
��CV�_???I�B�v�#�       @!Ъ1Z��#��pN�l��u�|�~�[��"��%���{���]���M
�y�Խ�����V�p�6t�>�7�jh���5��U��ݷ�FjZ�	���{L������P(��T(#��&O�Z%�N[0O��T>��7��\v�<>}� �+hE���*�/U��ĕyt�2�z�-D�FhyD�       �B���>R&��ж?g�QSUNۑ�/��-��6�=�}�I!�U}iH7S	Q+�9�˶��ٮ��Ĕ�x�Nyw�6��/:5ⓒM�A�&���n����1<й�,;xR��wѢZy�K3���em�Y�|����l8~NƵi$�*�5Ǌ�ۊ#� \%95U&|�P&th*��7�:�Jɕ�8Y��iɮ_�ꢝ�T��e���=|ݱsR�� ��>        \L?T�������Hyf�*Y�F����z��|w�<շ�Y|��\��W��'aQ����LO�j#�ۖ´��y���+�p�U)���ӰOg�C]Z�
z�%\w��������ۓM@���r��9��xy�^*S��uj.#��+�.\qjK p�Vf�~�~�ܨg���r�V��{v����  P�       �B��Kʿ�u/�m��{L�iY�����&����2gO�|=~�4����}Z��ۻI����K�
d�w�kb�=v��p�|�i��Nb�����-[O��ww��e�]��
���戞r���ʴ��[#{�g����
��"]�;��I �"=�Mඛ��J���w���k���	  \�`        .�Ґ�R��ץیON��]#_o�+ōV
���t�ψrw�f.߾��S�4Ԅ���_~�k\K>�W��O��V�{p�9%���3��{�LPS�:�ʈ���mޮ	9+V�H�VY����W(-��Ց��b X�+C��ʪ��7������IJj1H� ,�`        .ҡVצ�K���w��n��9wI����$y|�rӢW+�����jP��	���r�h���'����j��?\�C��x�$��Jqu-6^�~9O>���m7r�vߴ��ޞ"ɩ�|�[V����} �H�kW�qL�R�rK�
���E ���       �Z��Q=]Zmm��K2拹+�~�~9x��p��ٕz7�)/�*��`]��[�L��zh�����]�;�
v��s��-�'N]"��c���]��ƕ��}��˗��%;�L.ƁP ֦�>G�6+��j�  (�}        ����lY-��Ve��sr�7�%2>Q�;��������o�fUʻtۏ�jc*'��y���h�`ƃ�]DT�C/ێ�r�j��wii"���V�S��	�k�
��If�:b�Z���Q��9�!
���"cLe� ���.  ��>        ����C�1��˶�p�1y�����"�YhD��d�L��0�\�����c�ȁWLh.7�2������m��mS��̄��-\'����η8}[e������k�j>X�Cƶn$%}��h�ou� +J���4}�aS5;����3ע  W#�       ���޶�4�P�%�ZrV���b�A5�� #?�#S�*}�t�v�"��6U#l�!;�����K�z���>^�S�_��T�C���yz�*�\R5�����߹���|�\�Xվ��e�w��	�L�_��m9jZ9s,��-\/jU��U���;�2�3�  ��`        N��'z�uɶv��(w}��P��ⓒ厯��w�rI0ˮn���ٝ���*5��Ӌ��ʘ����[�]^\�^�}���D�<6V�Wunkg�>ܭ���t�X��#����˸6��E�
��$kC��/��g{��Uh�~��3�~̗1*�/ ��sT^[�I¢b ��@�        'ش�KZ��\
��_͕�D��SRLE1m����}�֑g����,�r���_z�&j���&O�\)�m�'ț��$������;�\I�nkb�����f�����6�}S�]6Xb�d����}�g�vP�x{yJIo)��+��%�[����JL<��n$*>Q^X��,>^^��;�^R�T�D��\��  \�`        N�x��N�Flb���v�\����?B+��f��~x�t�S�e����e�ً&e����[\I��˟3ע�i��?�f�t:�����C3���]RX��J^�MJxz��vg�&���YS�R�/�F�X�ս�BK�`?)����՘�|��mύ�XIT!�4�׬Jyi[����^I�W(-5�I��@���~�ke��1r�J�
�*/\�-'C��ūnѢ�f�`X�Ʌ�h�/b���>l�2���F��}=Z���y~�:�t�  �l�        p�&��I��՜��'^!�î
����d����1.���4,��]��{����z��C"M�%O�&�W4���ƽ�@�[����z�����6U]��Z���Y��[���Ѹ~r�����Դ�|9~���W=#�?�-���ؾ2�e��?;g�|��*���Y(-�s��=���U.ٖ_	/��vliV�TYՐW���]Bj�+e����j8qM�YY���,=t���A�2���w�:��k���;��	��E����U�e��]��2�(�������) ���       �$�tl��m|�y�L�qX�Z�k�W�d���JU�P��W&�7D��D��?L��]���?殖�6���lP�T�r�ꥃ�W���(ɭE�m-�0��Kפ(�^��yΆG�l�z�Њ�p���%��.-L[��Nz/ж���E��.�w̼�k�/�"���wh�ظvM�d����o
��i����֯g^?  ��`        N�[�Kno�ة��*}��ZPpN_����[(s'�4��+h{�5��\��e[�Uͫ��~�;��4�Z>���q&L����P��eE�n����`�h����ַ������U%�q�kW.��>��yg���֯[]��1��
rpmɬa�Gz�v�s��5�Z54�Ν�Wn������-�j�����[�����(ۦQ���Z*P�֭&+��  ��`        Npk��R6��i��Bu�i!�����y�������]�MW��~�yD^_�I�@}�u�V�+����ȡW�*�;'3wqjӡ��6��n���@Z�C\�J�0�Ѯ��w�VqUq���78�VC|wtoS��0i�Kmi����_6Ȍ���0
��mT3O����M�T�O�uU�sW�L�  �L�        pm��L?�:,kC�
�c�փҢj�Խ�5����G�-�t{o��U���tm(���[#���1���ϻ��h�@~ز_\E���g¤S휫�m?}A��z�KK�ZUd��P�o�q���P�Z�KC��Į-�Ze3�����w��m��/�|��ˋѭ��^|iK��/E�JŠ�ǅE�  �D�       ���]B4���G'$���_'p��毕��H�Ƶ�����ٻ����G:
���Q��{�ǖ��6[��l�n��MO6�W[,����;@Q�~��t��sg���=�<���)̽w���yS���ˑ�_ �N��|�� �گ�f�!�`-�n����\���)�&]EU1�}�E�}Sڱ�O5]���ܥa`�V��щɈM����H0\五�l8�U����
�J@������RaЊ
1���y�pŠ����x�:cX�F���Xz�$�����Y��?� ��n޼�jժF��j��0�GDDDDDDDDDDdf}C�k��%�[��4��h-��&�����^�u7�s1���H���֪��M{U(D��ܝ� Ε���Uѧ����xip�ە��7�l"��e���-C�¢-��p$���&��-:xg��Y�>e;37W,xlZ���g.��cɡXv���+���}v���`o��4:6ܫ�mB�d_�&Ui��L��7������*�y;i0}a�fd�䂈�233�����S	�U�^���[ W�����}DDDDDDDDDDDf�?\��7	e}���2����bݳ���[%!�'Y���+ ː}���{��Ю�ܾ]�j�դ�l��C�sZ,S;4U-d���Xs��C^A�l�<����;��Ʒ��a��c�ݷ4���j�qYʬ��1���FZu�>2�ܡ��/��~�����_N���#'��/�nT�h��z�OL-eofn�����p<���������||8��{�.�ߋ���F?"2��u������I�/=��Y�}B�Ϸ��|�U����>"""""""""""3��$H���|�6�Yر���>g-fL
[-��ߦ��i�,�۝���5��	�x�O�x/,ڌ�bvT,^�U�)o'�x��M.e����1�;���5�j�@���[��2����1cO4
$mF2�W0�������	mB�nc��2��L�E_Z�o��n��O�d�����=�,$�7����pC#�딒������Ha��V����`�5���kjr�2��mA�'Ko�ۃ�w���w.	���	���Y9��'������������+c6G�l�F']�����T��*�[$ܳ��yՐx;�.��]�cn�ش��e�	WT��*晞��ܲ�?w	�~^�x�>q9�g��Ǜ���fO#ۙ�L�`:H����L��ߡQ�1�WV�れa����a]w�ޘ�vDd>z	�Y*�V՞/�������������̨K�@�n[ڙ���Y�[kv�y�7�D4���1���R�C�u|��lk$  ��IDAT� ��R�A�����~^��X���9G��uK\?0<X��i%r��Q���m4�'-eҴ���(�ߧܮ����e?�>���Z���Ne��1.��_���<X�4���r�گ>����X����ol����S��9{cM���<�y���P��1�O}�az�V�vsUםJN��wa�~�7�UV��Y:�V՞/U�}DDTn���W��ȫf�Cײ@DDDDDDDdM�������Y���{|������Ն-���8k��)2M~���ǣoh}Mn�W㺚�^��P_!	����*����I�XV��X�I��5	�ɘ_c$H9o��{����	���X���H�F���E�#�l"~|`0|ܪ[�~�6k��&�ω�u�&��#S��߾i��I3�דb�m�ǆޞ�f� 5���M�@D�a����BnU��R�0�GDD�v�����)՜q�Z"����������C��&�+�0Q��֖���)?,Æ�&�艴*-<xd}�^��}-��B+��O�д�u���o��]�[!%�`���e�'�n	c�K��7ZmWG�a{kI�c��2vW��Z3�WHF;�l����b�)�M9s%��\T_˾.u��3�Ec�u�f5���޼����^�ˎ�R�jDd��Y;�f��[PP�7������l�SK�ۖ`�͛ 8q9�g�����=JL���/�҇��O�P����à����0?/5��4���㗯���m4�'��Ϝ��)&�����hP�ɸ�w.uy}�p\ON�O`2;/_�&Hcd�w� ����v2go��`_u'G�n�?�>��b|��R�;��aL�&xw]$��|,v�Kȭ�=_*�������������$̯�fA�_�yMOV=�7F�O}�A�d﵌,�>d��aM̙R����g5��ަ��G�;�t��(nym��x����w!!��m.K���u�gA�'���:��-�y�N_DU%AR{;�'0�?.(n��K�I�b��*��)�W�ӽ�u��*{"�8	����!3S�൓�rr�����8~�x�y�T6�������������Dڭ� �kU��ּ�r'���_�6#V�0VE����س��$��ķ�&$���%�s5#����\GƗ�_KCU1;*/�z�������,��7�����es�w^A�{ln�:F��\��o�ك�쾶a&����WR�~�c�ϐ.FF�K V������2�IJ+{"�;iii*즅��88�C/�U����T�8qB�����1�GDDDDDDDDDDd&aFZ��a��s �)�y��Z�M����kB�g��?˷Ö4����?|�2�nñ���J�V��ޚ�d�{�#����&����UjL��$}ip��f��75K�or;�!��Q1���������)�QUui�&>�L.�mb��}�_�:�l����/����)K����`�����6!""���#""""""""""2��]�N^����W�ۣ{����BSm�g���q�������Ӭ��ջTã��8���=�@�Bzv�Ю��=��W���-�WP�t٩���h3r�-�~&#T����m��n\J(�^}�e��P��lS"�(�qo��e2�SY���!.��4u�		B��5�i��>i�3f߹$�&^�_��`5ڸ4?�>��lj��&��h�Ň��Rӱ��95��	���rg�h���Im�ѵQ���_n;�#��&2y��u�7g'$ޟ2rrAD���>"""""""""""3�[�]���~�r��-c��bK�7��϶�Zx`��Kxg��sPgX�~��q�*�ݣI=L���*����n�m��z�}ǰ��EX���$M�}&ӊ4Q�{�6��c864Q�ߋ����@N\NAU432�h�O��&�	����֡&�h�,Gӿ�Q�2�^��UUgG��~#�˗>���l�˥��T�O�}C��:�l��_��v	�;�;��o
�[�hzv�[��m�"s�*��jS�}��D�u�r�����={b�0��:��bا��UH����vL�Wc����Q�x��M&�q@Gj� %A�A�̃1�GDDDDDDDDDDd&u=�����Ù+�����m��i�g�R�6�Š��6��j�����k�����
�e�4�=�1���a��Pt�u!`��S���Vu�;�Mn~O��)&���������O�-�Bg�VG�FU6�e��e�/{K�.9t��e�6d{��>!-g��ۀ���@S/��o^���ӈ�I�[�1�W����\5��W����4 =��OWg5�[.+�����M�>�}atOx�p-��Z�B�Z�hU׷�����	�b�������������$��V��{297+6b�,O�|��`6�q"��+��y��a��� };xA�f0i��R�@V���ai-^�]�
��ᱮ-�XV�����U\�@_40����IղD�\ۣD0Ƙ��ϡ*+m���W��'37K�����F��h o7W]&*JB%�OZ�I����G�*��e����=9�=��r~�Ͱ�F�M�����u�5
Դ���U2�W�]ǁ��;����˭`��CǡW���gugh��:YEG]ڢC.c�cj�%��/�ҿ��ڴoj���do����I�J�v^��g���*�v&�x����vM�*�7�D8J̊�ފj�S�r���>������':�\����r����7�d�O�!2^���PYHP�����6��O�X��yX!��Ր���IS�9��w//i���ఢP��,}j�Z�]�vǺ�G(� 1���H���^!�G����Wo�٭.e����.�~ƞh��}DDDDDDDDDDDf�����Jcَ����}m�`�Ҿ7��ABj:H��qM��<\�{���ZC�©����qG�O�����U�֪H�`d4������!��ҭ�ٯ����C�.��{c\<�b��{���b�u�e堪�ҡi��Us�Ɩ�v�-���4ԯ]���:DT�`_�`�~xx�1��f:�{+L�~v�b��=97xlo���gG�T(��D�V�1V�x��\����i��Jz%-z������}f�é������I�R�?k`���������������)t!��-[r�J*v���ZP,A���V9U��3��BZz\L~�7�j��C���\��`�섉�-EU53*��~��2Bq`�Xr�D�ok`�`��������d���B��r#'����֫�^��ī���QZ�����&$�붤�P���گ���~mU�Wס���z�m��B��|p(ڿ�s�;L���nj<n��X�������C��g{�V_�>����f=' �$i����2���y�M����#���i�Q��}DDDDDDDDDDDf �-���l��#'-�[|�D��.d}�ا;3�Dvi�F���{��������C�����e�ۅW(�7�}S��f�t��������f1�ƞ-������Χ\GU�'$H�&L�Y�mn�a}�o{��2��փ}S;4U�>S$�7�c3��>Dգq]���V��Օ;UfE�}}C����}zי�6��Q�խ����++v�?�2w�O��z6������Ǽ�Ǡg�����6�W3�9'.]��}K���S�J��������Ѿ�u��H�OF�UE��3�6��D4�cY����u��Z5�"�����>��8S*i�*MR9^�ʪ� �����@\�n�dr
��Ѿ~��Ƿſ�nCV�S�M�z~e��6��u�n��耏��U�Xُ��~�·Q<h����$|��섴�l]����/�Q��������ぎE�v_u���V�#""""""""""23�j
1�g{.[��!���H;Z��e��UTtr�SUC}�fF���{��6��t��2ocB�0��!mN���tq*uyrz��I��`#�l�u�g�*�8go��`_�}.<x��<Ǻ�~<���A��塚�d��݄�Z��-�:�l"���P���1!��U�I6�#	�U��[rT/���T)sG�EUN������c�����������������5l��oY�W�m�������̭�{�&`߹�R[�>�z U���Ӫ���~?�}�r�&�3z}Vn�� ��I�Oi2�ߪhB�P�1e��ػ�����ƈ&o[Zm9ط�Lƴ
)u�]�@T��`z�V����G!&��P�1�<���/(���&���W�u���y���<ܹ9&}�/pd/�4��ﮋ�዗5��^M�T�VH�}��x��}DDDDDDDDDDDf��x9Wg�m	�e��jU�d[���x��̭����ȌUX2}��r�c��;�`v��Uf��8<�ۇ�Ņ��B�@�`��i	NF�{]&�Jl�{.e�k9�o�{H��O;��拋��3iKÛ���Uѧ��vS۪]G�hlty�� z��B�uآ�1x�w[�{�]��v?�>��r������6�ؤ��`C�]�VM��������h�S����j�HSi���#i���s�a;^<}4z}8g���Țd_�dB?�/�]���a_(��~��>9��;������������� K��O�lΨ�M,v_Ú7���-*PA��U�`��,��;}%�ߟ��{����`��8�������9	�eƞh��>1�}S�����Njnr�,'�}-�U�W��$�c�������l���}2.\�)��������.�/W��.������,�6���s�v* .��?�]��K�����%�w-#��Z��K6�}�q/?1Z�����#�\"k*�/����d,��f����c#�Y��A�F�>6�ٖP��h]��"�4����F�m�bT������&P"���W�T2�hB�g�2���q�B��ې���2�t\k�=�]���'�C�dLޕY���ޗ4�98�n�t,eme5�C�R���{o!�����rz&|�\�.��.ﭏT������dtxg&�G��u �QiC��ٹ */	1I�I|������1β?��ֳB�X���P�8����xW?3^{6��޻8���E������}a��F���&.����:}Q��������������� ]����5`IYy��$�&�4/�s`'�A�%=Թ���kɱ��Fd�Z�q��x/��G렌����{��A� T�~7+2�h�����Ã��H�ᐈ��=��������^]�kb�@��񧺓�����U+�'�	��"��{		y?^����h�l��N��y�"l����qH]���^�'㯦��;��6e�t�~�&�����)���8u]�����g���B�\?��O������xm��DR<�>#2���>"""""""""""3H�������%������-	���>���k?��_Û7��ɇb��~�b��������}j�[E8�۩���#�*J嶝<����m2Rv�Yˆ!e��\��FǟBvj��\��%��ܽ����͚� �E���+ú��o7�]��`��1����1��,3'0�n.�C����*hjʜ��f	��
�����t�O~�m�����w߹$\�������vAu��Z��,m�r.T����2Ή�Λ
�}auj��d_�쯾���j�VZ��U���s��`��������������r�ԇ�P2&�ϲ�IH��*F�<����m}��ê�:5�Z���}iٶ���1�B���Aw}��g�Q�N[�QP����y���ҥ�u��7�}�
�t�jF���5Xm�G��3�; �V�*9�� ��{u�	2z[Ҥt�J*��H�>��t����6��2���1�蛻�t�WEH�(:�j�4ft�&xa�MZ��o��i���5!\0cO���lFf�m6ג�5��T�����R��~%޽Q]�y�	�������u�u�I������<c˓��(����������mV��o��o_�Vl_�?�i|۾`��"��^|�M�Og�������������L�n���y�}uj�P{�o��d��R�3��9�Ĵ�%�]������[Ѳ�/��U�O_����6���p��l�~032�h�O�)ǵ�[]7�]�
H��(��g	�7�2��r_��ܯ3�*����  �~k-҂�K��or�<�3f����,���ȣZ6V�8[!/����J\/��#��q�,�Χg���v���\�u�}�p]cm|��W00<X}��X��qW��KJ%k��}����.�[l��{�0�GDDDDDDDDDDd&��S�ħ��o�m��Ş�4G<۳������Ю������F�>9�haHDC8ٗ���}��?���u��2��.�D�o��1�9�Xr�$�ޕ�������������2�'�[a˜1��<�Y���3�����ھ�M�����+NB�Û76�'@T��	�XT�1�>���V:YF>K W�I��5s���V}ݸ��(��(�S��,��֑�+f��ղ	<~�LN��3�5��>"""""""""""39�����M���)�����KLX�}m����Xl���O��u5�]����4���t�"�1h�C�;��-}�	�hT�&Ƭ/:x��F��թ+)�.��{k�h"H*�r���yip�t<�dK�4������enr.�:�Qỷ�Q���	���o����;�y��uw�����j�{�om�s,��uݜ�0�Y��﷜8"k(�ЫI=,zb���h��1t�}��=�6׮�`��ę� �^�	��t���?O7W腌���~���,�o֙0�ڨ���m��ͱ�bj�c���SҬ�h��>!�i�\��ۛY͈��3�;|�r�˥�G��ʾK���L���M��I��;`�j��>�]C?�T������#�֨��\P�;���w��eo��2����u�g�w�j�Bhh�&�]�Fude��Y��[��+���QUH;o���7o�}�`k�#""""""""""2�Ce��Vx/x��+dC��Θ^hS�z�o�V���g��G�U�U���#�����*�c�<��TK�IW�7>I�P�݄�a����*��Ϟ���Z��<ޓ���Z)��]����lJ��"=�d�^_�S����ղ��\զ������yۆ�u=_�p6�ёxu�N�?��M���~0�Ec����h��?��~��
��E+iiiHMM�����v��ꢅ��^�oZZ�8fM�Qt �l0��`��Ș,��`gg��Ѽ��v��vi��;D@�&�	�ʣ����q�>�k-\�����3�8�,ي���6��|�~�}T���h��>i��`\o�g��lm<���ff���k����h\�R��;9bt�&�#	��		��سл_��S=Z��DJT����'I�%	�M�n	�?5�}<ѳI=u�P�\���D���¢�X}z&����\��f͚���I�/''G���f8�yxx��+{�O��I�F�ϴ�Vd������^Ƀ^9;f!���':DDDDDDDDe���Ct���1�m?б�}:ѡ�?��z�����y��
g�u��Z�;�i4���4 ]N���C������.=;��<�ڶ$@%��o�0�t8����z�`0���;[j�oHDC8��#'?�Ѩ�������Ҿ�M�_�������v2����Q����ڒ�g����A�0ٰ��]	��R�!s��x���.�;��m�R��B��Y"�W���$䗪��B-���:5k���`�d5��>""*7=� =?6"""""""�J����I������]���R�H��Oӆ� ��ծ������]����;�:� �-=|R]�z����#�\IEv^�B�CZV�=er�1[N�ǹk�7N��Ɯ���[�\^�p��R��UFS��so�!�«�+��Ȅ޽�vN\N�_��GX/u��A}$�����:6������*�s9��m���;�X^9wu��S��_BJf6��ҡ�B[J�5�ޯ5���{�o��sw�/H��n~No�#""""""""""2�m'/�"��ls��f�u�::`�CÊ�l���`<Թ�jW#�Q��:j��z�<,�|ʭ����:����^���!�J��'�B��Y6:N��=YBc3�Ѯ-+e��~��� z&!yS���4/8�.�.N��3	��4��>�}��ܤ��!�B���꿖
�Y+�W�V�}U�}DDDDDDDDDDDf$㭲��U�������ۃ�t�7�T62�����U]_ؚ7G�T�+�	������iAZ�,������[�x�w[t2BV�.Y��!�b6�8�����p+s]��I#"��[�D��鞭M��/�~�lĕ��ߦo%c�-�)Ǎ��㠝�#���`��#����N���<�i���hM�p�M���u��ڡ�B�j*��a������������Ȍnd�bS\<5m`�ۖ�/i|u�N�e�s`�
�o鉳�=~�6�>��ư��HՓ=ZC+�g���Ky{tO<ڥE��$�3�u(zyb��U����������m_��!ӂ�cU���#xʰ�
����놑_.De!��va&�����Yk,6��o-tn`t��*����E�+]����x�c���u���oُ�W�B^A��<��+�u����	og�B*?�������������l������][���q-#d�[6)W8GϤ5L�}�?���+z�Ks5S+[OXn��o�����A~��)_o?�eVd�ܧ}��ib��v�.]�R����M�ӳI=Lh�����2�����&�K[��B}b���j*�'�th�m��H8r��}�_X��K#������}u��5 �{��P_��p�����6��0�GDDDDDDDDDDdf+��Vm8��.����g{��++v��ס�?>�4��`�-��W�w�]x�^���:*z�:��;hzkc��R�6kT�~0�yc��9����g�ɰ�r�r
"�-7N�����!��������c{�1��IWa릴/u�<<�7G�P-��H��?˶���z1�y�;B}�Ml������@DwOZ���\w;��ݪ��{�`��I���SЫI=Mn����1;2�/sT����rǌ��v��bz��8p.	s��B/d��Ǜ��y�O�6�l"�]�g��Q���f�*9��'�R�k�����[��T5�mU���r	���s����ϻ��P�f&�qsv�Oӆb��lzl���3�4kdr���\�8z
�$�E�śl3�c����Xt�8�B���Y��>�{S�Bd7��O�`���i��}�x�����"�6j8;b�C���^�͇���0��s���7�Ҳm�Ld,�����/{c-;w-��u�\-{�����K�B�����T���M	�eO�Ũ/�bj:lѸ֡�җ9���<X���
��)��*��S���_%<G ""}a������������H���+ú����&��;$�Z6�Շ����]5|;e�x�2rqt��GGb�'��������>j;����q�$���A�L����	��v׳r��/k���ѥ�����Ixb����ks�ڡi������B�(m��7�oh=�q!�:��ܵ�G<��DD�1������������4 ^ό�Ɠ�[iv��]�/"1��|^޽�V!-l9q�<Jm�2'������d�M��ԣ�w1V�"��M���X�٫i����xsd��%����Ƥor���ҭ����:F>2�"c����'��x�{�@��VS�RG?'�gbc�9X��.=rۆ]nW��k��7DA��-5$Yp�a�$����`������������H#_m;�'��TVk����L��_.T�L��=ݳ5�k�4�X�U���rԯ]��WG�||#ABi��ůH��ݻ����\ﶚ���X�[�6��0���:	<}�e?>޼Ϣ��������'�Ң���[�]�[6�,�>������d��S�۳I=<ڵ%���:M�ھ���_�!�� ֲ`�1��>1���?���c��@��q�tint��k��hB2�����`�FN_IŚ�3���ukT��j���[6�Ec�:��E��jF&}�L�]���g��OE5m���f�_��_-DZV��թY_L�Y�����L̎���ۥ�O����푔vC5W	��B�Y�y�������k��؄o����{񷅛U ^��e�ѱ�um�.1�W�H��g��\��ˣVu���F� o�		B/���!n�=�MX��,����I[���|�c�x�cp�j#փ�nDl���O;x������5�1��ǉ���#""""""""""Ґ��i=���;a�$l>n��z�A����j�@�CY���`�O+p��HU	L}�1J�,�m�<6
c�^����iߚ��P�as�r�]璋�Ʒş��Cx/��዗��H,>tTyI������8-a�mƵ�,�пc��Բ�n�B~�BJ:�n =;�y�p��C'GT7\j�8���~�����F'\��r��V�[S�\I��@佒�����xWӁJi�K�O2�_o?�ov2��5��D���1�GDDDDDDDDDD������\�����>��0c�P�t>��݅N����!pv�����a�zl=q���_]���*�a)������G�&,i��@�4�����}���U�!�D����_��5����}J����G�H��\�[��d��͊�&>�4�6�c���S���6�UA��������������ղ1��h32rraiC�5³�ڠU]_�~�;�ƻ��`י�$""�4������������4$���l�?9V��qwq�/�G������
�P���I��%IXcvT��e�$���UX��	�m��$��O�Ø��bj:�|�3�+F�lb���~�a����<߷�����	�cN��E�I���ׇs�ߑ=0�B�ri$���x{�r��K#�4ϖf��cЃ�����at����
�͊4���tT�"��w�;$O�Y������#"����>"""""""""""�m?y돝E����R]Ow�}dF~�PW����ƧZ:Է��	��jW���H��X��}�ΰ	�~f<�~�q���J�|���c�����||�� �dR��RG��h�Ɇu��d+��Lt��_m;�׆wW#�---+3�ŗ��p�jZ�~���ap��3�\�c�&]��<H{���L��e�%�}���������6ùC�DDdi�Y���w����R0f�"�K����!9=d��������p�����/��kT+_Y�_���&sQj`����rǆ��ã3WcU�i�qӻ�Ŀu���}�i��B%�^5�\���V."=�ѫ}?�E��wo�F�ʸ{���Ė��@<��mߍ)�K�;Ogms�XZ��s�@4��ĩ��<��;F�Rvqt��6��p�^Y�}DDDDDDDDDDD m9�P#k�y��M�����g�Jz�ss�3��j�$i����2d���g6���_K���Q=aI2
q���ϥ[��V}������[�=,v	���`c��j9�A��@{�'e�)���y�f�����{��$^)���%5+[���u&A]�1u@X0�5o����^��o�|�ul=q��[i�|�!���5�`xI(el��艴Ή�A7�봪�k�`_#�Ze��[DDD��`����j'�5kh�ѯau����q���%8i���NZ�^�Otki�����S���i\�b�A��y���`I||sdti�g�Gj��a[ �w_�բ��+v�u���V=��K+�8���G	Y������Q_.����[�.U����?�.BF�˘�Fޞ�[����}ݪ���ܝ��:��*cue|��r%�-�u%()�ٕ�mӍ7ܶ�ہV��Y�H+���%��Ouj��������9��Q��`��ȇﯬܩ�R����럻O�s���LZ���:}C�[��e��s�c߹�����-ڄF�׳G㺰�-#"�[mG�.\FUu+���uma���<��_��B�dt�N�52�]Jي�'ATYH۞\�rY{K]gM�P��ا>�G}-����%1�GDDDDDDDDDDdA_m;��-��c��E������WW�����*j]��M�^V��w�G�=ݭ��L�iV==�~�(�Tk���Z'?۲�7Q�H0��)��?̲�м�꼩�_�4�M�n��[5�U�����"c�}�n;Q��v���������嫢OW�?� ""�`������������Ȃ$����u����pq���}JӘ�mS�Z���c �JBFOtm�W�w���e~׷[p �]��,�u-#c�^��ώ���,�ٰ��:�&�	�ӿ��2�}j���0�*�]���.A�d,��V��p۠:�i8�E�'�B�u�Nl�)�Ko�ddce�i|�yR8ڙ�tB�&��j!��<���+�^��Ҙ�gù�50�GDDDDDDDDDDdaq����5���!],z�2R�c� �a�:���#�z{�����F��z�<���V�9�EF@��z�j�6Fkh�����q�j����Ee5�]8��n�N�o	���>��ܵ��RȮZ5|3e ƴ
)����;�xc|���W�4%"��u��'��D����$�.m�rn6�˅h�Vu}�[��ݧp29DDD��`�|�iG4D��u,z�~����##0cO4^^��镫����O�l���G�}r��%L�~����~۱�Wp���Ոeg�4����<�1o�ٍ�v5k���j�8��1�U;�5HX�љ��f[5�{���₽<����YJ��:���Ԯ�Rt]����L��������K�BDD��YA^A�
gm��DԩY���?�CS�����=��&'��4K��F�J#�5����	�.Q#J�"m�SX��Z�Oȶ��>*!#��ƞ���0�#�[e�,���[m�%��-J]޵Q "��q4!DDZ���-�+�do�O����������͛7Q�Z5TU�������ܦ�;B�\� ˨戙�m�vQՒ�vO�^�_���Y����6�����܉%�N�d뚄�^�}C�[���bj:F���gh~_�����)����צ��=:{�����69�9ԯ6��=�8�Ỷ��������::�V��D�{1�GD1�MH��m	�?ѭ���F��899!3399��A̽�y� ի��=��|
���e�O?�#"�rk�n���-����Us���|�^[����j����'~�0�\I�[���G����k胧����6aV�		���W�{��E����!�'���Q��/_÷����h��΅�ի县�m�Z,e��5�9����o�����JZ��3#G��"�Z���N˺> "˫[�.Ο?�����������z}��q�ٟ/����¢�dy��ʱ��DDDDDDDDDz���(����f���8�a��Q=�����Ø�7֢!��qy1�{Ktkd�f��
C}��0>U�}5��񄾰�I�F�Zj[�ǠΘcؖb���%�Ix/<ٽ&����u}�|�uL�a9��l���K�oǩ������]g.����T�:�e�CD��[ح0ԧ�=��P��}DTa?��[RDDDDDDDDD�&�o��Y��O�T-t���^/��wTbs��b�㸚�e��Ժ�/&�Ǹ�!��
=�f�����hd����tR+$㞟��R]N~?�����q8�t�*����C#�.�ѥa �"#'��[f�Ζ�������X���G�!9=��{�V��/3�-~Dd~;O_�c][��Ύ�Y�^�nZ��
������##��>�b������������H�g�`�7����qj4�H�[�`uy{T/�p	���æ�x�9��,��j8;�g�z��O.n�#i4��"��A����n�䩱����ٮ_��A]�^M��cg�xl=qiY�}���ℾ��1�y#o��-=�0��3V���˨Lv��X�O&􃇫s��7o����5�Tä�>���Z�D��%�ջ�.�,���eɡ8���o�����z Dd]��Y*�W��ϗ�>�c������������H'��k���q�t����UC�z~���>�T�/&������m�������*�T^�����k���W�}���V��g1�W0���HH�܇eYy��Ӝ�����	z%��Ý�����.]þ�$�=��#�U���bmn�%���>��W��A�h���m)��&��^�UѧQ-=|�N^��f����Cg�ĜQ����K��Ķa%~F��y���s����GADT^�*#֧v�Pa�Ԭlu����]*P>񻥆���w���n��WT��T"[f����C}���|���ȅ�����|j,jUw�^�8ث�r)NBZ���|H�������� �p)((����j�����]UK���ʲ��yL�~��MswK�D%���^z'�ma~��er����R�e{����kY��)9��Ӱ-y�����2B�~m�=Z�0Է�@*3y�~�sg@oD��w��
I���Q=Uk�Eg�H�$�'�{��Z���<J�3��6���Uͨ=?���-�ී�=���������Mr^��9s���?���,v��ܸa�sK?_��l�}DDDDDDDDDDD:�xE��,xl��[׌��V��5ԥ�Z|�����"�W2δ��s1��������>��$���/k1o�1TU�څ�����cZ�����@DT�]<�W�����2]ߛ�������D��3���T��ڡ�B�|���������������th����W5�R���n��[�7V�R̈́z'c~2?O����!'?���N5DUe��k���W����;D��<L�h����AD�C�nqqq���fT���3rr�����8~�x�y�T6������������tj��K��|,||=�A�s#;W5�I[�-�q�c�^��F��C����+��z���rl9qUݕYfY��Hڂz{��^�Z�٠��4v�BHH��ǳ��T�8�Ϳ9��|�l��Xܥk���\�����)�1��8p�l�4��i��:s��WG~<d�i70��%8|�2X}
]�\.��+��R_{�:㙞m04�!j�pA��4̊���{����DT�I����u�(�����s�E�	}�.�F&��,��r#""""""""""�9	�X޹��@�z~ �Y}O�Y�������X�&^��ӆ �6G�Z���$�'�2���Ø�.��F����^��:5k`�Sc��۳h�\'#5G4���!7� DT�5����ڠ]��j���O�Ǜ��Ѕ[a鵱g1�u�ɟ����V��VJˏ�T*�ޮ��k�����#�$�9HV^>��g{x�pUܔt=��9�%�ـ��L�t>��S;4i++7/-ۆovR�a���z~8G5��l���9Q1���Mj�3�N���_.������^!	|�y?^_�K}����%B}�Ɵ����k���*�1�B�Ť�p��}|d/�j�D����?�7V�� �1������xs��Jҧ�a�a�� k�ȳ����\�<�7o�;5C�� �pv,�^nc�`�a�f�a�7Q�$��?�$���������0�{+ti�b��^MÂq�h�^��@�+�}DDDDDDDDDDD6BZ6����N]��c{Å#U5�t��X��	ɨ��eda�O+0�e��,ct!�	���x~�ud��'}�Lt��/�� {�$�oy{�wHP���H�xgݞJ�%��I��gK��
9�����!2>��S0��_���h�S�h9K��M{Ad|�\�Θ^�]ݥ��R�;9⻩�0�i�˥��Y���<ֵ�z�-l�$�#�/����
]+Ǿ �F�dB?�-���+��N5G?h�7�.ù���_�DDDDDDDDDDD6F��_����@Ow�yH�苭��ʝUbT٢�Ǳ�\��4 ���GB���q����v�J���.��W�?��^�5\q9=S}/c�$��<�ن�x���w��?"�@��MK����N������K���L��&�ബll9qWnd��^I�T�-�G:�=�d����|�x�O熸x����Z�ۓq��ۄ��I�����G��;3��?���Q%C}�Q�ڭ��цsA!�ˏ�Ī��H��EC/�~/m�uj��/����O�#6�
��>"""""""""""�7>I�T�6S�T~xn��*�\"���|� wn��br�!�����j�A����U"��̜�����y��A~�1m(�=܊�˨��.���V��@"җn��bh��*�t��4wo,N&�-o�_v��i������<�.D��W�څ�v/i�l����א��E�����aB��r�\��:jo�mƗ�ޱ�g[`��T�IS��/-�"�l�d��Ⱦ #������R����|�e?�����<\�������|��}DD��͛7�������#������.�$�NDDDDDDDD6OB*�[�ک�ӫd���5����}*�Uܼ�ov���'�úab�0P����¡�%��9�j���up#;W���?:R�ݮK�@�p:��w4�ɸ��>�j?8~�����'�u��<�(�Q�/}�ᥥ�������߂��)�:D!�0�Y#uNԫI���㯦iv�0zlo��Ƹx̎�)w��_X���#�&�	i%�璭�v� �}��1�Gz#����ۊM��aVdt����{�.�Z��o�	it~|�D�m�:��  �C��~�G�U2���HOO/
���333U����M����������r����H�ޘ�%�:�4	�̉��k�v�bj:H�����`��cxmxw����M�g��ޅ/�TMQd>׳r��H�&i��q�o���3=Z��p_���X{V}/#�1���ֲ(8����6D�M{9���ԯ]���������\��ԫû����ycD�޷��)l>~ckm2E�!�Wvժ�C��
�I���P�^�M5��y��oP�B��ϽF���ϗ��O����)�pK��� ���}!��R���hSϯ���v6�nzv��uD��q�C�#""�IS��P_q����5��HDDDDDDDD�������r���֨��s�2N�=�Y��	W@wZg��l�;�)���;���NRYx0ΰ-mǹk�A��`c�\���^mT�Pjf���w������˼-�)����n��;�����튺�����MFoC>�}�G4�F~A����w����3	w�+��'����#���S�Ğ�W�Ʃb�FI[���u��VM��Ĵ*������edݱ~���>�#6m g5�tƞ�jĜ��AU�B���޸�zlr���s�b�>W��ȘƖu} ���O_�;�"��8����Ǻ�������O-�a��cg��5�q,���9;�f�q�CQ���
Kk�4�^622Y~����������T��7n�2:��e��:~u7��Ύ��M���fD5��?�i�ֿ��'��Q�9�N��;5ã��+#:�s�UP�ջTs��\�G�m��&T�fҶ+B���Ʒ�����f��k�Z���?���U�)o^�Km}B��券KWU����U��v=����}ۣ}�?/�E���{���s�ܮ)�wo��'���r�<�4�N�_�c}iYZ<}4Z��+q��;���8�r�X���G�4�)r�/蠂}�:?e؏���+ۗ�9�-	�ʨ]9��)���?��c�a8.��!B}��ʝ8k��+�K���qӮ��mŗK��HO����ׯ�څ3������=�p��j8o�s���2��d8����v0�GDT���݂r�E���d]Q�"!�51g�l��x�W��[d4٫+w�P�N��~�}D�I���
��l�BGt�j�>��ʝ8|�2H[��++v���G10<>����ˏ�*vsv�/�o}4:$�Q��um��DQ�%�eX70,$Ḿ��UP�9k1w߱�f=4\�9,$���֡��� ��\�Z�
IXm����[��:	�N��J�}2O��
�����cT���~yhW�
	o� '�����ľ��z\�o㋉��.������s}q@Gu)N��|��ܼ�y�Ѣ��C��ƈ���swqRAs	̍3<i�-�{X��XD�{]'a6	���?��)��e%(���0X�^��I�m�K�b���iCKl��xB_t��g�/���&MYų0��عA ��d��WH�������.��:g;�6���X�c���J���k��u�Pe!o��x�c�z]:�D�3�vM�2<׀b-Zr�_��W��!�-P�B�z�}d�
� �;�{�т��\]"��P�f�ݷx��c��a[�l�!�����Q?S�\���k$��i?�T��B.������x�
��뫞W�wg� Q۠:%���H8S������4mH�&&!�A��c�N����:Ȱ�J;_��`N6&˰���>�9��ٷ��.��G���㋼�|�� *JF�j�S�rl(���E������"�ܣPZfv��_-v)�a�%�?��>"�J$77�%�2�GDDDDDDDT9IS�4<}���л�j�*O�2�<�4)I0C>����mI���K�d$�P�Ƕ�>���t�5���$���6�a���U��4�.�j36��vcZ5)�P[�P_qP����*4\��&��⡾����)���E��գD��8	��;��
0		�|=y`�P_q��U��ﭿҒ�?�ؿD��8	ԭ?_Ғ��4�#��w��2<�s�QJH{]�P_ql�z� �}�g��+�+N����������8���B�a�72U@AD��[��ۮ����j���Vm�[Q8A6�Gd�
a$��=���ⅻ�.�$w�K�z��=���w�[��������?L�����y��z�ð�۽�	�i�L��A]��w�~���<��	��������Q�+���9�e�ᓕ�fچ�liP�9�}�x�����C3�����0��/3�YR9ӝ~���N�5Q~�l��[:lC}�n�OV'��k�.U�Ӫ��w��j^��1޼6����_mC}����c��˕�?[ƅ��Iuia*�ixЯ�P��u9��7�o˴��d��=WZUQ+̖W�7�ӽ��̧�Gd��_�sYO�Y�;�T�,�	{�C3ǛJc��౶��+}�g�r�����p�~?�{��rZ����kHQ[���W��̞_m�_R�m����+'�U=ii@��}  �*+s����,     ��I�<��&S���3�ɼ�}�;��޳t�!yf�.9�$�F�i8���{�Q���)�Mʖ@�ku8}���S��W=�1���uZJ�ʕw��˝\h/ݩJ�J+��D�UF�����riyYi��u�O�p�~>�d��^�қ���0[m��]������cW�����`���j�䨡9m[��XUm�5.:�T6�p�Q	��N-�SMtY�i�K�΂qV����}a^Z��Mh�E�bpe���1kl[�!�����Cl4��\�=�=���]dYM4D�A���v�ڎ�&�� �|�Y�㴂_m���7�2ا�Ě��e����s�`��K��c��*W�Z�Q�}	�Ι�}M�����6���j+m����τ��1!f���؅,Y��
���:� ����;$Ѧ�^]he��^Z!o�3�|.�z�lN�*�'3r�k��5�,�g��������a�p�1�w��G��O��)R�-��	����n�Z�[U��!2T|�> hFZY~Upf      �8z!S���������Ć����4e�X�#Q^�v@.��K�$��I[+j�.�hU��&��Xް����e�÷iu�����T���Ҋbw��@�Rk8�ku&3��o��F[�*��^m][^�}�j��е>']����k#��uj O�YW{�v�/;c�\{m.-n�}��?�����c�	���`�ڸ��//�+���պ|lX�Ӫ�U���.W�W����i��,���}��c�j]�o��-��˕�HmC/�{�{�Ξ$�u��TC��g��=M0���N[?gɲ=�ek�S�ӛ����~<�zG�ַ��9���Mx���}��dKOV�}�oH�k�4&�-,�^�-����R�r�M(ܺ?�'!8ۮ�3�jX?��@� �?˗^i�k����
      hi���
KO��!�G��oM�R�_������	��O���9uN~�t�i���>��4�GgsP����_k�Nʲ���e�t�=���L�1�~��mťe�m�?�ز��@��?�,!�n^va��&�����9Eŵ����Z��om�
������������c�}�<�̂���ٖ�S[E@�c�.��su�h��ܯ�c��ۮ�.���U,�jɻY{NQ��2WSE@��]y�:���0n�\�2n��RC����=iSM�G�6�y�mhU�ްG^�~@��Җ�Z)s��x�v��.�u�V�|��]���\	�ۏ��6-���|���M��z�F�U}��p�#��N��]����s��j��ۃSG��N���,iض����������L#k�R�o[������+�V�z�� hF\��f�      ���5�N~�Vzs��1-���/O���7�#N_j�ơ���l��L����f<M�ݥI�~.)+���O� ��
�t1dߤ���}������1�~�s�:��M	�3��<miX[�T]��rM-g����#'�e��jj��
mI�.��x�	R�T�NەZ?WL��_;��Ǿ����3�ty��O�=㝷m����R�����Ԉ��.�!L��W[�S�gLT!���ױ��>�gM����gU�kM!O�����5�O��[[�j�r���2��q��$�[����2�6�,��t|��_
Uj�M�������Ǯ�[��֤��ʬ5/�jCC��t�q�g���������,�ߴ/n*�2��&��Jۙ��_n3�������u��Z��9٥1i�O�}�y��Ӷ�^���~r��&���?/l�k���g���G|Ui�G�(y��)ru�nr�KV����0��-�x�sYKlMnض��{�g�~W���ߙ/�n�c���{G+��c�t�+�﷞�Q�Ueg_C� ����`)))�5ܧ���     @�;s�L�t�9 ������A�b}��%4Т=7?#��2m��{4��Җ}fҪ�{v6��i@�Ɣ���g/�j=�����3�-���{_�T�ϔ&�l!���/�o���]�6�ۼ״l�jP���w�.����3uF|����Z��M��W�o�%��uX�M���[_��`�Wn��gMp��ܢby��/*�֐�ۻ9jhP+�Yi���㇘�G4Pf��m����6�q����#)�ٕ?�b��w��N�����ZX�Hi%��Y��_o����Ӫ�VZ�����M�őӖ�^���;ɴ�ӽ���X�s���p��_����#/n�k��R��
�-�#z�5��!�_��(�9i��?���ʿ�[�7�R����������/� �@�~�9�jE�7w$V��ہ�1��&���olO4aD+}��y��n<zZ����<}�zt���m��硆v4ȭ��t{��/�-x���~6�~^ח�o=5�Y�ż���w���t�e4����y��Lx[���f�x���F���g���$�߹a[�P�W��ߘk*q��˃SG��*��J���_
����=� ��	���\��>��&      @UZ1���m�'ˤ�=Fu� c{t���:��C��`�?�r�|�:�!I�igJ�l?�fR�i�k �I��p��N�2�s;S-r@�s0ϓ4ȣcI+�lIN�/�������NE��d��u�6�Ӿ�	������[.�]4C&�����a;C�x���5t5����E3�Z<j��o�o7a8[������򷛮����9��l�Z���q��Z�C4��k��U�;z!S��39b�����WI^Q��u� ��V����ڵ]�j�7>��<{�2���6��t�!yp��*�g�reγ���f�*TV�y��58nK��i�(�t��|�B+������U�-��к����	����� X�����Տ�Yky�JM`�6L�G}��6A^}�������rݠ^v�Ѱ�w�ZeתR?;�s�}��ko���7&؅�����?.�r@N×�|��ih뭝M0�9�M2+m9��%�W�d��6���ߞ2®B���r�mj}�n{i��c�4�:ݖV|`�g&<h�}���m�����C���!C���7X����Ig��V�[�����gx�~��>�b�|�;�s�j�u�z�5泹�~}���ϻ���Z��J��߲l�	�����4L�Y������n�ݲ-�c�}����X�w�H��U�����	���ǷU�?��+��` 43�,?�5�W\\\Y�O����IPP�	�      ��),6�IuR��e����6m�4|�)2���������V���4�v�d)+/7�TZ��Bn��e��ٜ<�8��+�ϥK��l��4m��ku<��4����m"MU��1��%:B�C�$"(Ќ'�DZƗ�����2�b^�	ꜷ��t�e�jEG�h�/�&�T��O�r���f���FVC]�|�	�9�-g���k2�WgS�O�kZ1鼓`�V3�V�W��f�.��g���)tkH�o�w�+��˕}��mF�|\�gYiXO�?�f�L�'��~�y�<�氕�V{���weh\;ѥ��\ޚ|�Z`��@�E���7䊞�M�W�iu8ga*�e�c�"],۾ޟ~�8�^�ݘ o�:$W��*mÂ�w�VH,*�������]gB��z�IH���?sQ���:|�Z���W�P�5`�=%ͮ�-}�~�-x�J?ť���ipD��O�b���g�~��<g��4h��th{s0�?|�ݰ-}_4L���d�s��,�{[r�	�U���=�~l*J�����4|�l�j��<��y]4�]PR&�,��>&G4<=�/�D������"Y��b�<M�Oj5�O-�3�>�f�W�Kao�D5$�L�MUS�|�����~��}�?��i�y\�Ε��X����=&�ix?sr�V�Ԫ������2�����\�&�l��m��Ͷ`K���Ă�?�"}۵1�7-�>��`Z����j~�:\�Ĭ�u���E� �����!>�       w�.^�i�������l3M��tr���Zk�Ք>�%�aKCb�T�pWm��R��M��U���$�`�N�������.?�i��Uz�^+v�J���N�|U�s��yU+�9��U]���
�U���DC�u	�$}U�����sur�~�۞ x���̤�1"����|��=i&:ĵc�z"�u٪�mm�n�֧۫�4S��d��S��P�m��mZ�	g�yZ���������_D� �'��f_yպU��۴          мi�:��z��>x�s��)�7���4��dw�,ޙh*�6���\
)k�P������54]V��mUW=T���k�V��O�r��l�Ʊϲ-�s[�+ml���D�U�  .K/iؗ�g��c         �n�Φ��Wʃ﬑�{��W6-�m�t�
��_5�L-�k���u�`�.�-��Sm���M��w)̴/��������j���:&�RXO[��ԎW��N�����Yתw���pU߮���7���k���J�:���\�mHC���`            �,m���=������#��mcJ�6v��#?�v��욱��D�	�9�Z{u_���W&&�ͣ��5�
�
;������w�XtTZ�l�	�Z�7�������ȺCBB���@|E���l۶��'��[�o�4g�^:-�yK�)}��+wΪ����V�lL�            �,9�)O|�U��j�L����f�i��Y�n�J����L%e�Ҕ=�z��8��y~�:����/��-�MR�	,���]:ȷ�7����d��?���\���6��dggIVV�������|=��o���2�p�Q���bn�i��36Jf�%��Q��`�;|�Z�"���*--?��7          @�PV^!�&&��mX�,�_n3Pw��[N�oV�������Ȓ݇�Uo}h{�ﾵJ��y�	���V^�s�����L������������4�W\��Jj��QҪU+��̔���竚s�oh\;39SQ!�▽���k�e_F�@����/'N�8֦M�z�          @Sw1�@�ݰ�L|�e� ��[.<(P~}�x3i���;��=Ir6'_|�ۻɾ��icd����U��j�o��3��}��BnV�&����8�>o?__	3z}G%:4X:D�V����\6=m�yn������h������222̿��          4'�.�#n��?�bBp������u3�ym���L�͙$k�N�;eٞ$�<Fm�����6R/��_�Ą�v���m"$28H�KL�����%#�P|��CnV�c���5���0���p���'�-<��f3u��1��9:²m���ʓD˶��[� �(��\��>M�GDD          ��\����K~q�˷-*-3A=�:G�ˢ1�ht�􊍶[οuk�>���k��k�������N�5SS�X!7+o����6v�BOJ��3�H�4e� ����.==��K�         ��y`�yx�s��=I��>��z�d��_Vm7�V�����`D	
xGNN������o��;�g�X�
��} Z���B}�D�         @K���9���������́=M���>]��+�>+�igfO����P��>�E�@��_R*���Ϗ�����ʖ���~          Z�Ry7ᰙ����k�{
���B}Vڦ�|��Z�}�-�4 4{��pAC�ޮ          xޑ�i���4��!7��� ���ןopp�TTT|�>             ^��Bd��PG�              �!�              �!�              �!�              �!�            Фu���y��zl���%�Yb� ���           @�6�G'3yJJz�M|I �[�             �C�          �Z����� �-*����8���$-;OJ��]�]�_k�mä��\���KyE�  ��        ���'􊳛��_(k���H[�u�
�����9I��%  ��� �ah�&��L��E:X����d��ۻɓ�wHVA��۷�%��P����=Q�ߔP�2#����ʼa}�mX��WV^!G�gȺ#'寫��ٜ|��}d�D�gy.��b�}��v��>�b��h��&�ʿ7�����K ��`        �i�;��Kw\g7/��9�����}�ʑ2gHo�y?\�Z^"� �1��&ӽ�ݼ��	
��Q��ëGɂ�dγ��؅�j�����]��z?k�Rj��ʾ]�;gITH��[��KxP���c�e�����o#g�	j��Cg�M��{L�|k�p�ڿ��xf�	��i;��#�& h.�       ���͟o���u��{_   o
�o-�E�|���-��Hai���w����FI\t�	�]�ԛ���3?zg��;	�%�Kwz��q���{�7-�5���Ǜe�ᓦo��`�9Vn�Wr��WS�o�Z^��z�;|>C�o��W]�a��f���S��]�|$  ��}        ��[F�˼a}^׷}�}  ��\�SVL6U�lie��}􅔖��Ϯ+�;�ʔ>]k���Ɂ�}o]h0�_7_cB}�N���g�KaIi��Zeo��Sfrd���&����}���P�Z{��������i2wHة�H�(  �
�}        ����tzݠN�2�s;�{�   xKmmM��y�	��aq�jm�[W��2�A��e��B}����~��M�N�jU����������M��Ɂ�� �� �       @#ӽ��S�2��(?w�   ����RZ^n*����v����7�~y���`^M�Z��ɽ���Շ���dӱ�r���rU����'�  ��`        ����k]��������L   |��nM�O9�Y�����m"$:$ȴ�ݙrV>I<^�ͯU�V"W��l.�HI3�j�y��H�p�.,��#MV�;&�����=&J�.E"��e�3�Φ�`_��5�d ���       ����o��q��UkK<��;^�P  h��H�oVA��>t��e�0wr�y�����֛��Uu�7!@u�b�����rۘ�'C��9�r�����'���U���9��麈�@s5- �7�       ��0��9�l+-;Ov�<+��������  _0D?�=������[L=g����Sg%%=��=�s�9a!&4X���Z		𗗶쳻���`u��a�%:�T�{m�~��u|s�0�*o�;Wf<�Dv��ܮWO���,(t����*/�� ��}        4�;��}{�!�|�L�`���%.:BNg�  @c߳�<�p������ݘ�p9m�;�W�؅�mz{�����1W��o#O̻RV<a��p9Π������?���
3OOvX�;IV}o����s���.��M��_���R����:�� ����r�U�Z�2�;��狆!�       @#���{�U����M7��
�U�V�����o�w  @c�P��{o�� ���۫�.[XR�0ԧ�/f����~�H�����O|���������"�Y��2�g��vQ�^�K~~�8�����ɌK����˷����l+�v�*��6h��~���y��\\滁)8(���RT䛕2���$,,�m�k
�744�p�!�       @#��U��h������wv�oOaw�m��<�f�9�  �M�P�V��t�����GRҀ0��Ȱ��Y۽�	���*����lN��,�Ⱥ�'M�O�k_�˲i,�ض����0|Sai���t�����ӧ}.�VVV&��yn�)_}�����3�>��}        4�֭d���j��<Xy���Ղ}�c�e\�β����Dp�����n�V�ْ�Zm�+zt�Y�{˘��O�6,�����˾3d��t��aX_��^��iy�r1�P�^Ȕ�����c��D�����YZ֠�O+�����n^~q�ˏ{P�Xib7�йI��u��W��*Ukh|q������6J��'S�t��b$�r��z_�-0�GNɧ�ɲ��)�Eۆ��ܡ�eB�8�f1��w��P�}}���
$%#G�[^����`�E ��+lB}��w��>0�u:����]���-�^�/.��� ��<��Oɸܾ7ڦ��q�J�U�m�mإ�Ҳ����>_�YC}��k����!�       @#�ֿ�t����PZ^n��Yi�>��74���r����`��޽�F�y�o��/W����Ξ(ë��.i%��\�^1�[Gyb��oU�^XCn:i��W�2�{~�l���������<Sҳe�^��:vl[m�Zqhܟ_s��ZUhΐ�v�~�t���e�K�_��y&j��o�k��J�7���`�j����12�L����w�i�xo��>yN�A� �s\0����9\F�N��rF|yh�x�jy�l��NJ �oխ�,��\�����yOr��S�����>��~�
c��mu����Sd[�/_���}���c�=Io?���,=YM��x2�W�W�K+:�﫶�p?_	�y:�g���ԩSR\ܸ�B�-�A	��.�}        4����6o��s��;��n�W��u�W䙪2��[��7L�oN��u=0y�<:g�Y��Fv� �}o���5�����]ݯ��x�uv�j���O��@�y��p����c�������gy��'o�:$���c� P7|{��Lܽg��M�y�m-k��J�YꀃʭZ�U�}z2��ҵ�^U��^>q�@�}8oeb�,/3���~�E��j��q_� ^y0Y��L��E�5�+��'�����y+�gեK�F�]
��V5��`        ^�-J�Գ�|�6�VKw�G��$~��q��ahyc{��[�V"���Y8���u��a& X���iRTZ&竄ᘆ^�{v�B�VZY�;���}O�>Y��d�D��գ��t�iU�y�/7m� �g���x�}�L /1�������_�����S�+���՟o�ʴ�U����̛;�g׌5��Lc*���}��^��I8}N��ϴ�^��j�O+�j����ؿ�(	��3a�W��]���v�Ϫ��}����}        x�B-J���G��U[V�MZAf֠^v��'�}L�0�w ��$��hZڅH\t�9H������tx]qY��:xB�9%�Y�&i%m��-��!F�}�4yx�FA�4���lC}�%����i���93�Z�n%q��yr�.�mm������2�/�׹���Pv�++��uGN����~XW��ѵ�\?��� U�i���d�3K��  4���\_����,�:ݙ]'�V����ݳ%��D��:d*��HdH��le�7u�5�-ۓ$_;]m��
�7�߾v��;a�����^F~��,V~ey<�,�m%e���w�W����&���%�/�a���IJ1�y����oOa������}��nS�X�>+o���5�        �2mWZջ	���^ߞX-�7�g�􊍖c2�]ڄ�C3������\^�b�<�n����qxm�[�����MW�`^U�8.?\��a+�o�cn�a��=�<����Wj����%$��a�>�z�<�1A����p�Ӗ׹G�(��]�D�w��?����}O�'���q<����%�ˉ�l���(`�y5X���~��ko���x 4�h˾�U�}����Ԁ1����D�-[��zm}�>"T~:}�ه����������8����^%Q!Ar̀��{���~�<�f��i�p�Q:�g�U�o��;�g�Ҟ/\C�        /� ��N�+�i�9gV&&�*2�n�JCs�F��c�lv�cӃ�V�E2�?�Ɏ��o��y��Ӽ+��e���>�����n~�}�����+GT{\pL+��Y����%�˨q�GNɬ�#����TK�uۘ���Uۥ�����ՊGO͟Z-���ۘ ?o�Դc�z�FSQ�;fU[�]����^ �'>�jB��8��gγ�et��%�V���z�-;1�r�e��s�Ξ$9�vѥ�����r�؁�R�V{�j��{y���
���w��ޓ9C��M��J��().-�#�3���VFӥ�<�����Ұ[RR����{d����RT�z{qO���

��b�8F��       ��44U�V3ے�ʌ�ֵKv'ɷ&���hL�<����ԝ�J�d�s�eϩsu���ԛ;�O���=j\�zh�S=�Ѻ�XNa�����.W�9��+�|��t�uv��D���d�q�c�j��ҷ]�j�������R������������7k��{W��;^�P  ���=��V���]��XN����u�7Q�}��M:hZ�������Yw�~�����deeɑ#�����狚�       �K��e��~��/�y�� ԛ������U}���N��a��8�	����\m�V���w׹�R��O�����u3UyP��?�T�Vtp8��#q_U��խ�K���&�6O[�{W^Q���󛾔[FǛ�N����T$<��#    �R�       �K��]���f���y���j������mL�[�}�������u[mշpd�j�_޲�T����9���{�g׌��|n����@�o�����&ڇF����-��/��G߻�<�G?�,�|�����[�q�Ǖ�   �	
�a�[Tl�_hz�       �%��Tm޶��E�+^�q@~?g�ݼY�{K��`��/t�cԐ��⭏�q����Iz<�j���
���%�:_m^�6���n\�N��iP�!��N���<�f7|�8  h.�r�U2�[G��׊ڟ8^�rZ!��W��[F�K�vѕ�s
���}G�5;���t|�'�� ��2�C[k~���V.U���~�d�4�        ���1�2�w�j��LtyKv��Ξh*�Yi�<m���M_��q�;|�޷���Ui%��'��Σ2%1��wl+pnkr�ms�IN�޾7ʅ��c�W? �AUG��+��}�����յ��nժ��}  |Q��h�*$[��u�m�䭯ϑ�b�]aٷ�et���O\�Z����o��ܽ-�~�l�&����9�>��D��}        x�mcJ�V��2��=�]^���Zu���سں���}�l�o;�A������Y��S�������z�V+�T��bU#�Vrj��r�=ݯ}*�   �څ�H\tD��g�r����Ε#�U��ɿ��_��A<EO���b�ż��ת�oc��_Rzr��6�$˾Sth�|mx?��+Μ���i�B�|�;��>��8�5E�        �0�4�hL|���B(���N���U�}Z�`P�X�k��29�� �+:G�U�� ������e��m�*,)�6/ȿ��a"B�����1h�q��::D��  ����dr�Kձ��e�_^wۺ�4L^�~@�zf���WH��,i�M]�;nY���cV/|�W�5A�,�տ����2�O����W,�l��-������������*�Z��)"�       ��]շ�t�� bU�X��/�6��v�o;P~��zi��bi�(U�2j�����_Gs�_���R�UƠ���ꂓ1�BA  ��L�ӥ2ԧ~�|����q��5����&t�tIÇV?X�]���я7˕��%ZuY���G/m�'@sr�S���ʉKm�ni*�       �a��J�j�:Q�uik��������_0��<�bS��n�50�(ؗ����V�h\��*$��a�l7�W�N�XF�4�r  �s�5yx��g���]�m�e���
aC�ڙ��3�{J��pIu�kl�t��/���돜r�\yE�<�a�<�h��[���CsS�ySF�  �h~�$6$���)+�p��e�����2)*s��~f|��6>�K�   ���� ���6?-;O�3eD��Pm^lx���C>�{Tꫢ�a�+4�UUIi�4-�|O��V�%nx�4��+� @ˢ����^��?����5w��:����͔�#��_�Vr��x����k��Qy���k\���ds�AÊzřs���T���  -��vQ���1RRRb&G���%;;[�w�|z2S od��vq|�7�<��   |��#�;$�k&w�m���J������ (�-y�ߣz����*2��:2
  �ֵ�=*������In]�3�v�`��ڿ�G�}R,)/����U�رm��)i5.�!��s2�C�ُ���v��3����c[h��       �A�9h��)چ�cd�����W�pT]��"�}+����ZZ:-��V������:�&  �٭c���I)n�����99��+���ex��`�,)kxEj[O/�&��u�Я��KJeGJ���wL^ݶ��pS�V"}�EW��\C[a���&ا�;����G���`        2,�����k��ߺ��<j��}�Ni��W]�D4x��c"�}�r�]̫fk�����Z4佺��(��  `kx��}�5I)��#�3M�/$�_������ܺ��}���l��I���������?�UO8�mX``eJi�6�6�t��WԶ-|۲-�t�-4W�        ����{�>�l�`_b�E�گ�ݼ���JCn@8R[�V��*���n���[϶�!<wY�8hQ���   lu�
��|2#�#�q.'��r{�~��T��[�o��ϐS�9�_\*��CeB����}�v�!�����m/��O�v��@��OAIi���_|��YxPëk��Ҷ�����E��BsE�        ���#�W���D�y�c��ǜ!}������k�F���$[��x��E;O��6���Z5��X�C۝i;���vp��A�dy�J�תmL�N�'ReF|�y�^i���������[Ց��_(   ��C�*/��jr޲���U���-�	˹�r���I��sx₶םk����׮��a!�׺�<w�2����؜�RV^�R��B�}`��4�ڶ���������i�����\�       �f�����[����貄$��)v�V�k�`_JZ�y�~~r�����yׇV �i��,�k]^QaY��Ѿ��Ⱦ3uo��A�+�v�l?Q��փ�W��Z�Yzp~ڀ���+9M   �

�{q���/�˾������~��o?��:�T�ޗGL���[`���,�H�M*\��n�b������>����$�u���Ee�;�p�ڶ��Ͷ�!����r[��0yⳭ��       �n;��<m��b�Q��G^Q�|������n���������r��ْp���ko7������g��=&�ʧE����	=���?�?�x����ܢbSі�g���f�n4Z���	  @Uy��x�O��Yoz�����O� �nL�Mm��9�W�`�m[]�U�k�l�̭gUm���^�o�#?�6��=s`O�}        �~���pX�����Lʝ��>T-ا�oo�G�<(������כ�}S�t���˪:���5ԃ6�aê������������+��A�e{˝��͟5��y��9U������N[m���˶s\   �J�/��u���}t����L/���je�`_|��ծ�-*1�
�����."TRҳk\g�p��big����/�V��;����`  �(���td���Z~X�z�J�+.����7�oʒ�9+Mn�_QQ.��[�{%�sϥJ���^{��n
s���>;>�7���g�3�   hY��m�W�%���~_�:!�
�U(ъ���[��<2k�	�z�kSe�3K�LV�K����,��Ǵ��IY0��ݼ��:�ʆ����`�o���>S�#��c�N3��Zۏ��|����R9����z�J߳�^kZ�V��{]n�  Z��92�S��<�w�����@�@��L��e��;����V���|1[���6w����ݟM:�.@S`�-heJ����|�>  �1�E�20q��W�KNN�T8&5��Lז�j�5�����WB��"��D��������_լ�筌O   ��[4:�����B����IkRRV.�&�oL�oY;�W��6J�/f�7e�c�l�?λ�n�V1\~�<���%�\F����!F^�k���;���'��	�����ir.7_6=]��� �o�!W��,��m���)A�5y��|}�>�֍���#�F�&mB��7O�kt�v��nc�*+ ��C+[+<k�h=Y���}'��:�'��~��'-�K����(t�fW�y�`�иv��1���Z�o�MPQ[�M��Z��m���&�O�>s***ڈ�+]�rlA��n_oI�nR* ��������P_s(������$	]L����ӗC}́��|�p   Z��}�H���j�5\�΃����>T-ا�5`��O����gӗ�`dSϖ���h��{�nyk�A9x־BȀ�m�Q���M+�J8��З����;��	C��k����I^۾_�؞(;RҤ��������d��^r��A�B����4Lp��>�l�&Wm��+6Z���ya�^y���jKd[Z�qް��ëGI�����_+�|����_\"   �hef���ar�A��/�t˺u��W_�>l8zJ�M�G�R�r+�Um�k0kP/s�J�o�g7�q����;V�쒘v��j�@c��򶐖��b*z�kB***~o�g��8��t�����כ5�k� �� ��}��\G����  �����h��S�&�1�ͪV��ut�<��VS������}�S���_�NQ�v�i@�����t!�@����"C��V[�S��Ɇ�ԣo���6|miٻ�6��L��1V��g��5;��	����ݭ/�p�~���oY^+�2�$-+WJ�˥]x�	�9jY��������� ���@��u���������I!��P���I�ep��ʿ����6������]5���6!F[�?&��0��WM����j�ɑ;l~���pX���ڶ�tRZ
�}  ���B��u��*:t���	���0	�CBB���XJJJ��yyyRPP`��N��Ȑr:�p_�B����S���6��I�   �XtH��ܻ�|mٵ���ݯ��^���	��Ҡߔ>]��$mU6��e�⁯U�Yņ��ə��3䎗VȐ���x�
��o|*��c��ɖf�bB�����M	��G����J����^&o�s����n:զ��L~�t�,ޑ(   5����?�"K����'��}�\��w�T����[�3���MGO���.��Kv��U���V��ǂ�����<�*�#z�������L �O󮔻^�H��߳��2*�\�}cg��5mڴ����{d�aa�RXX(�ē�744D����W趰˲-��a[��nO/�f�L+�-|� -�>  �6����;J�޽�K�.fҰTll�DEEI+'g��D������ٳg�ܹs���&�N���'O���~�s��B}���ϟ���T3>uJII��I�   ����%8���z_�;��U�8�)m#��>u�|�\����E3䊞uí<xB��SI�w�o��v���ȫw͖.��Ry��M�/�;v!S���m�ͬ����CĿu�:�ckr�<��j9�zQ   \����%&˵�=��}۵�M?^$�|�,�uH���\^W�p��+�p�����;���a}��;�������ӓْ]Xl�lx�i�{����ճ�ȞS眮�7����%*$H��#/�1K���I:�.A��wʣ�O2ժ��lv�~����F���)z�(++S|�r���1��deeY�s�+Z��<�X�n��:%=[r�JL኶_m�T���l�O:�4 ��El�i]y����S��]�.�ҽ/"������D8�RB �_�i��H||��~�ի�	I��h�J�I:����ʳf4,���/���&<u��q9v��߿�TO��S��B�����ٳ��k��+�S�C���   ���h�0D�x���vi�-��t�R/<(�T�������=Vg-�B+�\���2oh_����2�{'qv.Siy�9�������J:V}�G�������+r��ar����;6��9�Ų,!I��f�	�YeU{<�2\��?��D��K��u��뎜��¶����U��V{>������E���������}����uU��VUPRjƿ�u�i�  PW�����������p�����7�&��]�d�T�~�Y��[`�=��Oi5�>����.�ej�nr̀��7�_��^��Hs����3<�j����ŗ��7Ը����L���� ���^�t����Z��)T�����E�i~�df6n�OC}ڭ�Ӭ�%|%�X�m��_��nM��D��Wvz�V��z�����������IsR��4 ���X�>mYھ}{7n�<؄�����f�P[���q�c����*~����9t����+��K�S���   �w<���F�������e���疋7��m�S��Ps�cd�t�
3�A2�$�\��:yִ�J����j��g��2��ݭ�����))+�y���.�R�:��!ʆ<��4���wŝ�U��ǂ\փ�:i՜>��H����j._����~N��{Ϝ�<  ��x����孯ϑ�V��}��\9B�##*�������nk���&X�N��R��e�hP�Xs�#�o�'<<�n�l<zʥ��;|R&��M��SL�>(چ��^Ȕ?��fN�u�
�YEDD�+��P���-��L��ƴ�2f������ݻ-4'�  @�x;ԧa)�r6q�D9r�8д4�j����l�T���J۔)S��t��ٺu�	Qy
�)�����ܶm�<���O   ��:��/�&&��8��m&x��Hu  �$ݧ����M�ͅ#�;].���L5�O~�l�,����8�w$�I�L]�DJ���v�Mh�9�%5+O��9oNF�+�����椕!��I��0���Y�䔦�ۡ>+��aoW�k��y�r_cV*�Ķ��ޣ��HsA�  ԛ7C}!!!2t�P�:u�>\���|*$Uwi[`�g���ѣG��mǎ�z�j��Ӓ�S��5��g�m߾��	       h�K�7>���-L.F���Z�&�s�/��g7�1�>O�Jd�.d����yhe��F�K4F���R%;��+�g�Xaƪ<�-4u��d��]*�Om=�����Ew$�r�-۞�DDE5|}�Ŗmپ�F�U�,6Nд�y!ԧg��������eҤIҳg���iJ���4�ԡC�4,�!0�%&&�G}$���n������B�������P3>�z����Ǐ�����       �Q��s�7?��}�L��E&��,:����`i,A�~�UX$�y�r&+W��H�/����)gM�^x����:��V�<ߖ��C}V�3�nHG�ɨ(+�r�h�
ˇh�=X45�,�^EY��¥�^_y�e��I��|���y0ԧ�L;w�,�gϖ	&H۶m�}4尔#���6��X����HZZ�|�ᇒ����jI�)���P���?~��n�Ƨ�M�RSS�       �&AC{o�<h&�._	�Yi%;�p_cW&��p��"�  �ē�>�k����M�fE�10�Hxx�������p�=��˗/w[��%����Owb|^�JǧV�[�l�        ԛ������>w���k�T�B�  �̓�>��w�u�Ɍ3�M�6-&0U��=�ѣ�٩///�{��TH{��$%%���o��)Ƨ�9�Za��W_e|       �:р�/U��*00ȭ�ki�G�����EEEҜ��;n����gZ���� �C+T����)(��_�>�aq���wy*4�A��c��M7�$�{�6c�%����h}�����)((����g��~y�7L���h��)Ƨw1>       �;���.gB�kN�8!-ALL�	���� ���vQ���]�6x}yyy��hzz���h]\ �׸54�a�={�e	f���:���>{��y��x�	y���O>i�z�Sx���x�         �g�  5�����Ŀ��m����(���k�n���h�L��V��ܹ�	P�:uJfϞ-�G���{NΟ?_��6����9��?���;w���$�       �E��H��6�+�UXZ&[�� ��}  �)�ڿ�m�д
Z�^�L��'�ִ�����������{L�/_ޠ�hM9<��P�a���G}�E�O       ��}mx?yx���WJz���K �B�  8��P��Q�2e��r�-K[�z��VG���VG�;w���Ǜ�h��>�bx�ݡ>Ƨ{8�4�%[��         �`  ��ݡ����˼y�L�N�P���i߾}�ĉ'O<��������z��)������y��כ���e|6���Ԡ_K�         �;�  v445h�J�NB�C}�Z���={ʝw�)cǎ���2��H�޽���Ӓ��)���o���_��?��^�k
�K��U�_Q���q���o�!�V����	�       ��x��<��&��Wva� �7�  ���� 7�����ȑ#��_��t�֍Д�h8�K�.,���r뭷J�N�L��>�/���곎�{�G�w�������S[��|�ך��       x��if��`  0��������M��m۶R^^.���X	

����0a�i��OJIII����)w����g;>������⺟�H�         - �>  ��P_hh�L�6M��.S��!�B�DDD�ֲ��ɦJ�#�<"�=���y]��rg��:>��nHH�Ӌl�g\\�<�������^���뼮@�}         h�� �¹3�.�\s��q�&xCh��4�ֻwo9v옹�裏�o�[��֕/����ӟ��,T�����̔��]�u�        @3F� �̝����H�9s�,Z�H���M5"myګW/����7�)�ޗ��U�u5fx���<9����u^���y��Rq�O         h� �B��R��7�����4<��ю=Z��կ~%���u^Wc���9>����>���Ԫ�����        Uu��)}�H��hil�@�֒UX$�y�r6;O��H���礬��  |�>  Z w�����ԩS��;�4*��<����TFkժ�<������F


굮��?K��S��W_}��~��O��I�       ��{'���H�vm\�MNa��:tB�ߘ ��� hl��d�Aޢ�")..6 �(,,4Syyy��$V�۲��ǝ����`�<y�	���A����Ä��r�/�KS�������F������6����S�p       �\�G��?�x�Ą��v��r㰾f�`�Q����r1��'����C��A = O��.��4T�������O�URR"h�MiKӑ#G�Jh�!4廴j]�n��ĉ+>����/��{��p�e���$�       -�/g\!?�fl��3gHoѵ��}v�����' P�  h!��jݺ�:T��.���1�O����H�ر����ʀ��o�ŋ�k]��1>[����[n�7�|�^�"�       -�}�9��e�Ɇ��dǉ49��+YER\Z&ѡ�$C��ɸ�M��u�V���!��'W>��dZn �F� ����)իW/�?�t��U���MC�v�Lܴ�4�3g�����_|Q�u�3���`��g��S����������ܴiS��E�       Z���m��s'��������������1�l0a�d�h��]I����^iF�6;i�6MҤ	ً��3l���{/�:H��C�,Y�~�|��ҽ�}�Œ�:g���/��O��)�Uu������k��Vr�9����Ğ�뚜`��o) �k�  ݷ.���P����84���*��6����cǎ&�w����;�W=5������d۶m�z�'R1��F�G�3:,�V�����ק��>O�������O~��U~�Q�>?���       h�~7u����8��]�M�|�+))�py;�g�O��R>۲G^��|��7�_;<]��z��>��?O^�X,�Ԕ����3�  !�*�������d	2m�4BSJ��v��Uv��!����<`�~�]���7�>��S��9����4�����>�6��>��q�       ���qr~z7��g[�ʭo~&�}[l�w���b����KL�>�{��~�9��2�����= ��㏪�*%66��֧�W����?��aLL�>?B�  �D2�����}�{Ѽ�IC�N�d߾}&���P^x�	d�g�n�(�ݻ���'       �{n�OBCN���J������oh8�?�6ȏ�4���+�[&~�m-P鴩C��]�OC}���M�S�����.ܧ������ �  \ңG���K%99Y*++�-11QZ�j%���2v�XY�~�,^�XU����K.�>[����U�        �9�w��W�o4ᾦ�������g��`��X��.Y6�4=��S������C}�?�  @�4,5~�x:t(#N[�:HAA��ԭ��*7n���	4Z�:�wذa�g���O��>o��6ٴi�dgg        v:&��)��7Vnn�u�ΗŻ��^�����)���_�n�����E��  �
�~���ԩS���B�r��V�4�ٳ��4����K �ǐ��N}�@��ܽ{����ˏ�〫O       �w�Nm%������b�y�i,�{�)ؗ*o��"����:��܏W�`��g�  @��u�fBSqqq�8m����%))�tB4h��5JV�X!�"--��l����#y��9z�hY�|�        ��$'8ί;x����ή����\a���\�\��P_` �  ꔐ�`ƛ�^���\�#yu����륤�D���>�D}�\�۷7��#��>���       �������EM���_��������n�r����  ��X,ңG������J�r���Ijj�>|������
����'������믿.        $D��喔6��s�O7BH������n�ރ?��|�x	��}  �V�3f���V^^.h�Z�n-YYYr��q����/�����W���ر#���s�������u}       N�����UV���Ա�������^'�|O�n۷o��$���)+k�@hc��^;v��ǋ��  g		1�ЦL�� �۵k'{��'N��7�,�?���#�Ϟ={��ɓ�� H�	       �n��,ѵ���WVɎ���;,$�q޳�`�B-����噰�7���[��B�_��!����s�N����/F�  �A��;VbbbN���������1b�t��M���#��^�z_���(�	       �V���_,5sq�Y��d� �v�  @5���&03n�8�����m���ݻ͘�k��V}�Q�'ڭ��^ڵo׮]�>���:y�G       ��>ݼGn~}�����ңM�	��{���+MO���$!*B����x~��T�
�Stx��M����䕔�1��H�!`DGG�7����$<<\�}7[	[�՛WUU9.��ׯz�y] ���-**�nhA(..Μ�������HfR���;ʘ1c�� ����9h� ��O       @�>ٰӜ4dS\���vH�[Fh�u���o���dx�v�?��$��:Q���&S�w�!�R%>*��=y���1��j���r3!?����"�B媡}e�m�S���$.2��uN����%�e��#���!`���9�[�]���w�'c�W� �'f�W�?�!?�W �K��Ν;�ȑ#��ڴi#���)�_~����`��Q�FQ�A̹>g̘!�?��        ��B}�ܾ]�)h�B��ult��{���!���~xh����Μn7Pny}�l���4徠A�箚���u�1���s�z��ǋ�ʏ�*�0�C_���3����kdd�	i�O� |+55U�j�b����SBB�鈗��cBt:���ѣ�}�$%%E�B}9������'        ����	)m���v�K��X�yN~���l8t\���c�w��=;��}۵�9w̐�Ov���x�/�iPo���H�d�����"ӹ�k�x�ث��O�3����IEe��f�b�W� 4�:����v󋈈0'�i�O�,ҕ	�ëA.F�B��<xP���e�����K/5�]2cxG�M}<8�W�	       @c\��l�{"ףul?�-/-� 3Wo����3�?�[y��i�&.�t,{���r�����\g��x�/䗖���Α��IvQI�׉������'6�w�=D^Z����������v_�w`�N~��OC~�UC�=�5ޓ��(}��5]��ǟ#8%%%ɑ#G$++K�L�"���z�@��Q�p��p��a��O       @�q�GA w���4��>�/ێeI}o�/�sXnzm�̽c�Y�.~�S[�@ �R���cB}�*+嗟,�]�˰.m%�b���䟋׋?"��/i����"s�N~����E:�Rǜ�Ai�T��8q���رce����v�O8��lժ�dff�E}       ��ӂ=��5#˥�i3u�ޮ�Y�)U�!i��ͻM�OuH�E���� ��4�g��;�� ��hu�i�~�د�кuk�Ӯh�~���O�&99���>/���}        4�PN�#�!@���:���XA��+�} ���JJJ�)**��ЄRRRd��fvUU� J��z���7cp۶m+>��'jc�[�^�����ѣ       @ J�����*)(-��6��It�����0��/������7�E�@@r���Ę�~�Ӡ �ip����dqǫa���\?~�����>��'꒘�(��Ŏ�|��       �@��U���.m%:�d����R��?*�7��Vlj�p��.�G�$s��j�o���<�}!<4D~7u�����,�;xL��yP��> M�}eee��R�� �EDD�NW]�ve����}&L�y���D}j�'�>       @�ףc�娰P۽�9�;y��������m�b��q��O6��������������/|oP/I��4�S⢥cR��۷�t�}Uک��Wf����"� ��XƢ�"����5c�JKK���u�֒��.@m4X��U=�j��z�)���Ԭ����ˑ#G       �@�5#Kvϖ�9RTVn�G�w��:뵱-������W�ȼM���;��M���of-����/�ts_����wj�3.?��/���D>�n��W�w��`�C�����Idd�y�_G6j�@�����W�^�9E����͸���|>|�̞=�gۦ>ѐ��G}:T�̙#        ��w�l�?\(;�g��=�7}@yj�df
�]��5�����+�E%no뼾]�i��ymLv����`N� ���}aZ������^{�~�U�jľ`����|�DI����?n�G�@�b�qu<��k���3�y�{�՟��@3
		�V�Z�1�t�D]4�w��1�2d�ς}�'\���gdd��6l�>       �ߛ�jK��ӷ�g}�Kve�ȗw^%1�f��m�ɟ?_��v&��$��<MBC,f��-�O7��_4�/��xz_��������}aʳoK��d�G����)I&4{���#�c��-=l�����W� �H��)77Wbbb�y���)11Q�u�f�Y��u�cihh��Yg�%���&@�m�'\�\�	       �7m>rB���:�o��|Az7��}����[߿X��OF���T��d� �f�ѓ�����.��ھ�_r��EA}$�@��yP��b�||��&����e��O6�D�@�VTTdF������7���48���F74��b�Hll�鈦P{��-�6m��v�O�¹>�V���#7n        �v����o���ui+���R��L=��Jy��U*�����v������/?^(/]�Y�s�P�} �\�˓��̛�t}N���S�N�� HkpJ������$�G}�U5�`       �%8���8j�z���7��1E���ea��_�F�4o� ���!���~hP���J�CCdh�*e~8�`����}�?>>^����h^�:3�jp�cǎ�� 툦��)o�>�_�'�O��t���2�[�
 �y����m��x��q���k�����%,$D     ���3��������w���Z������k'�o�L��#����of- �ٻO*W����VT�``��(	������fc����Idd�����C���������n�O�b�MK�0�ڵ���p:Y�A���&lW\\���	w��>\��3p�L��E ���2\n���|�n��=�[�˜�̐.�	    h>���w�	�yB?llw8�@*��n^�;��||���ul�Y����̸Q�%���q��m_��1HBT�$�
�j���R�G� ��WPP`#�p���_TU�DW����,m��i�U�S�pEHH�#���֭[ˉ'��=��p�O��ۦM����)�h�@B} ����x������}��/,���\6�P    ���&5_	�5���s�P����n�6I���Kj|�Y~m�&������,h	̾0�y_8��:��n����3L@D�@б��bbb̛���F����2�.�c��������`�	wլO�}h*S�u h.:Nv\�N2g�.�ktt�y}�    ������é9�WX�u�5�篚":�1�:����^�kr�̺�{�.!�,�\�E�y���kժ�����+뎍��I�eHNN�����m_8�C�Yֺ�ג��|_7"]>Z�S������}���/�X�}�_�������>����
AG;Wjp�ڇ��x�4���իW{m[�'�U�>W�Z%       ��G�������o�*_n�+��<(��򤠴܌m-c�u�������h�m��h��?t����~�43�X�TT��<9���"۶?X�]��6��`���%//Wrss���t`�z��������ҫ�߬�uk�~u�hy쒳e��=�r�9��o֧��:&ƙ��}��잝�Y���p��j�c||�c|L��T	N�Uz�TeeeҩS'�&����>;v�(@S� ����1 �RPZ&Kvy>Z$�TVY勭{�'�    ��p_uQa�2}@s���;�o���%�FU[�#��t4���>��k�ޖ��h���Hs����Hnn�>^;w��/]/��U�1$1:R��ל���}����ד��> AO��LHH0��������`kyy� ����0_�IEJJ�׶C}�1����W�O��4���l�)}����] |���R�z�k�)�y��~��Bо�tIN    ���p_YE�<��2	f_o�'�RZ�1��!�^����t1{~�ZY��_�����O���\�>_?^�G���}�}��Jme��6ž��W+���i2�{GI����:�[�琼��;�h��w� =����'���&@��@��Z��\��j۶�׶c�O�t�*_�'�OiE�\��咁=et��Ӄ �mG�
彵�d�q���t��1+c�x�|2�o�d	�y    �Dϔ��_���5��}o��jN�|�s�xI���ֱђ)�%er4�@6�4�M�b�ïHK�됛]s������C��m�~�v��,�hN!�tk�()���H����S�+��GOHQY�dB�������������ҵ�@eN1�����P�֎}�
���p�s}�iӆ�2�T���K��^ |z p��1~i�    �Nh�E�~�yru#05��cy+��dω\s�I��}s6��p��}꫰[s���4qrq�4����5�]�9����)�+,,���X)))!��MG����Q�p���O0���	GS�>�X������Q�       ����;��o(ܧcyU���pZs���|���_�����;܇�� '�@��JKKh���Utt4�)�MkG����?�=�mP�h���y��       ��>4��������K�����k�����L���ᗘ�ܥ��***Oj������       ԏpܡ�w��}yo��௏W�}4��?� ���J�:�W�UUU��
�|d�X�=]_��L���_"##��n		1_����r���Dc��>       #�W�{��~�l'**�I߯
�����Zh ����t�+..�`�!<��[OMȳ��K�/��V�;4�t?�VQ�h,_�'       �5��А`{�����p�v@�;���d$/Z"N�;[�p�o��O4�/�    �!�u�X,۬V�&�����5$��vyveEUQ��Rj����KeU��]�"}l��m�X��XR  �} �x�� �(--���h�}hq��Uhh� �wD��^�����E}    �c�Z�ٞ�}f�ZT���/z�G=Y_��O����L��c[�b{&�$  �����!� �Б�f����Z
�<�S�j��ܵ�>�)o�'    �a�����O$$䵼'����L�ɞ�<�-�/zzA�|&2)Bη��F�V/�m'\  �_"� �#� Ю}:�W��@K��L'J4��8��)=>zk:p�/�    P7��g{V��k�������wyo���]�#2�vnV�=O���v�v�X�  �w�}:�巄� 1�} � �����H)..�%���c+WكSv�f���)ù>�    >��"ևr�ߔ�V��w���{�ؾ<����l)���*��Y,+  �����T�>�} ��> p�v�������P3�tZ�tDCc�"ا�I����    8���U�e)�U�����'l_~�����QQY�g�Xn  �W��k���4A�>��N���|�M볢�B wi�(�}    �}V�.��ȏ��zώ\�?'�z�aۗ����[�ˋ��  ��> h�> p]�Вhh�`�ѨO4�    ��V��sy����]�s�O�37����W�f[�H  �߰���BCd����^W�}=R��X~��ye�Ȭ�v����w� 7h�$<<�`��raa!�N�6{�.,,L���������n�E}   @P�Z��%���'��Z������=����#"�P  ~A�}����~t@�R������g����Y,�.X# ��` �A����ƚ��}����Unn.�)��>"WCS:�Wá�@}��4ا��5��P    @ӱ��J��Oܹ]�Ś���%��g�VYe�E$Z  �_�p�m3?3�
��?�[8��h�|�e�l������� 7h�E��ih�1�M'6�*U�|L�1�*/>��o�R�%F�>e���4ԧ�A�\z��ګS�h�w��	 �ԽM��R�u�**%��Ld�ɾ�<��.�{w�)}�J��8I���]fF��/����g���w����Ǡ��n���R�b��:��1;vGsd��#.o{R�Βe���~N_m�W���c�eB�N�y�vKiř��_���;5�����
K���)~�hX+[ML�Ն�E;�:wWz��ҧm�����|Y������'#��;��o�/�ťnߗ�����v���0�V��q��8�i�WVUɬ�v�7����~�dp�Ts�im�'*�X~��+��,���1?�����&��,#���6���#$��TrKJe��l3Rj��ò�D�x�t�vo�!u}�tt��.!��e��d��c�.o�f�~�~� �����0kŅYO�wH\����8�g�L��X?�X,�  ���b�������` �I������P��T_�/Z*%�z��;�j���F��:ՠ�*�Z�48u���o滋�Dc��>�����U�r�D����X�m�#/-� ��r֠���)��9K���Lw��������9�ǹK\
����N�����Ͽ�r8���L��N6C��K��7n�.���f��;���Jm%��8U<����҂3?�t�оr�9�\^ONq�|�i���l�|��� #�sӨ���i�]��y�䉯V����{��玨v���=���}�BC}�u8��7d��l\���.���L���v���K**��/^�������ޭύ#�KEU���z���k|���E.�K��������t�Ys C�Y�M^[�I�ʚ���_ێ���B����Ԟ��c�� �m<�)g?5S�\�*q��^p��$�}p����Y*���z�i!r��{a�=ϝk���vx�  ��@u� �M��:K���HUU� �H�Z�ʼ�<���c�4\b4GDDx�#����U}�?ӮO7��'׍H��Y'����brQ����kΓ�Sݹ\�3%I^�y�,�q@nymn��%��7�ף�K�>�r
��n��cR���o���:�:B}�~���C�;�fx�\=,]^]�Q�h��W򼳩]?����~���+�)���Nw�L.��D|E����;�q���c�/>Z(�B��������z�|����;�l`/���2s����?��n��� am�vnkN�M!�|��g�w�/th#��%�Щ��+BB�=yw�	���=}�ğ=s�X��D,��!  ��p_����[�
 �!� nr�k�"w���-������1��)���e}@s�ў:��YdX�tk�dFp�iW�;�b4���u��y� yr�9ft�������N�l�^�+(-���9�C�t`O3�NG�ιc�����uv��v,K���qrܤvs�3ڐNm�c�IGW��B�g|��e�w5�;�_$�s�].���y�tVt&i�	ҧmk���5��� �ar���Mgd���;����h��idٞ�M����2[O:̹����쪡}����:*�גc���^b�x:[�|�n��4�a�yi�wH�7]�����ԱC����<b~~�����"'��m���dվ�f��*,���(��b$�]�\�ޭ��[=��t�P�
��_]0Z>ް�0�%�j����S���ܧp�ӷX��X�`  ���?}�F�90��.�} ��(**�`��:=z������}.).>�&ttt������=OP�p�s}�ܹS �%ҐP]]���M6c{5hgw�������^m��!O_1�Z��[�7����ce�E�Ż�?l�aJ���v�[��Z׿}y�G�ʹϾmFv֤/�.�}�tԨ��M7��B(�#E��K���ۛ`�ܕ`�v��**�-GO4x}����X���ϖ���&I�dB�Q���kF��߾_�4���8 ;�tI���0��񲩂}��a���#�拷i����}˛���~�O���0�֔���v�{�W�i���-�k���1��q��a����1�㱃̱JO_<޶O˛+>���w~pI��{O�ʟ?_!��f�,��nkX�vr�������-��Y��2�
����j��yO��� ���1��x��m{�/  �{�oWf�����}�E?��� x�> h��g�Xǋ����#G��Z\QTTd�j����)���"##�< �����H޸ez�`����5��!1N��jJ�P��_|k�g�j�>9��we�3�xK�� ���:CL:���Ӏ��N��r_���9�}a�Z���q*�{u��h�1�,���.��3s�Wf�q���Sz븁�����.t�Ӄ9�%ĘP��Q�~�P
K���k{x�Q�Mg�='rś4���T�U������S�~�n�=���=x��j�������t��/)�?\({O���߾7IV�Ϩ�3D\d��n۟�C}�/���\�ކ�!C;���O�y	�ԌsL��h���Γ�v'���}s�))���X-���=q�W$r����j��b�   �oh��1^� ���` 4REE�x���)��c��[iFF�zw��	wh}��Z�Ǐ7� �H_���rn߮&ئ�t�hF��{hH�y,�v|ԍ�5�s�K��{�3�W?{��.��#g\��]�-kh��`�	�u;�r�>�lP/��^�$'�����:o?�c���re�?���/?^$���p�.���dF%��Y��p�s]�c�W�j�i L�}o����m�~��.15��~u�h����7]?���DW��A�6y��LGڶO�3�ms�j�_�2±\QU%W�<��P���/Zk�%�qF��'.�du�`s���c���s�>i��Z=�\a;�]د��=V�i�2y���Ͳ������_-@��Z�̋�zT���X��3�UV�Z�R    ?@� I������C���V������T�V�(D�|9�׾=�O�J}�^����td��A�w�
5]����j�G�Kvy%e�O�����s�8�?L��s����9�[3Nȉ�bim�uL���PuJ1ݶ�ѼB�q<یHu������z�}�c|Ւ 	�)���w��@��4�y��xd��� �v{ӟ���l�Q��}�F�u<	�iX��n6��Ռ��M�j��L�%<ͩ��;k��Ns3Wmq�4z���׫�9�([�v�Z�^6:��z~?g�L���щPC�C;��52θ�?~<n�cYǄ���g�
����uަ��/����Gv=y\��a���[\*�'l�^l���M��ǠS�����{�A��   �����i�T�=�@@� I��?����	��+Z�.]�c��>�ח�){}v�ܙ�D��@u:���S�0��ͣ��Nbvo��"����/�`:qٻ�]Կ�tno�i������g� ����t4��]�qëct�_5�����I�\�����|���R�t�;�*o�,(r�TR4�>O��N����1���j�jmjw�_�?�,�J� =S�Lp����ŷrͰ���e��"��p�\��,�+��1^��E�}j��l3Fvx��������U��?�#m�����i�E�����2�����G�0�v��m��g\W�z��p�v��Dn�]&�r�9�*&J�8T�t� ��#�O��?)V�}��W�{�f�X&
   �.""¼���t��*���m����㭪�4��p�� � ��!=�H�����\ٿ������P�b���Tll�lڴ�'۴�g׮]�O��<��ܼ��v �����\Q����^��-kg��*,-7c|�?�dw21�ݳs�ϖ�:��i7-�[[�-���;�[��G������$u��������v�� ��@�S I��狽������ڵ��u���}���2���u#��Cs�6z[:��_K6�]�����u��i�e��#�Ԯw
ͭ�Č�{k�VG�O��jhQ�#_�)����E;ʡ�|i�7mǖ�N�7>�w�Z�W�8��
�<��Ŷ��W��ɔ>]��g����F���ʶ�r��5�5��ٻ��*��  �/t��I<�wa7�i���)}��y(**l���� <����H�}T999f��I�����􉋎///�;v�d����8�ɣn����o߾]  ��m�\m9��t�7���ֱ�������l���`�۽C���Ż����q���j��ctud�v��@`��x3:��\ڧT��ܮ�ӱ�}ڞ����BA�i����eBe:u@ܗ�'������N�:���O�� ic=��J�iTG�8Y}��ISJo�ڶ?�:���3/>r��5Oi�<_�F;��J���Ε:Z��)f�m|�	-�r
4j8�y�e���
�:����]L��D���玐?\(@cX�����ς~�s�Sw�O��7m���   >�oa7{��[����C}�?� ��`�������RXXhZ?3������Tbb��]��g��>�c�vc�����8���ի�� �Jk/�RN�p�.*�ݙ��o=S�c;Ն��=�f��F`fP��Z����	st\�Ү|�.Xs��4��p�×�x��r|O��j�O��ݾ�`߸�-ۃ��H��0#[ݑW\*Y���T<����`��� �h�6�����:{c�G��}b�L��E�غ�����/,\#��p�Y֠���i�����T48h���U� ��o�n�#��i��7�����&��+�;������1�׹j_�#اuJ���/)q�G�뱧���~ s��L�x�N��U��`���&�
�igށ�M�@`UV�c�b�A,"   �		��8Z}��������o� ��0�4(���%�w�~���}�Ҁ�JHH0�)_q����t��j�� �1)^^���j�}�yO���=TgwЃ���ud�m���s�U���:�����w7�ڕO������� �s�M���>a�9?�g'y��3�k�w��v����	o5����o��/?^$��q��O!���L�aO|�R��F�W�o����v�q��6��/�(���fYG�z�S/,Z'?7�t�S��h�|i[gS����W��X�b��Z�:f���Ǧ��\�����j]m�@���dW���q̩����[:�0���5�����G��o}!�[��G�ݫx�}J��wmM���,b�B   �3�v�u�-�/�G� <���Y,s��Uvv��ܹS@p
����碣�M�>_���ѿ����>Q��O �5���4bVE��IZr����&?;��Z����/����^r�=���!%Kٷ�U�u�:��iW>�U�������_}l����f'��̧4\�<�W����SmjwM*W�[�2�tn/û�����/��W�-�͕�y���	�g���X��f%��mM��n��]���T[�j-{ҍ���\��j�����f��6��������Ҥ�SW�ں*�/��S��G��i���}�N��ʩqܪX�y��sq���]Я[���0��Gş�<�c~��.�W�+O/X#[���%V�܂�7�X��'lZ�  ��
�5W�-�/�C� <��>�}d�`5��蓈��R���3��rrrė�O��^�����g���' �ڳWN1'W�?�w��U��*:<��rY����=�fv�u%����|��>̫�>F7��X�˒>m�͸Ԟ)I&�bׯ}�j!���O��
56d徣r�����6���һ����l�����싴�檡}����=����6�g�.�	f�W��O��)�U�W;
�i@W�s֦��J�[���5:���h�tƱ�[�ê���B<U\#�Ys�vV��65(��S���(W��_�>���W�U���z�n���:F�{e� ��������6����Oݽ<��g��E�   |��a���������4lb������\�9b�Sݻw��Q��TRR����;>߾�>w��%ݺu�>Q��>[�j%����?hHGG��M1���t��]�~U�њ���"#�)8w
�/-�s��#�&�d��v�{a�鎫����m�Da�l�8����݇M��ܾG�j�>�nj�.��}�.X#���X����r��5�F�w��}���X����7c��M�x��Ι�}�B�q�yfYCu�{u��F�SG��۷�c���;������Vnv����u#��O�/��r�р�'kt�����rS���a[}��d��t�P���QGvm/��;"@C,byMP+�X߰�|   ����n�r���� i�D;���رc�a��ի�)T��)/kG�E��'�c�Ϟ={R����g��6Yn=���N��+z '�t��t����.&�MNQ��K̀Lchg3�YY�u�vt,��ӽ�ԸK�����o��x]�Ֆ\��|� s~B�N�R�ztr��@цC�����n�Ni�s뚜 cm?��S�ei��;����;G>߲W�x��qH�T��[���:U����l�{'w�^/���;k��ݓ�J�v�����i�Km#�]q��t	��tz�ۤ>������3e@�6f�Z���l�O�T��%Fy~̩9j��q-������]k�Wz�K?���wO}�Zn5@�O�@���1r�Pۑ`Sޓw���b	���D�  ��h�m���RTT��GEEIii��o?���H)++�} �!{�> ��8qB�l�"%%%��S�SAڭoժU����,�C�s���r�EQ�pp��իWK^^� @K�]�>ٰ��e��ԍq��
��(�+������=��h~�/<�x]{�O:ڥ�ޝn�S�oI�����wv�׎}�9+��@�������{��1��dަ�&�X������Jld���#A'?�l��4�N�j����[��8�}J��m8�У���?}�\޸e�Y�1ҷ�h����<�wV�	�6�M��z��	�|�����E����gS�ȯ��wj+Y�x�o�cN^A���5:vk���z��ʤ��:�rۮ���������//m�5�<����z�~�d�Ou�}�=��=����F_  @����w���u���[��Bş���Ik�����#� ��Q4���ѣGMxj����3�<�����o��{}nڴI�B}��� _**+?�����e�1�m��rﶭL׸�FvSû����ro�c����.}��`ޘn��y�w�V�Q����L�;I�;5Y�edI߶��ul�����Wڝ�Wg�?�LBC,.��8U�~j��$�����UC�g0�����jh3�ٝ mm�l�eF��hTu��ڊMn�ӣ�ڛp�]�~��׻ܾ?�E�o���A�np�Tywm����z������2�}_�m��{�$��㏵;inqpt$x~�Z��؁�j;>��]4V���/|>
u�Z,�џ�>    >G <D�(�:�tݺu2l�0�S05��
���rY��q�D��}���éO���~BO볢���� �>}�p�E���e�9�OW��qW��i_���::���XӼ�2I85*r\����7�̨K{0/��Č�˲݇L�Oi�?�Mpë�3`�Y�〼��;��؁fY&z����sAz7G���b�d���?Z�yg���-�On�ܜ�n��7q�<��2��q}�.����m��eyw�ЊA�����׳�i����"����ێe��rM���;�ͳ��
K�婯W�c��m�5Ly��^MR�h��R^nm�N,�2_,�    #� M���NC2۶m�H���Mp�+++��@۶meΜ9&<՜�>�n�J}�����LMM�ٳg7{}@��t�ja�F�kt�O�u��tq,痔��:��X��{�ѳJ;��S���O�4�SUχ�t�5���y�����Uë�O�}6�G?].3�6�2��y#e�-wk6Z�M����$�h�A��}����0X��d�˷�.���K�BdX�\9���s���o��ǲdω\�8\�68:����?sV���z��9y���%ا^^�����!��/-��k|�-��_ڍY�ݝ'�WyH�7�V>d   ������c�>��e˖ɕW^Ip*��q-33SBCC%&&F�͛'��������@�Κm�i�L�.���&��$��ttퟦ����C�]�ф��d�!G�O�Հ�]C����9�}��}Ў\v�����A��k���5����!��g��������X~k�V�}��n�����u�5��!1N�x|���T&��b¬���rߔ&��K���S�.Տ��T�[���m�~���?�v	�fY�o��i>�_�mػ�);��=�_��r��t�rYee��_��{O�Jک@����v�[w00����я}�B^��\��+��\;<]��,�A����ӣ	�=�c;t'	    ��>  �]�֯_/�'O���DFM���3~W��}�嗒��/���������ꫯ��>q���0y�����U[��@�J�+L���a�5`�����yϽ#�nt�ӎy4r^�߸����잝��4��y<G����RJ\����1.����k�z���!���?�0،+���Ԗ��a}͘i���ns{��nc���XL(ꉯVz|��8&�|�S.=��|� 9����37�8�Ү�s7�qk������M'75�c�9�xlo���ͦ���뷍$/.v�[�߯>O"BC���j�9�F;�j@���e��x��2������\��[���]��J���f�珔�1���� ��E��m�)    �C� �CK��hW��˗˴i�Lx�G��i'�V�Z�'�|"��������9k�,	4����[/3���_g4�M��ȓ�x�K�̛ҁJG��2z���Y��(�>����[�>����km�u<�?�Lf��#�F�j��+�T��׳���.��<.��\ܩc�/4��4\��H�A#�rfK���Ϯ����_��ѵO���9i��q�RAÜG�f����^�7�:£'י.O~�R��%�G>]f��z��5�v�a�F;ύsW=g��F��[���S���ph�x�v��������:.{�ҳ���B^�vS���P���O7���g��og/��v���d�#��3�}�&˧�w�\��&������G>[.��t�Y��a�f�*p�E[��   �S� �C��EKs��1Y�j�L�8Q�������<)..���dY�t��b��I�&Idd$�d�;��>u,�ѣG���>E��s~�_^3� �J**��o~&���J�Qú���� ���X>\���Q�r�����������v�.�������{�8ƥ��J{����>��9�^�NkdHc$FG8Fw�#��ĭn���ٵ��q��EkMPuٵ��C��Z�zs�֠�V�%��m�dtZ����g��l��j��#�=�Z�놧W��ӅPi�@���g��i�W�c�y�Z�lc�Fj'O���g�z�.r���fY�?w�s�Ü%��D���࣎���gK���奧�_�s�{�鵹��W�P����>x�m��`F����nh��FK����Ns<�ǡ\�5���P�j��j= �   ��� �j���dϞ=�`��>}:]тLFF����H�֭塇�\�t�>����Duy%er�S3=^�{6Δ���@���Ŏ1����u��ߛ$��C9���~@�62�K;�q���r�;_��}�g�ռ�KwמE�v��ZC���y� sr�Cs�ʓ_���T�k_ld��=iX�]ʂ��#�w$kl N�8^{�Oi(�)�}�ϟ��+����������uNcxO�׶����q���Q�|rL�L�����]x���f������������Wʏ�t\�#�����1Y��-�؈pi�'{u>#��a��_�#+\��{$�@�}�]y����Ki��{'7'Yj�-��3�N�ᡡg�k:j�ә��h�����sPz|���	P��ҵV��ŒO�   ����&@�(�4��q�#F��6mژ0Z���l��m۶2o�<9r�?G_j}j���ÇS�AĹ>?��S��O�Ve��ho-�w �����;���er�.�˓�#�S����5���Jyv��F�']��[�״��	�)�ULT�����f׾�(�/\#�E�3E����z;�u\�}���a��ٝ��wi 큏�Х�tl��K7�gi�p�t���h��F�W�s�O�8���}ME� >�����f�*������h��������ۻC�}�������1f�:��1�zj�v��`��]0���.�q@�NZG@MV	!��2k���    �;�  �4��k�.��/��o���2A˦�8�fF0��������_�7�@}�@�O D�����}$�zu��'6���KMڝ��.yf�j��j�=�a�_�G+n8tܥ�k�x��æۘ�o\��]���r����ˏ	Τ������{붋���{w�v��y#�y효����fi
���Q�M���G�ڽ�AB��xu$��'�t��yG|X{y�w�1��ġr��w�<:�&��c�u��썻�M]�v�� ��.�7��m]�TM�m>rc��������-�/{^�Q����XI�fb�3��v   �5�} �!	H�>�D�kݺu2f�IKK�+Zw��q3ֶcǎ&4UP�߯�k}�]���g׮]���f}���T@p������+��IO:tDZ{�/mb�%.2܌�<�_$��d�PPSЎc~���q�+�=����V�E�{��O}�ʜа�Vo5����g�ͩ.�̜C���~�b�����>5��t�3o������)ޔWR���vMN��:��Q�m�M����g��W(��1�ME���y��I�����t�L������4���t{���M���\���X���Y�ގv�l����u\ֈ0➮�O���   �[� �C��`Z�ݻw��}��z�����Tff�鄦�N�̙#�@����?�>[8��,))��s�
 ��J**囝-g�- ��]C��k��t��YXei��%U!�b}    |�` x�`Z���"Y�f�,^�X&L� ���СC��]�����3�j֧�     �����s�U�d    #� �`_ee� -Ձ��>�>}�H�6my�����H^^��������eӦMH�ϖ͹>,Xp�ِq=:J~IY��z�$9ΏLk/����]���|ٝ�4#1   �%4^�����
   ��� ����%
-�v�ܺu�|��'���P�r�����i�_�u	4�g�U�>_{�5ii^�yZ������5��'�Z)��L���v���RYEGc   ��UUJ'�k�֎b�e    �"� Ҏ}t�BKWXX(�W��~���رc	��:�T�]�t��\���%��3==]ƍG}����ڵk@�g0�,(6'O�m�,Q�ar ;_N��   �^Uo�k,�G    ����4�G��b�޽����˿��oY�l�dee	�Yg�%3f̐��dٳg��]�V���/� /����Ԭ�5k�HK�+3G�0gI����}G���0��<|��-.�A��z��;$�ɭ�����D�u4�{�Ʃҷ]k��;_����,    �����ˬb�M�>    �F� <�cx	�!����Hjj�:T-Z$eee��ӦM�>}�����.������%�>[��Z�v��������%�����:��.!V�9g�9��ܥbF�   ��j��s���,��$    #� �Ё�ʛ�Z��	M�7�Z�b�@���������|�2e�<���-ft-����)�&M��{L�    �a�X�J�����g~�#�Sxe�8	�_    �#� �`����r���5�^�z�����AG�_r�%���b�o���dddHKB}�����k����    �b	�
��3�u�)    ̀` x@�}������"S��{����B9t���i�HZZ��^�Z֬Y#-����>�J�։�)�Er$�@    �1,9G���j�,4�   ��@#�����UUU���|	�A�� Uvv��i`��ϖ��d)..�ٳ[�k���YRR"'N���`���=:��n�f�y쿒]TR��Q�a��G���-X#'
�k]�#�L���w�'�Z)��L    �1,b�j�r��V��=�M��G   �l���>}��'Yll�yɟ��E��@#i7���J����t��#dɒ%�;��v@���$::Z:u�$�=��{}6���c��ٹsgy��G�%���Hs���Qa�r�9����}���`    4��������ݫg�Z�n�Xh�  �\��CRR�9yoy���#����@Z�jeNޒ��+�����@� ),,L***fV�U233%%%EF�-˖-3���?���� �����;��	ABpww/R�n�[*m���֍��z�P�P�hq�$X�"����/�af�$W�ӽ;73�!g�w���=o�ܹdggGaaaB4��Qn��G��au���@^N���`GEť�rf6���Z��0�ʈn�X�g���0�0�,@�WTt�睜�]�L�gd4�������︸��W�"fd���}�0��}�0Z⩔�����>}��[8�___�?>988PϞ=���_o�����)_|||4�>�Q&�=]�!4"$H�W����]J�5����v�삛?w3��;�C ��13Zm�2�0�ѕ�ͥ�^z�^y�o�F8?�A?*#.��0�0��ف�m������ӳ�i:�Jԧ���E<6����D}z f,�?,�c����Q�]���3ʞB<�w�^�63M�~�����$JѾ�����͒��>�����	Q��ۧ����(؄����ɰ��K�
ik+Kb9�
lύ�KF�$+���k�����ذ��⍴��yRZ��a�a4�N���qkѷ��(�x��a���BG�Z�S�@
��V�.�hkM.v6TRV&���t~>5�N%�Ҏ�	-=jKKr�)�&dK�K1��);+K��M��N�.���4���Mj��[FѨ� �,�����J�.���h/�Y)Y���#�y����i.q_S����ũ���1��.��0U())18�0@����i�вeK���[� �k׮��oj�Xp��U�'���P'��>��վ�г��(����{t5��I���T:��NydeiAn����� `�p����1�X��~;CJ�!�>�d#-9M�0�(���饗~�W^�IO	��>�He4�t�0s�<9�'��#T���0����4�|G��臘�m3":��sF�������I�@�6�s[�6��l)����.%ӟ��RrV��1ǆ��gG��-�D'�\%���h�p��+*��R���I:x1��$�=0(���K�N��c�`߅+���;h��Db����=6�MoG�nΕ^�N�F�8E_�<B�E��-l.Q����i-^��a����<��e���2))I8���S�2MGpp0͝;Wt�۵k'DS\޴n��O��	�isd�1�ԕ��:Dn�%%��߇諝G(�̄~G_O�t7+"D88�7}�>wY1%[�����ۢ���k�ӆҮ�	�%j�aFA�tm]��gf-&�,�,��,�a�
������G���M�~���;}0c8��?�n�~���B
97�ooKm��*=[�N��ā�ΦH���Cf+P����l�I�`��ɬ�4�W�J�n@w��L/��%�?��R���+�π�o��{h&���_���ib��I��n)���~���1Ű���m�������p}e� ��w����x-������i*����e���aꈕ��p~�2�c}�SOOO�ׯEFFRz:w��N�:Ѵi����]|���^1����|�������E����ۧzAV�w{�7��IN#�iN0����be�f~���Y %����/���B�L*|�ޓ�\���Ny��~n!�]E��%T�;���o���a�a���H���h%�rg>i�'>/++��n}�TeNώ��-���I��_�"\�P�33���r�`cM.����L!>ԯuKjY�x��I��M�?ZBq��4?�[�ӊ{�Vr�3e�_�0��"6�YV2/��w��O����_�0�\H�VR�Ջ��g<z9��_� G{��'�,,�˹���@L�5�O��E��&�G��;S�I���::�L���������{��N"[��]P(�9�Yzp>��o|�W�zS ����p��YkHr���O~���a��X[[�_5.��'6Q�P��F;�<�%1�D/�B'���t��Q���'�� 'Q8Ѝ1B�9MMM�O>���p�lZL�Ϗ?����.l�F�S@EY�ǖm�Q�g�׻��}L�ό�@/���leLj�Ȑ 1i[��FQ�1����W�?^�a�a*��%+��L��H����,>�L����0�� ��iC��UG��7F֩�*~�]�=�?�
�%;Q�v��e�4/5}5o�Aԗ_\B�G�������Ԇڵ(w�C��5̠i_�0�l/w�=]�ѡ�?/���������|��қ�Ӈ|]龁�R���9t��k*�܅3��[F
�8����6���$7p�!� �ϰ�R�Z%�?��i�!���M���ıA.tW�����n�x����wn6r��qvv�)�+�x��>F^���a�XH�l�ż8՘��Ⱦ�ף�<)�ڛ呙�)�lv�֍\]]��ɓBT�4p�<y2u��U8�mݺU��15������zZ����mc\�ʸ`Ҭ��t�4Ξd��2<$P<���J�����c�tnώ��I�@�_G��Gd�/;S���ǋ�Y�@_�y����0�(t��\���#���G������0S��t�-��yk�>��L=�8Oc.�E��e}��׹��\{� ����L��ס��ri��EU
=/��I�"B�I����A8.�}h&M�bŧg�Ҙ�#T���v�Ta �R2���;��K�;�!K����ѼEҡKI�>'5'�n�~-�X0W�R�ߏR�jfX�@���%���9Yj�.&Vzυk���?w
�n� Ā���D���+��7܊dl�cccK���㵳��2���>�a�:`cc#n�|3c�ړ��/��Z�nM���t��a!�bʙΜ9�����K�.�h�"�|��.B�ϛ	�Ϛ5��>���;JH�������Ĝj_��i�0L�ӣ��x\y�4�gp>5����I��-[�^�g��H#��߂�}�0�0tD�e��Ь�F���%�!<��(����\��aS)O�:w5���ذ�U��,�J��Z�/8��M��ƤA�А�
���3�?�ts%Q����C1��L<��	"�����x&M�|�+	Jʵ��~���������u*�Q�|�;�3�� ��>v��
�x��.�=�������^O��&%0�c�a���n����H,���A$n�����؋7�o�ں{��:��>�a�Z�R�p���!�a��������AC�⩔�b�Oxx8M�0������Ǉ�}�]*(( ����'�h�>n�L]�vv�`W**-��W3(=��#��v�M`׆#	�B�֮�;ɝƍ׍�a�Q:�siu��L�WH+���Uq6����<�a�nN�Nf�� ʸ��G'�\��|��Չ��{�[_\j�?y���P�t�����;&Ш� �]8Ӛg��3)��%e�IsZn����7~�]��˸</\��&����C"f�T�9��]��5���}�kLj�-*��VRZ*ڇR	�o!��8�9V���<)�}�߽��>�a���}�0�n}(��*z��8wRSS����z��M�O��Su��֖Ə/�S!!!�s�NZ�d	1��}��y�������YG���]�vq����l���X��Lr�i�,tT"�CY��]0C}<�S���v�Di����1���;(69�Ԇ��#�kM�.b��M��Oq3��ҹ�DvJV^�?6�٨ܶ�o���e�a�<:������we���&� �Y�KA$�a3XVL\4�����T<b�i^<������ߋ2��~�'-�m���tu�?�AS�\A1U��䊓��x�O7�6�`Tb8�W����(nv$7 �D)�����C��ў>�9�fw�Je����6��_sբ�����-*��a��1����Y[[Snn�l��1�#�?m۶-����ѣG)=]���Ơ}��4q�D�֪U+���o��5eL(}�lӦ����}֞����!�e*���Ǘm!5c!��?wy9�������M�%:�<0�Ꮵ��Fwe;P���ee8h���}q\?ߩ-�;�҅k��{T���.(�,�w@8�6i �ZYV��S����=���PS�@�jQ�x�?��!��H<��\������0�0
EGTZ�����z��Ӥb\��p���1�T�Mp��ߺ�H�jh>���-u���W2�W)ꚑ��k����c�y�����&�W?mY!�ԏ�k������a-}5oMo/9W�?]��N%�N4��H�۪k���=(�⭎Ԝ|�d����Z���GNӮ���ڤA4�G(�o�O;̣�6�O�Rw�mE�6��X���|q�ï9VA�i�{Ue��z����Rb���\JNN&{{{8p �?�����������4r�H�ѣ�DFFF�ҥK��9p���>����D}`ɡ�ﱶ���獩����Y��524������gsF��~%��g����GfS���Ṷ^n�̨��+ȗf~���#�ޞ6���w���U�O�q�щ+W��V���4C����ɑJ�6 �����0�(��[WR�������p�R!�O~<���;�j7�0����D=})T�?6�}��`�?⧷�5�e���Dr�8���š�%H�6��)��G��u(��Ż^/D~�a~�����/W��I���X>΍�Ć��^y��±������V��f���	hFDzx�f:����[�è��^KGE��{G�y�0L���>�a���:.����/c�a�N^^�pG._�N��+WT9O\/,--�gϞ4t�P���²�����C�n�Ճ���}�;���<`¬Tf��0?O��&�'tnK!>b���t!hÄ"xc�^Q
��>��K��'�%�=���ǳFD}��y/�Õ��nI�:Ҕ���	�Y���Y����t��U�=�gG��v���3�c._�0�0���N����r��c���	UYڻ<�a�����R�l3�0L����=<��p���޴������L�������b� @@w�b"ɍ�	ׅ}][� ������]�k9�XS��[]u��������0׳��i�,�a�7�Ċҹ>.�fߓ�[@��=.�/�eV�yn���b�9�q���T�}�'zu�@��Og1���ٴp{���^!�T*������$e�s�Z�W�t�'%����9aa�0L���QAA��1�M�.W�^%+++�����'N����4�2(;v�XQ����O8�%&�o�G�p�4��1c(00P��e˖�豉�$�#C��IƷ7F����~&�l���:��X�� �*���m4�SQ�vh�V���molXk����#���Ng�в�'�+�X�;�ӥ��]�<�{|Z0�'�����I�ȏQ�A��U��8:(��EC�2�0c����YY��x棱��~,�T�����+�؜�a����N���MoL$~�ޭ�آ��Qd��MN����VVR��dceip��8����v������n�e����r��OrL.mL���L���.ec:ӊ#��B���e��������U8��3�+�$��<2�/�$Q�r%#�_��V��y�����lR
���"�%���#�]7z|X���  qIDAT�,}7�.�B;�*�۳���̾�n_~M��Q�q
�t5�'e���4',�c��kkkd�Raa������Ǎ��������LP�� 8d��i||<�9s����HKѐ!C(44�<==i���B4�4/�>�����`2�ށ����Q��orû"�7&�����.@�ci��	���b���E�bp��+(P��u�+M�c��w��"~~a��J�>=o�����
��p�ca�<���!�%��X��0�T�ԍ�T\B;���`l�;OĐ�q]��T*�����jW��a���ۢ��kʎ��eh=�.Ptޢ�B`%W�%��Oh�(���UT]P+kN��7���{���`>���G��A�	=�����y�;�#/(/��A��B�׏�؍�x�	�ůw%����j�.T�|��j�7"$Ȱ��s�a� ��a�e322��C� vl����1>�+J�2MG��B�+�uBZ���	QRR��ƊsQ�����N�:���[�l���ϓ��*���ξ��gp��=U��֭[)::�䎾}R����{��-�)Dn'���P&�[[��{҃��������R�x:������?�8;J9l��3���V.�E���i��]<BėSpc���>s���ѽ�L<͌�  �a�aF�舂u�;]��h~滏m ���K.Y��J��&cA�0� �����Q�iB�dgU�����y��c���(�$(g~9p���fg�0Y��Q����9��]P�2�M��k�t*1U���kݒ����HB2��q=�j����}��PY�o�֠ς�uV�P��ϼ���dx�e��->M��)�m�70��B�Dr�(�\�5\�������>*Ɯ�R����4>,�c�1�.iZ�Ǩ�B+;ҕ�Q��JCH
J��9s�����,4��ģZ4q��ܹ3��Ӈڵk'�Ϯ]���p�e^-������+���)3��g����q*C���%�g���%/,�\l1�>��!�[�G3�W*�����_�7,��f��d������ӳ��^�䶵�����mʇ���W\�x�6+����\J��l"'0yY۲3�!!]ޓۍoMe]�B���qߴF���'Ή� �a�Q)^�����>�$#��)��>��3L��]/�,�H�G�0�w��i=9�X�y�� oj��.J�:�X��M��WF~���ٔ4:��F{�_����]~8Vl���JHμ�z'ui�%���oN��RjN�!y�T��������}�|V/W�}.Al�N�J�hB
��x����ܘ�5�����#�����:�7���}�������E6vt$b2i�2�?i�b�2�dꀅ}�0&@�Xrrr�a�@��QV�pJT�pJ�^@u��eqN�����Ν;'J�6��ds��ݻw��={
����TZ�z�"�9yyy�<�����W�}fs��	���U��>���ű)	�@r��ޖ�?<K�0�����(�?�^�8H���k�P�����C�TT"��%>�\�ӽ�������7���4���/-/��LjN���dcc�u�q2�`��Zn��XZ�q�����w��vVZ�W���E%�tC�rr �a�Q7:�Y>��Q���{��T֖�nO~4�����ϮV"�0�	�:��l6�\[c���#�Τ�7j���|އ[��Sq�7�O<��]+�y�7�Z(C�X�؍����a�666�����%���H%'.���w�R|A`Z�hA������)T			B`%g���E�.]�w>�����ʫ\cJ�::�P�C�K���'��}6jm����}��3ɉgG�1��0I���YQ����]ۉ���{���%=4$B��W���MK�b��T��d��z����I�א�:�[��ٞ*��� 69��LRf���όCamq�(i���<-�(���b���%j�}�(�a�a��N�dI�G]|��M��)�=,+�^�g>
().��4��M�ӎ{
�0�0�Ctb���a��1�T��,)U\�0�(����2r��U�h�'ʠ???!FJKK�K�.QJJ�,��0a���+J���i�V��{��ӧi�ҥ��0���y�v��\1���N�O�����cy����ϐ����kI������i�W+(���_���HZ��L
����[<���Xz�͊�
�~�,B���m���[�Х$
pw��G��V��B�ߣb�\S���Q���l�c	)$g+h��f�u���ח5���w+�^�R��a�λ�_����l@/��_I�w��c�aFS���W`W<�����pL��^y�Y�����۪�pAq	=*��a�a�aF����a�����A���:.� �K���N�]��W8�///
		΄P�y���o��*�}�l)R��P.nǏ�}���ڀ���=����2n�@�s�399Y��m��DVVVt��5:v옺��І���$�Õ<�ו^Z������������O�� ~���_6P���T�Q�7~�g��-�k��I�ɣ��6_�adH�8����w g�_�*=\�����<��������|ţ��ay��Iό�MS���;��J��I+��&�aFti�B�ۉr�{��uS��tAT���%��_��o;:�{���4{�}���Jt�ORY�=���}�0�0�(�1�T �"� �(���
�w�x;�/��*H$R[p�^�z�𳷷7�nݚ���E)Ԭ�,!��{p��Gċk����(� �<<<���I|[p�;y�$��8���1l
K�Άbh�e�Xi�}����'Ġ�>��}��(�1ы���˦�茟�ߞc���AI˻~^O�Nn���^������RR��5���t�'���2�r�\j�(�kgmE�[���q�O���zR~q	m?O�|���!�;�i��C�f9�
�o}h�^ۗ�tmO��~�Ҳ����}'jt�d䅻���L=})��C�]�l��ƚ�KJ)���2��lJ:E']��5δE%ʻ7��;�X�NI�!	�Q6�n׊ZH��y���F/%��/]/��'�s��B_��	;+K��ҋ�����#D�H�iN��c+��?�����ɏ��~�1���ZZ:����/-�s�ʘ$ݘo�B�ú����v��YkOW�y6A$v1�}�6^�T"��H
õ�*p��ށ�ukO��B�|)-�6�\��F�q�����?$����W�R�ʥ�%���JK)#��Rs�)�RE^H�mZ�Ck����r�jB�z8�ؐa���a�\�"���QL�0z�:#������B����q�S���������=�����>�g\આ籏�������o111�5�G��PqİF�\n�$�&���Y���#Dj�݇�ܰ�.�a"$+�tu*��s)�T�X�w�E֚Z{���	Q����)�����Ax�R�ؔ�^��ӆ.;����kv	��RJ.k�W��q��y��/��o� ����n��@3��o�u��ό�M��#+��G?��}��X�e�Cowzql?!d���.�>C�Ey���C��~��},��f�4yS#����Qb��e�D'Y,@��F����t� 8��Lˢb��6��ցޛQ>֙%]��� ��K���P;���H����iBh���9�� �~yB�g@8Y[Vn��e�s�vК�g�Q�>����8�|����ăk�o��靍���ݼ�t��Gz�%��g���O>�(�	��XYnI}�\\�t�O|ڹLW2��heg���N�T���ё!�[������米�L�b�ӷuKzo�P���ex�5�V�M��nH2����4�]@�ߏh�M����O$����r�<1�'��*�51E� I滽�i���j�
��������b���ڣrgY5�3�¸Nmh�-#���O�Ҿ�+�fFK��߱�Z�g�T�+߽*<��1j�3��R�|��jF~��p_�����aFb&��x!�Q;�eu8�Q���h�E1+�%p������Ν;Gnm;R�Ļ����gȱM�>�}֋��3��'4v�lt��e�����Im,,b����������0��G����u�H ��w.}�Dڌ|y@:��Mh^�W�c����a4�?)�R21�aX�@�f��t������ z|XOZ����zg���|׻[ֳ��l ���Ή"fc�z�	!��mQ����	��}#���p���	��ʿ��]G�i���Hc;���o4�F!��d�H��2�L�v{�p�ڵ=��fI��5JA�t��x'�\��(N�H���2�EK�'��2ˊu�e��Y�e:�*sԕB�W�#]����~}V��yBŧ �Ypq�bCr�M垻���.����h��Sn8O�����c.���wO����f?+�͙V�?��~�X�%�8�~5o�Vq�pL�׸~4�WGzP���e��0�(
��q*�M��ni07Ѓ�͉+���\-?[�<�'�GP��-?c������P=:�;M��A��� �8r���L�ܖ�����c�	�YE��AGR(*>�dPQ��}�h�A<Q����DJ�l):b<�:���-���eQ+S#��Ll�ի��g$�sS���S�����'Sk��}2�)0q�RBZ�:�ˏ���p*��̙��z�~� _zdhQzJ	h-��{�=��҂�����/�O���kpYa�&y_�8��3J��:� � ��p-SL8�\����X��ws�N�^�}eס��su��Τ��F'�\%����lU�@�v�t^�	���߭NuJ�iCn�G��O_�֞nQ�9n�����RƎ��	WJ�鷦�e)V}}�@zxH�}���#�������!���'Mo/�Y�Y���8z}>g�h�z��|1-K��<\B"�e�~����ϲ�gI6�nLy4e�:�2ҕZ`�,�.]Ż����@��+,����½liT��S 6�M.�)�3з���`OW
��w�	?q9� ��y6���}�b�����%�o�O���Kߙ>�A���	\�~�c|��	��d�:�Mz�X��?�rP�.�H߇�k�R���6^n����4��մ%�"1�0#o�߁��}�E�����#C��q狫v��jB� o��/��O+����o���l��N�݃�$h��5��q�E��C1Ͷ��>�a4D}��l�h�6��rҩչHr�Ϣ�\�����L�)..���t���"K� ���([���z�����g��>��}27R�}�O�����`R[�pW+���aZQ�nf?���-)�����<R��S�	:~Y��Gk:��Җm�����ӗ��{}=����Nm��\Ey)9���~�M���*���HϏ�k(!��UG���kw��]F�`b�� eԿ�u�>�r�΂�v�}��	D�7d_�E�?����ڼ@L � ���Zn>�o�1���E-�sy�t}�6@ؐ�����4��v?��v��W'��kʂ�� qGx�����w�Vn��}�7����J�1,��;m�(���K��V8�up|>�5� �h��;i��X!�M_��r��-�D�<y_���7�Oz��������ā�����Sy�̔��n�kyeh�g~����{м�a�Ѭ�4�GG:\�θh�qZ�|K��Dֿ�?E>0C��kE�=]����(����^�����D�zpo����R�	b����2�z�X�_��?Cڷ�?�9����H�`�aF�����D��Q���D�/$��i�4Ni!�I��l�#���g��3�������C�#�퍑����}���N�o0����op!ĆD��lc릆�}�h+++!��ӆ�Ø��э�v-���/�u�U���$*Χ�Rm�L!���Ա�bH���8����RJ+(�܊	s5�X���Қ
mtT�e8��SS��>m�S�";�t��>�A�,�h�EZk��l�`���m�j|����)P�u{HNh�O�"BDY����~��Xd�B308W#(%!�J��rB�8�1A�D��rՙ<�qٰ�G������+,2E���F���zw2,�c!�M����BL�&���4[Ƌ�:�k�N:v9�e3�w��~�'�onH��LJ�p{�`�p��_g!���Wd�7(�b�x�)��]ڊ�w���q��NW2����p?z�0�� ��ڇfҴ�V(R�?�G�X` X�xk�>�k�/H׬���42$H\߰�2��?o'á�ѥ��sK/!&B�H�ȡ�S��[Q�[��O�� L�{ߗ;���?��2mfH��V��<�T"G��|�^��s����y}�����v6tG��bñ�=*�~�<I�|~ʚQ���	3��Y�z�i��;�y҃�#(�ߛ��r�q�6�	X_��Z���E�6-e'컥{�!B=�u��~=pJ��!�G_{�m�x�]1N��ǯN(\|p�g� �ߒ����y�Kk�L��a�K�h!^�S����Ʋ{���b�5�E{��1�)^\�S$+<3����+��.�����&�/�b�58h�O��j���8�AꗍY�L$6%,�cFs�+/D}%%%,�c#������Hk�����{	78s%_Q�;33���N��.���h�}F�J�sB���7��hc<�O���b�?�v����}x}�c��}��?���wue������fPJv��>X�w�?���o��ū��	�	)�տ|�e� hDɅ}q��G)�ڔFP(ɌE�u3�݂����$_e�j�.��%������kv�^�gd� D\���Қ�4�{���Ey���-ѳ�%J����ֆ�o�$�ӳ�\�(��ռ��a�n8!A�'��Ձ�� b���>t�����=9���y��B�j
�� �Xx�H!�-}�
�	���Qp.{t�Z/�,�k2��,���W�GJe�Q��W���m�����c�_�����牑'8�����?w��nı��K��ώ�CO��M;�Ƌ��k��y�k��iN�'h�����;�|�,�� H�� �1�±��W�v܋�@h��?&�d?�Q����-��p��=�}!�[)�'��� ��~�CC"H+<=���j��#������-�XFK}���[���f1��f�#޷�6����0�˕t$��15�����:�~���Q�����^�a�XI/OJ׭祾DS��m8cC���.�� G�����{?SV~!5,�cFS��rs�5(�2���o�l�u��Ud�a���N�f6�>�}bB	l��H��~C��A���m�#\ກ.K�biўc�/'�I"���@sNώ4Oڰ���E,�`{o�0Z�Xp�v���<����ݿ�X���w����P�;�Z�u���$��wE���~b�+�ֳ�B~����k�ff~!�LL��93�D� 69��T#��.(�۾_#J���&��?�N3�^)�)�V��s(��x�`
�~�s	�~��"L����#�l�$k+K�w@W��G;��+�ۿ��^�t��
KJ���5���C�B����%e�{���B}=�X��>���C2n�!�
��p.aga��f_~�̉�������sWkN�D2�1.v�#��a\\�����8!f���n��`܈$�^Ac��p?��!�0���M~5o��$��l�pQ�/\�Q�C�:j#�3cv�/���0�A��]����Rl�Қ6	5�~W@��*\�1G�;*�4,�cF3@�gmm-�����YM��9�QI�V�0�0j������u?6����7� %�փڝ"/$���D�޼"����Kp3{m��D�p��w����tZz(�~�b��pQ�1n�70��Ss �,<�"\�Ԅ���#��}�!�����Y@!?���:�F�LkK�J��4e��T�b����D�E%tW�."�~ŽSi�7����h[.��lPOB���3�On5vDr���pb�gWn�?����g��e�[��L�,ݬ(Qf}q�8.1R̜�ӘcF%�=���"�+%���kM�ڎn�F��p�\E���I����8C�c5���t�_�Й_�ϒcõ�ڔ�[����
��㱇����Q��a�ajˌn*�� O(\�j#�W�����&�\ '���YK��l�}l9(�BՐ���.�M��3������g�c~��`�9h���aM`aa!D}�(�E�a�a��?p�0�lTq�����Չi��XZ|0��\�&Qc[/7Q6�Q��ⅳH�B!��b�;ta}폣��u{��QMh-^F�ħg	��aZ�Ih\�Ή������TM�� k��[�DsC�+]�k[GN�U� 0�����Z�U܏Pb�����v5m��ir���ZZ���_���T�t5;O|'З�Z�w� ����Uܗ�]8����,�a�	zq�N�ȨVJ*�xm�=��u�;{�ڝ�<�u
IAؐ04+��p+�;w��>b;�xM�c5p-'O�z�������a���k�����'3_~���A�8�����>`����~��$?Qr�Q����[�cfC�+�sG�\Iʺ����~f�Q��������[F�\Ij�q悾���5���߷Т=;��zu��n�W��16F�c��16�����62$��R�Vs�;�ck��O�M��ͮ#���nbNgv�P���CR�7���Ϸ6���("��"/\i�[��t�a�F�w!�C�ݢ��3Z�a�a�1����@z��.~p?K��#�R��Q_6�Sӊ#��$j]K54��'wmG�׏�x]_|����p�2�-Z�%����}�}^���%JfS�Q�3�ӕޘ4��[��ޥ���",�����\�[�Ҳip�	0�����wPAI	-�S��.��$���j�;t���G��1��[ou5G�}��p/�=*�>�e��{�����b� ��zv���ڀ=��Ƶ�\�ҳ�33�+_L���� �4?'�\��^A��l�L�-�C��;��gm�K�G��C���Z�\�+mSs��U��5<$���RM.�w��^�/�D<���G�y�2O-����_9^�qLc�-�{,A�cC�j�����J�P�#^�u�*�$�����!�>�5\�q0_9wџ�ԜO����mZ���a�1�K��������i�P�a�a����N�dk--��
�� 2��,�4Ʈvp�B�{u4L�A����ؾt��kUQ�S/j|c�,��1X�]�ʆ���=����'��������hԥdzy�.E�:���P6#.5�u�Lr�D�3����Qx�7��y?m��X��v�M�Җ�ot���F���z��}���8�x���<����p����յ����D��	q�]�i����j*�T���su2����^bk��m@Ojv�e{��#?��Aύ�+%��*���\�7��(7Yb~ώb���u��cn��Q�K%'�0�A{��}π��4?�M��A�~�s"������Bť�b,xπpန(]�1�D��I�K�+�r�c��Ù��>.{���ʅ�'Ή� ;+K��	4��Dl�����[�d�γ�7��X����q$>��(��~���.-�{4Ak�jkqD�I�!ss1v$F�%�	������Ԯ����FT���4�:c�.%�}A�s,nX��0�*�C��
E�ݲ2^g�aF~8��Н};�?�uB���/�eQ1���t������G�/v[�^tk�0�S:�p}��M��S�N�fP:����N_WG�3:��o��g8P�g�>Zr��q���xmq9#��Z��>�e�X��׺%-�{�(y!��J����lQ��z��.���']����-�}zpM�����r��3v��+p�*�`b㮳	�=&��8�Ҭu�-�Z�[X$��'��Dm����pބ8b.8{Ն�F��K2R��ĸ�T}2k�pȂ�����]�Y��5u�������,8�U��1M2#�aԁ�k6;�5?���Bq�^C����b��c����i�����o�t�B���g��K�!+
hA3����n;sI�LˍeQ����^Ծ�����6ێ�񔒕+�M�fM��V���z�Q���{���8���-!#��~W��7�9�{�ZA?}h84u��T}?}'S}]�|\�Ԝd��q�>��$��~�<��b�@f��0�K�p�ק������u��I�c.�������(��f��>�aT�N�#KKK!�����һ�0��,<~3l%�zs`���t�O�E	45OkL��	.v�R�j"�A�hh�@��T0��֔�b�p��ㇵ��v)��/�~ �).)�Of��l .��B��Vb����/�Ҳ��A�0,��Z��۝�� �:��]�������aB����nu����-,�w�5��+�%��0)������Ld\ӔSjL���.\J����'�21g�p��rTW����#�}��Nm��91H3�����潿l���M.� �=[���"8E�� e��(��`^���LfQ1=��v�#Xd�����g��Elp���A�0,̛bj�v�b�C��H���,@��j�� ��J�.y�o/�/�"M���%�3�xa�
p�n��q�r���ji���gh��bLW_*_�����=FyS�i��$-��3�zӼ�;���#"����8K��!�	��nIc�Z7y�������f��>�aT�ޥ����rrrإ�a�Zq�j&�^�Kd���@)+���0Mɉ�L��tg-�g	1�Y���9�਀n��K�t�B"]L��1��GF?����	rd�b��I�o`-��`cMS��ei�	�$�d��#gh�Y��W�/�X�"^ĭ_�h�(����#�$�8a�hcMJ����*+^F�Y�sQ���qO�pJ�f�1���I�(>�E{ϗ�����'��p�ؔFrV� ������q���Ծ�}�J�J���"A��,Jp��^��缥{�CatR�b˶b�����B�ҕ�:�x#q���p*N��ֆ��%��9�W�؇���+�W.�a�ȁ��4�ӥ����"�I?�u���g��U;�c0������14�K[�����Ab���m�>���6N܃�c���x|�!V4�ЧI����� �5���
��Zq���q?���}_%�3���uC�ZK�b�&gО�U�熎#p~/���E��qS�3ƕ��bd��<���]-�=쪭R�fo[��ɯ��MK�"~~i|1�jJ�@�ݦ쫰��a�A\� 䃠������LH\��%��#h���\Xc̃r<��>N��0�0��M��uZA�圞����~B�7�G�,�Erk�������={���o��Dj�[�7��og�ѡ���� e�0ٛS��id���"&Q���Yr(���bn��PSP(�-V6�B\��Lc�{�����g����m��;x1�~���[�t@�����?wR�����{�	�
\��-��;&��

).5�b���޸˲p�
��ش��vY�Z��8����7@	:���/W4�g�%jił\[�JUN�j�(�G��+���<�r�� I�ޱÊ�X��m���y\mF�@P;E�Nc����U��`�SUІ�o�~��P�������V;+��r.n���&viK��Z��n�v"�����(J�a<�y\{��ҵz���]Z�g��V�<�����mk�LӒ��o�w��(�;�㕞��KD+�z��/��s	Կ���cz��hj*�ňzG˦��}�(}�]l���TP�tO�a�a�����~B4��{~��V"�ȼ��yZ��Q䙑������рZN�����<P��J�:q[bf��p�q�	:{5�� �4Q���Q��diq���9(1��7E_P��2Ė��qi�ūBd�o8%��O@`��qYSF��mD�8�P�?[)s��%�^^����w�bςb�c8|!q��'gR���h�Ԝ<���Iؔ�rV=#6�a�aԇq�#�7P��J5�p��<Q��!�>���ݴ��Yb��p�m����4e ��QzA��
��.�0�0��Ҧwk/��Q�c�n�nmb�Ȋ��N��,��щ-[A.vzqBCڵ�Tj.[b.
q۟�ΒZ�S�s#�k�����ȓ�Z�b�a�iL�V��a�a�a�i1Iׄk�{�+z� �f�B�O���a�)�Å��ׅ�h�_���i�yOE�릀�}�(}�]�1�0�T� �?��g��7�<��J�:O;��!A���v(FlZ�6⶟��e��@un�(A ��{�����P��ۛ�7����PBf^��¡��ee���]�[Hq��ϑ'��e�^˵�=��=�C|��hj�t�sY3�V7]�~�j�p?2�۳���>��Nm�|����h��(�=�k;��-�C�ͩ���{ht�`Q5���'�s���w��JM~q	E6Rŀ���>�ad���.��%wY��0�0�	�p�;�0��˶ӗ��/�C��l�}�^�97!n�Y��p�<��b�DOIim��@?E���N�5�m3Ls����4ʨ7�:85�=�ٯ�X� +���Q"���J)Zc��=��w�
ڳ9L���ʎ��˚����q���*�W�����n���_��땢Qc���p�����k#��1����R��B^N��𐈛����8�#C{~�q�	�+*����}���3��S^^)��0�0�)<*l�ZL���v�4/�,=}�"J�bB�)�M	�Ջ�Τ�Ӳ�r㥴,�2(�зuK������;#E6�P[�8�qs�c��Am��{|�6�}W�5������U_��|.k>��ƒ�Ϥf8^�WMp��W1BxŔ�/�{3@�Ýn �����и���Zn>55o����vmO֖Bط1��M�w������S'{�sna}�� 5%,�cF�E|�ǒ���1��1�0��+�3���PCp����y�V C�&�P(W.g���_�����I�H}s��@Y��MXn����颔vrV.��WJ�̩�������Aݪ����bzg�~RZ����+��o-��e�/^�$�a~�tk�0��=�0�kLBz�h7��i�$����+DLPWq�~�4�&]#5S�㫦�A���}��V��c||�t.��9Ә���ʛ<� ���Z�<e������Jk�i����ʨ�~dL��*����׫ʨ���)FS�Vi��vS?��_7ж���@��m~���y��b��Fcp�j����g�.�dkC������k���H��4\�P��?�o�u �1��@�g,��cii)���a�Q=zqL� �}���5��O�@4������ÿm"9���9�i���Bz�ͤ%��n)Dn���o�Ֆǆ��/w��³�����L�K�C��7Q>(_�y0q;-�=��ّ����zF^�;y^����qbRW	�5�����㭌�UK�H�	�p�p�H63�q���7&���GU���U����H�l{���w]�m���b\��\	���Uoe8^�ū��JJ�)'����e]�Ȧ��V�/wN"g�0��Yb>��/&QjNe�H�yj��D��-Du@���#i�Ԗ��ujK��-�\�KaȀҾ����f<��˶�Ģ���}�b��t&��Q���|��=��Pb�>�#�0�0���q6A,6��r�!A�9����|� �<OJ��ʒ
j(�9�c0=7��A��0r`Z���qk����?���ǖV>���|r��F�'�nrfj����E%�SP$�@\��?��o�b�C��)ĨL������z��R�hǦx���}5����B���:�1Jȼ����������P������bD�֦��� ���^Eƫ�s��^]�[\_��&�{�<8C,�U�G���z�CK�TZ�^iK�ݗ�ڿ2��G�h�zeea!�@�_U��^)-�֝<G�'�h��c7�߀xo臋�9�hH�V�9���VH�����5��@B2�3�Ֆ�>b�	�]�\���}��LF,�c�_�����R}��Ղ�i�ƛ��A��n|�0�hd�틻,2�>�1��,\&��-ȟx{�Q~
ْ9CrDw�Jsz���3�E��O���[�ӥ�,�{�����}`bIO��Āyk�|��V�'��S:>v��)�UT}% ��;XZn>�O�����*,��L�!�(T:��vDV��Q2��D9�����!�t%��E�������`��F�j+^/��m_�Z\��ѷ��n[�������.��k���)�I:_�f��P2�U�H�*_�^?��!&�gFt?�NNS�GMq�Iq�H�"B�ϧSҨ@���}��f���Ԯ=��+>�:�d�_5���!����GM�i��7���e*7E_���b� �Ӆƅ��V���u��C����o�Bfc���m5�����W����.�2sT|?2Fk�9�r��@_�H��I����c���	tw!-���Y�v�i��1�?��"i羁�B���`g򽨈q@�~�~8�~��m�
	�ٯ��n�R�G�������IGR��#�6Jc�����>F1���
g7������2�0�0��嵻i݃3E驵����%��{�9e����aM��[[��{�������:I���4�K[���r:��J�zu��NB�o��Y��\R
(]���Q�޸+���--�	��7�Ǌ؍�K��z�sl�E{���1.���Hs����D/��/JT�rF6��ϝB�)w����t�rG2w��B���-H� �6�o���5mef�Al�k�};�r" :/O@ύ�+�Q���cg��Q��߹�X|Ջ8�����焐sۙK�'��a�C��9� ?Â�����P�x�*�=�����V���B�@/؃�����^��_����O��U�������sl��G�{4���7��4N:��o����۪F+�����Q�x{j��q�JI�����j�^�h욬�3]����otߩ5���eе�|R3H�su��"�j�!�kj�����>���$�e-,t"�s�X�m������ǿ���z�����Mi�:�a�a�a�	�{�2��=���~B0����\�9!k->-K8`9�ڐ��uiقF�ьn�7d���zɕ��5�� z��FrV��d�ws�w��Wg�Lx��{OA_|�;�ӽ�-�{�p�3�o�-��$��/b��XԗWT,���ʒޟ>\L4�qT�.� �����C������Z!|��Q��~DS9z;;�gۣHδ�r��(�Z_���NdmiQ뉬�Fo|c��,�x��)�}�u�.~���u"]d�c��$~?�;aR���ˇ�t��ҵخJ�!܃6�\�N�Y�J!�ߛ*�չ��!}\K�v���YE�UWjs|��=�/\���ڳ9����5v.�9���t���S��7�?�x#�8r����b�^���6q��{h�o��*�v��Z;��ڿ2���C#hR�&�� f� 0�	�]�"Z��;�3����zEJ��Ʈ��@�dlL�SZV&ܱ1���a�a�a��w6��PϏ�+J���[m���=��%l��&����Y쟽�N��Y%� [t�-���� "�����6+rЏL�����p9�v�1��O�`!
���ߕ��U�������t&%�m������AB��ߩC���DP��Hό,�a���ZjN�(���&pmD�yB�x*N�Γ@_>��ҫK�%�=��b���
�ڻ���lK���i�x��oJ�rKע\6�7��c��zQ���a=Ć�}��8-��i�(��y�U������Җ��KJdV�����������Z�W�|���e��RpW�M�P�������Ϙ/v���>(�Pz��Zا����ڹ����X�:�E��U�����Zc������ݝ��VX��0�0�0����(w '�Q��7�E�
\�>�E?�?qC	*9�����,x��*�� �׻�н����]N��_���y
kbP� Q�<�t��(���c�c�<zzd/!x�j�w
Q'�����	�����"�!AB��T��bE[�8q��V�����"��R����	dci)�Ϯ�Fr���̪��u���1��9�^��gEk-޺`\��ݹ=;�-��452�?�9�^�4�^_�W�g�{� JŨ��%�{w�UW\uEk߃Z۳9�p|�#��p�v��5�����x<�\��C��db�p��rr �����m5���#U��{߯i��x�ܞ�_���6�0j��}�0�0�0����I4��(��E��B�/G{�ǫk�yt*�틻,ܠ�,�ӣ�@���B����{I��7D*V�p����Q����A����������1���A��S����ד��)V�'�>��%���g,�3f�����P�p+�ß�I���~��B�X�s�ϵ��\��ޯ���(�b�=�@��9.\ˤ�6�[�R��P���7nδ�ީ�5��\��s��T:(w����UW��=��=�ÿ"^C�Cƫ�ҳ)��U8x[[Z��X��[�'���!���[�K��~���mU��s�-ޏ��;E3�ן�WT��+ՠ����6�0j��}�0�0�0���k�b3v{S*�N]�2;�RZ�a�p-]8�
&���KITjBu��U���Nh�<!�k��NJ�}w��XQ�!�D��]#�}�Z�	�>�N.�qbLOG{���E�+�g]�׺\�x:9M�]}�v�ٯE�m�:�oc���J.����!7'ש�ZY�啱�9u��XZr�E]R�}�w���B�xq����XZ����Ju�W���~�t��=����Yz��s��_$X�?�T��1[b/Ҁ��"1dz�7$Ȝ�r�z�R�V>�J6����N�^b�rF6��]�����e���́����W�׫��b��ő�W*mϵ�?+�z��F����a�a�a�i4�®�ZEF���哒��w>S�d�Ǥ̜jK��D0W�L	�K0�	�ju�M)/�l�ӑ����ﯹ��+��=}辁���o���p�A�V �J9�x�ⓨg�/�;�k��=}���s{��8�x�Uzn~[b.#?�x��	ɴ��tg����-^C9���s[lr-?+��j����u��� JƵ�>�UW�;�j�j۞c��ъ#�U���y���e�	��G�^�8P8}���nx��ȓ���;�t�������ː`$���֮WZCk�Z�W�������:o����x!`���z���WQ�&3��`a�0�0�0�ԓ�
�J(�B��W\Z��H^Q�x�N�'w�U�q�����Y��ݬ�惡�~�q!��3��?W�R�/�������\e}�����l�Mvg6�$��;$��"rA!X�U��r�V%VI��4�V@I��hZ�
R
�`�"+
��@�E�	���n��˜��I6n ���3g��y�I����>�y�s~��wbm�/���Sw�{��ba_)�^�����q���o;����_v���^ˮ�wד�/os��vx�mć-`�"�fOr�{�[�#gI]����S&�M.��c��g^��:���\�s��}�a;���5/�/�ي�q���ah^[Xp�����YS'mן�*h�l����
l_2Z/��ɒ�~#ͧ-Sj��O>�����{�'����_-�����E=I�����x\�{��ێ]e��.>w��?�U��t����͕}yPR�W;34���x1�;g��`L���} h��־�0�b~U�\�vׇg&lL\@a     {����������-Գ'.�n����;f��U�UZ_\��^�cJ��mE�;��ޒ�Dun������������8�t����_>��K/U]��zO��Ж���ӯ���ے��œ��{s���{�cG.w�O��+vآ��cSe�>��_~M_��|���Cqp���ݷ�����<s��m��\z�/>h0ח����:'�uҐ\���:d���5R���do�?�����'�vٟ����#oߺ���>D��>|�ݿ�w�;Uf�r�����ϐ�v�߮�_��UY��_?<�����KO{�4�>����+�������uڶ�e?(�&�����̵�M��jgl�����/����ھ6��*��h�Ǚ_1�:���և����    "b�,��#%���{����K�#��������^��?���/��g�Kq�՚u��������U��'����{�����3��?t�R�����Ŵ��O���=�k��uK��������yg?�lW���{�(�ٓ�ϯ�?=&�If�X9|��r�����wV\EƲ+��_~�T�ߗs��]��y�v��~ڻ�B���>ٚb!�yǾM~åvm!�~�F��OT̊@�=[dl/io������B������f%�~���Χ���y��b��^�)��Fʵ߃�{�c���]�+�}��wl�{�����}mQ�?lm����VXݜ�1���.����#yh���:I����v����T�	��´��#����?T�y�q;�6;�z�Z^{i��N���P��_1�a������a i(�    `=��r��i���{t21�y��C�|���g^�$��)�좰��,�WʊnϬ딿����O}H������R�ӓ�od/k��%{��R����եv퉶�}�x�;~��v��F�؂�{#K�{TN8xzqE���W��0j�zl����K��GW�7�j��7r��3�k��ھ;�Ƽ��6����ü/vy[%K���s[ v�n�מ�\|%����}ٞd���wʇ����i�?,3���@��>/��ò~c�$�k�k�:�������$�����Չ�l�]�_�8^�j�\�y]{� $�}    ����KZ�eWΊ��7t�4c�/Mk����sR=�J�e&�Qaߙy�L�_<�o//g���W���n��{E]{�T�G�����+��Ѯ�vR�M2�#��ǿC2�����׬� K������*r���}�� ｏ�?Yqy����C�ϑ�7d����g/���KK#���v{�+n�K3�C/=5#�;vՕ�}�yy腵R	�j�������H��}�{�.o0�}��ˌw�>۾�^ִik�U��睱��� ��i߆��U���
lߤ�˶p�ގ�oo9��/�kWﳫ�>w���ƾY�>�~��Xt�� ۦ���0�H�6^��8������θ�z4�����Ӱ7W�W?_�����	�\{� T2
�     "����|��dw=�|�撏�ǣ�����*��Y���*�S��aW;����Jb?���'�'߸��r��{˱�#S3d��q��n:{z���s��^.�F�W��Jv�wJ��4!Yy��Rۊ�6��O>�%g��/l���YS'�Ǐ:��R�-T�dCs͜2Q>dJB��Jj��L>�kW �7�"�<�v�$E���G�y��a�\�\����k�مף���_�k�����o���k}�4�    PF/�p��0m��߾��T����m�jvA���[WҰ����wk�y��Y����ʥ���������-�+�Ԯ~54�=�S�ݻ���7鿇�炟܊��~���~)�~`�����˾���+׸�/'u~�3.������0����*1\��@%��      �z������oF��P�۟x�xK���)�~�嵫����oI�Ǿ��:��x=J4^���?'y�����
�              �
�              �
�P1������GTU D����g��R������:           ��Q؇�a��@ycb�-           ����             ���             ���             ��� �0�l�u�])jV{Ƽb�Ԧ��;F7V�����x����N��'*������m"��           \��Y)FV��*c�+�'�Ft�=���R奴ƞsV1��?0��Y��33�g��AŢ� �&Pџ�{���6�5���j�[�R��`��MN	&iY          $��b�
c�F�ޮ����xK�k��ޥ��V����(����>  ��1&L��G<������QS�mw�7>��۷dn�غ1�`������y�          � �WD�c��뮾M���_��.\8�%�+�r�b�%�dMߦ��D��9Uk� 0B[W�*c
׽��ܳ�o���K�{7��<�}�EK���&Q3GEk          P��:#ڪ��\{Æ�����sr����-Ӹ����*�IQ#�%
�  &c��*޿����~J"_��a�Us_	���4-�2��c�AU&           ��yUE��������l*Ǐ�om^�]0���(�|�9+�
�  �-�/F��9}�evKt��=��l�EK�
W�].          OF|Q�w���b�z^�K�C�7�_
�2����^����S�Aa  �`��o<�l�U�Hm]�����%�������          @��&�}6���1���+���in���,ѽeGa  ;d��F��i��-g$�ϻ���K��~���?( 'g:�ؚh.^~[�^����W'?%�!GO�&�Sd���RN���=���ap-�� �*�F��*<q��ٌW�Y�x9��F�~���WQ��x�[�oD��*<��"w
�����*r��B��	sm�O����^���↛&�k�7�67���eEa_�3�HGG�$I6��t��]s���ſ�<�x�������ߍ;v��+
RUU%�f�k���s-�VH�r����?#��~������ Fa��N����Qmc���D�ڨ�Sʫ#¼�1��I�и�w<y#�x����X3QV�z��b�Ǝ`���Qm���*4��"�Z���QXƓ7r���������OW�b��x���\�2�
K-��u2^�f�y�'L�gs����cr����5,�
�qIßd��ӳݓ)�IDU-#~�[�*�}	�aC��]:555;-�EE��b_$H�tuu��L&S���b��
&W�I�ֵx�j�Hj�-re����}#�̰� ���z�&F���=Y��7�'+7��d�F�p���*)����+JfۗQm�bڷD?yC|�r#o�OVn�����0߈-�{�#�7�'+7��d�F�p���*(/U`b�\��gN�-j��T��r"��6�=�y溠U)ԉJ����Æ�ߣ� ����ߧMᴎֆ���mXT������}5?Rլ           Bg�S�@~Q��p]�7d�/y�����5������>  �X���Tո�:�>''	�����L����_�*�          �Y]��n\��'I�ܢy?�kn��/zW����,
�P1
�5R3Ft�8�B_o�祂W���M.���.�k��JY�쀗>=����A����d�?,j�`�          @�c^т9u����ڰ���Mmg��rQ��JnE}�hT���ϐ��Ӆ���Qn}�@Ƽ*���M-�*	�k��7Ӵ��U���	          �d�Ȇ�I���>�I����g��><�7�x�TvR�gQ؇
�BQ��
^ ����ښ���˷���ls�;��_          @��~��u��p����6��CT�	FoE}�}  g�/�[�G�j:���t���           �Q3"�s��$��uW����#��	��n��,
�  ��;_�q��d�TӢO��~LT'          `�C����\;�_Z�1����f#7��>�¾
� 2}�tI���*�0��#��Ζ�/f��/~G �D�	�}��+�K�ͥB�xq/���J�=C��
yGǵ��1��X!��7^�;:���c�ϱB��!o��wt�/�7��H_A���B7��ښ��4�_<��`d�Y�gQؗ �ƍ �󯹖���Q��y��4-�d0�~� @	��/�6m������S�.)�B�d%o�H6�탥��?�3Ǎ-��k�)%m_���8��;e�Ԓ���Ul�1^�&����;z�76_m�?ǀ�x5j���5�W���y�#�����Flx̟G�P`�QQTZ��?%���v\��x~��8F0<#(�(� 8Ƭ��v.��Q��^|��`��\ ��كRUUc���v�a�}�I:����ޒn7��������{�}�+`���4�yKݾ�?�mVW��Uq��A�0�7��o�9��m_{��j���W.�k�����ui�u�}���1}=��R������t��4�����'���b�*3�^�\�;ձ��a�q�T�?�J:�|������&.[��7K����+Q)ݥf�j�E}'�+H0P~���	sS�{㬣o)�vٷ �V�f�+���G?*PnQ�o���7� (�8���e���E��ГVa������fa�Sq�Ѓfa���;X�����}-ƫ�z���Z��-/�oi���_�+����R��3T��\6�W�4�Uٸ8^�����e���K3߈=5�u�.�����>�mj�5���-ع=(���*Ț5k�
Pwf��F�{�w N[�q����y*�}�OO (��|R4�"�Aq(���� 7۷��y�8h��7����Qe��^��k���U���l�i��E;�����I��w��v�}]�f�*�^�\���둵���7N��F��Ǝ����7��x��ϲ=F�f{X�g�� �a�kr��To����t���6�� @	��`C�'q��X�<y]k��<��(���N9�2^E�y]��e|O����2>�.M��RKӟ#C��ӼE��_����]1��*q��u�����;��g�7��>�� ��.�=�����*Ba��+���rQ��X��y]k_��ż���3�U�(�Ny���w*�9�o���92���Ѿ�9|�N���#��o���Fd��7bňl�PS}]^0����x�mg�E}�}  '���9���t���_��mu0՚) PbQl�CE��2���Z��7,��-�'��£�E.���J��e|��9<�/�Fy��v�����aQ��K3߈�y��9�_#�6���y������((IQ�Ea �	��/�!c��`~��Dq�AcTDa�W-�7��׵�%o���|�JO)�+�t����[>�����o鑷|��7-M.9�O����a�)�[6�-=e��[�1�v@�jۍ��K�u%*�(� $�1O�jzT�c��L.�" {��P�(}}��lƌ}cu���,���������O���a�/y�˵�7�xUR�gD)�xUR�y�-+���eE.���u�oiMg�-+�򦃼�о��xU^i�ee�y����"�7�=s��ۅ}%,�(� $��_�N��?��x����C֭[ʶ큆�y��׋��Ǽa��i�%n�[:���xUv��g����~��P���l���a����;�����kO<��U�L��x�h�6^����4����k���W�3���P�;��t�꺪qU������A��Y� ψY!�5�+��(�}          �#*�
vɞ�WQ�
�B(�(� $����~��`�L0	U��	          `{F����'�5�5���T�gQ� H4#�����y�.Uyރ�/          �72+�[�s��II߃�T�3B,�(� $�������澒ij˩jV           �է�����R�iI���J҅\�gQ� H6�U�a	&W�wG	          `5f�`Ԩ���ջ$�"(�(� $�Ê}�et�(�}          0�����"HMna_DE}�} �D�|]+&�b���          �m�x/
�ň��س��Y� ͤ]�a	&X]��`         �2�s�y�����L�E}�} �D��c�5LFma�          ����[0,�<�\��>��> @��}&X��?e�ďN          ��3�e�+q��T�gQ� H��*�$�ф}r          �=QƢ>��> @���F0,�J�          �P}�~�`X|�j�$\���E}�} �D�R���S+\�          ��y)
��IE2R�bP�gQ� H4`�5l��	          ��z\)n�Le���IQ�Ea  �|��aQ��X�          ����+5�_Şw�QQ�Ea  �Te�`x����          �2����eDfV�Y��Y� ��&X�T�,          �
��Ǩh{�-(â>��> @�ӆ��5�q��hF           �QU�;��K����F*IL��,
�  ��Fߖ�ⲉ�+?�)ة/��
��          D�V3�}����;U(�	u�9�E}�} �dS��}���;L�N          �����I��[;��승
ő�,
�  Г�¾ݙ-          ��P{N�¾]2��*�*��Ϣ� � ==�R/ءL��C��C B��r���~����Ǎ'qs�!�H�Pe�q�k����
�}���%N\����Z�q�We����۾|�p��l?��y���e�q����L�Ҋc^ƫ�GF������t�y�[V.���xU2�h_aTN+~5�7��o=<�J�UHQ�Ea  �T�mn=�kq�o�^�\��؃'N����P�'��������ky-��fy�C�CA��sl�r�������a��1�*�|��\�G>�|�\�Uy�y˃��<�[�����Q��.Zz�����Rz��]�Y� ��IqAaߛ�~n�N@ �Ԣ:�be2��lp-�e�}��о�#ox�[.�W�Q��А7z�y�G��d�oDN�ϡ!o���F����0��%�`�yg
��Ĩ�%��Y�
+�(� ����dn{�,��l3���=���`��� àrl o��򆏼�q-�k��:�F���#ot�>��Q�s��򆏼�!o��o�9{��4�]8g�`�l㒓��$�*��Ϣ� ����1�ɜȵ�m
�M�����T����q����!o���ϵ��Q�sd�>�F���#ot�o�O�ϑ!o��򆏼�a��cA�d7vm�t�p���<�/qU�E}�}  �\"\'2��4��U�|X ���y�aP��=򆇼�#ox\���?G���!o���F��Fx��9򆇼�#ox�=�;c.��������z�sz�k%v*��Ϣ� ���j�?�%r�@RF�̭<���A�AQl o�����[>�-=��F��eC��#o�����[>�7JO��eC��#o�����[>�7�,h�ٮI��D��1�eǪ�
/�(� 8��t���?|���G�mnW0�9+��+ �)N�y����G��!o���t\���?�yK���7�������Vڷ�ȋ=��We��[:�-?���!o�1�x3��>�͛�-��[�in;Z�����	(�(� ��.M}1�_ �Z���n���mAJ �<ϋ�A�A�`C.�+�6�a��&M�$�lV�&��qn_{�����d���c��)�ƫ�����r*�k��a�Wq���W��g)�Ul0^a�*�}]�r���}cc�}��y�#�񪒩Ⱦ}�.~Q\u��)�W���U�R�gQ� p��%����uU�*qP�{��/�8�I�R�S���������׵��y큩��ω�b�J4���5)_�ț\�M6�&[��F���i�?'y�͵���Wɖb�Qa��n~ۍ5�NT��+�wJ�$��Ϣ� � ��Vκy��rvAR������\�/�2�H���p�T^�7�
��D+оH��o��7�țl�ER�/$y�����D#/bK%m|�V.��D�vN鯻c������:휰�>��> ��T����.ȉ|Y\q�5UFzn�O          �����|E^d��bn�X-�M�R+q���>��> ���\�ij{ ��p�8 �P~=�Y/          ��P5M٦�s-����cLk��H����Y� ܥ��5MKN�n��R����|��A�/          ���Q�^����\K�c�`��%sD�?J\$��Ϣ� ືx��=��t~�Ꮢ@��K>d���P�          %��sW�Em't]���$P]S�������	/�(� 8OUg̏3��Oʷ6wH���o}����AH^�          ,�S���1a^ۉ�4�I$ۼd�1�!S�Y�� @���x�x�'6-:��e��� ['W�Uu�           ¥rh*-�����Ԥ��gW���ܤ��$)�(� ��/H����KO�l���T�LS�9b�u��j�           "���/d��Oϵ�?&,۴�SF̿i\j�*���K  &�I�4_
��6�������4gݜ���K����6�           �6ը�/����\K�-Ri.��*S�s��i��p��Ϣ� �7R���q0�Z�뮞/���
0�yٔ�y�� ��� 0Z'L���u樶qr�C���Kn��KV�L�r:%�!GO�&�Sd���^m}vо�Ԑ7��]�]E�H1^�'y+�ƚ��7f3^�f9�U�\����[;�_Em6�Uhne�1"��o0^�g9�U�Na~�[�_En6�Uh�7	T4|�9��v}�)�y���G*�ĦE���sS��x��KE}�}  ��,����|�����ζ�'%Ʋ�m+����Ǟ* #��'o��'7�xsŊ�mW�ɛT�M6�+$�
ƫDsm�r-�k�V0^%�k��k��m�U����*�V0^�R������3K?�o���ĖѺ���}і�t��� �]Qy��~�mj[�N�^���K�$F2��V#K��          @������6��� M�-�_��mZ:ӓ�o��b��>  vG����/��h���|�~G�����G�вO:��Wc��lc          _*^�弔I��mn�Ƙ��5�]�]�)[�z���KD�~�*A�P� �0����[�*s�6�-J{���
~['V��~�q          ��S������S���݌I-�r��(�����zF.5��Xe�?� 0B�:-�k(��<��~{0Ź~CMǝ�p�@�7�qqu�����|1r��          P�T'�ȿh�Y�������Ԉ�K��=a<]���&J�Yb��"�x{����FaJN�f߰:' hqż�Lp�vM|U����VxU��ί7�q���`��ݔ=B
���<�����t�z�s
           )T�_�0�wF�ѶLS�}�fE��������ow��1u�&�����̖��w/���z�Y}q�}(9��n�� p������D�y��J������+U�j_�����1y#^W��F��5د�%5A�ϊ/ۘ�Ff�.sX�8;X�W��*          ��NT�3�g���=���s6�+ŘU*����2"�g�SF�
�֨�5��OR#�ՙbd�v�C���������<���1���r��lm���-��Q��R��)�l��L8������Y����          \�"u��c��cdH��}�F��f�!�=x���_�$/����w�~�Զ6O�	             ���1�!*����            �-�HN���0�h�C�,             0�<&����0b�S�f            �=f�����P؇P�I�����Q�j            �=`��bݲ��1�!믺�+���?�ÿ             ���q�}���?ԣ�            ��#SUշ��(�Ch��we��U�#             FB�՝_��Q؇P�1����U�             ��1fӀ﷈�(�C�r�?�4��P��             ���MmMk�Q�!t�x_��<�"�             �`D���v:�Z�EaB��2oe�qI�x��             ;c�f�x��}�0
��|�k2�mǩ�             ���ɧs��=.������q�g2��ͪʙ             C�8���F�}��-g2����K�T��             �J}F�9�ҰHPDa"�Rks�,X��l��o�@             �˘ͪ�\K���P؇�-\8��S�����Y��5            �-F�ѿ۰��1�v(�C�t-��~R��M]!��	             �~1r����K�-��[�&���:Z�_���6�}ψ^�*'	            �2�F�z�W�[��v��>�B�����L�ң��?)*��            PٌyʨސN��ߨI�[�!V�ms	��곛�G��lDߡb�{y��f            @|�/9��c�S����>,E����������z��    IEND�B`�PK
     t$v[Ìs�    /   images/01119c27-1bad-421a-afe4-dfb48490a906.png�PNG

   IHDR   d   1   ,�   	pHYs  \F  \F�CA  �IDATx��|	�$�Y�u�]WwW�=�=�3#i4�[��e+�����Ƭ/XL�a���B`vp�^0�k������XcidI#�Gs�1}VwWWWu�w&��2������z�TV��|��?�����;Z�/|���N�tc؀M���5-Ð����j,Z�Av��-��.?t��/�K���8�q�>v�쓱Z�c����5�����3��곎�����z�v,�0:Ͽ���n�5�
k̪���<�E�Z���-}q�e_n4�������÷*���b����p�c!��v4t�Mx�XA_ȏ�l�ZCM�j'e{s���\���/��W˭��B���/B�Z��`w8Q���J_>�?�F��q�ܨ�����P��<^?�͆0T���E%����a��Ɓ�ga�Oӛ0($d�0�f��h���vh�\]z8��.}M�g��*� fG�.s�?_~�ݹ�:!�ނfwt�3���G�G�4�38��5l�F��������Ş_��_H/-<�s�[8�z�\�k��ƻ�?79|�]s�s|�+1D����'�S\��M���F�Q�u����5O˖�T�Γ�l����4C�X�����!T�i�e">���U�#3;��� r�*�C!l$��߿ٹ9D	�J%��6�f����Z�<�����'p��E���3E�p8���yLLL`rr���(
h�8�==����A雙�B`x���J���^<��0+��E�h��ge~������8�t:�J�0::��7&����|A�G�J��������(xB�)�?�����j5$}��� �o8�t��B�G���~�ͭX�
JCL�D;8y��-�=���L���\���w�7~�M��;�**�3 :�u�v�!�7rk-]ݏ���ڰ(}>��H_[W��7v;��.e��n�k�&,�4{��J)�!2�5��g�1,��x�!-K��Y[�Q׹�����m2��DXb����[Z甾%���K�X�}GP�Lc�>�cQ�n�
�gX� �����?��ba>㫕~Q��w�&O�w@b�t5�x��Wd�b�'��FSm�V%%��TJ��|���kS(y��S@S�p��)�#�=�B@�K՗�� ��e��h�L��BU�M������8c�0&ײ���U�h�<��G����/aT�Sr�)c��v�Ŵ�uazmC�@V��y�\9���h�TAB�o�V�^,)���3MQ��L���������_mZ���0�ޖ��@4������c�` k�u����V�#�ׇ���p�ʁ[�doDT��v�CSV���[������|
��S��\@"��QG1G��ƚHN4�n1W����}�Z���y\���qKo�I�a4�z�*ĵ�WL�KKk���F�eq�M0��)-�e��f�.��&�U'����9aT�e
BE�p����H�C�����s8��$�_�`D�Q��!Z���ǔ%��9�u�QJA��pF�x�P/^^^�W��)��g� �4���3H� ��_��f3��5"���S�6ӱ�	�@m���M�{���dM��r��L��DЅQ3�
Ы��Qj�@�E#S��$Z��]��<�*P����9ݵbY�a]��3a�ߨ�j���zS�Hk�\U�E��0��y�\N%����������?ǒ9�Q�m�9�zއr�<ޏ~��c+�X��F�D�E��E8EZ|�1�Q=s������u|��Ś'��[���z<��dʺ��b�a� !��5!a({ɀ�� �t�.�r��coԇE2�0}ۅՌ�.��-�Wkj����E�Ma���i.�v�w���1m�5�Y9�����J��<�<Ͱ�O�b�%���8�ܚ0���zՆ��$�(�� �|�o�W��T&r����P���f8e���/�������?6�ی{]�O^J�^?C8��l��`�9S:�Vj-3.�$C���{�Ȗ(r\�ms�����t
L��e! +� &�u��>�NŨV�V:mm��W}�������3K�ܤ
%�6�D��A���~���ʜ���ķR�tî��R���?$2��3T5�� R��S���p(��S߷��J��eٻ�ĸ�h���6`����/�3Ֆ&F`%y��e�$�q�%W���7�1�l�d�d	��ޒ�xb9�PdN�8�����c!WFYƦ��~Ś�g��3���iJ�Z��@��\S|м�3j-�GQ�#�c���C�������I_r��4���oX������#~�L�|�t�{��;'��&�A���!�kkO-�KL�'X��p9	n�<��!��&˄�n��Sb̸F���]��·�^����%ARvض��W��L���E��c�]���}ne�h����\��/5���>錀j��FA!1m��d��)3Z����!un�b7�o��c�5L�#tu�:��ǚvE�i[�O3��dM���s5|e�Kb�k`��nÍi�SE�X^1^�I:x�$������K�I�җ����c��:�t�M��7��P,�K�4R{�;`�1/w\?C��F�i4[�<�W6���`����A��E?!�ib�L�eݢ�$;�I�#����7:��{�V�.+��)&�rs�'�퀽���EK~Y��G_1�0����� �� 4�-�tzv�8�P�s��za�����ϡ��Ys^E����d��vR��e;�]��G�{��Ag�W�!LQx3�����Q�����:U��Q�8rНYa^��1�w��V��t��;;�Vi:~�~q΃���xj�pE���7���K��-2��
��hKc	��V_��g%A�@��Sp�J�ߢ���rw��r�1ix���s��/dU�=,afװ��|����/���l?�G��l]n��"�i0���S
�a��L��I�_�	\�{�JxP�_����s�W�dYΟ����Όn/�fU�Ū/���F������l�\���(EPu_�)ߖ-e��g�`�J鋻��i�����BA���K�1��
J�@�[�[��^׸�É�Պ���h�P�'o�nce�o��}��"g u��V���g��zO�|?��BX�ޥ]4#�6���i趽�sZ��D%�+Ҹ�!?*S�~z۽��}�J���:/��p_9Y`pR�C��7�	{�ư(���%�45�����A̷}�Ӧ,���H�6L��k|chǕ���!�����*81���f9���f�D�*V�:͕f���}oQ�p�hk0��ӄ�[��L�0�ef�RŲB[��w��gU�X,����aa��E��Gp0EIh3����L&� ��݊m乲�~�W �p�i+���0���ʉ�r\nV �H�C�)�h��?t��%��JC��L�8n ��l��*�Ŭ�6��p����!�[���~�|��423}��{��>?��|�1�u9�Ae]���!�w�"X+����������<[��Um���\�ن�-	:ͣv6"�+L�RW����Q:ն��N����0_�&V&qܞĥ�"�#T;��o@��~x(���pO��"dv��6� �<�_��	p�62�Q���XTqX8���^�53�*!�c�=��b9t���ﯮ�A�vxg`/M����Vwy����)�k��D��2�pV#�i�<�2g/ �o�D���=R��4�\RS�a^���e�ޜX��6���O�oH��)��k
�6���࣯W�I�����H?�m�!|���Ԛ[�Wmmػ^��+�j+��[����Ѵ�:^��U/�k7T��eg"A���Sj�r/�J�����e��؞�A��/�w�7�3�׶e{��%8��:�- ����^�)��X^�U&+[j�,��%�h'E��$��8�������n9���8\3�낽K��{wf{�`A�/.� b��U͐�j�NL/����*b�VA�R�q;�����c����G|J���3��X(톽��ӹ��Yx�2�1G&2�g��L%Xc�Q��EK6MU!+�������5��0���YC��Q�"�LcW�w)���zS��*f��B����m�m
�#�,��;/������X��4���kSKW���W{��d{u��-5n���ՍvL¸B�q��:�(�f:d��&�5�r�]�\D�_�X;�o��P�?sI��?��z���33�li�5�v��ỗ�ϋe�{k��C��.�E^��P�{f�Y��!�������W3��GY�'�k0=#���6��Z�a������#f���Q|��8�T%M��U�_�2���o�/��f:�Xo���;�wө�1�%fqk�CP`�9�ʪ��낽N��S&�?��0�!�O9��w�ϕ�X�q�o��JW*�Ğ�a��H"�_{���0�%<�͗��Ϟ�;�<����"7�O~㟞ŋ�)�|��?��验��0U���"�= c�H�����/�������ٝEKpO�s8��\�����a2�;�xk������qV�}v��t�ƛ-�l��KS5S"������N���z�&z����^���2���IUZzl������m��[��ǩ�e싄$�+�ҟ�ۅ�lq�]���؁Q8+.��7��r�ٹw��k*S@hW���^a�rVP��R*\����}4%�)�;���~'�t���Ԑ�m��C�QlT��ҙ)��G��W�����*N������Rk6�k���~o=6����V�c�Qe��BC�7�X"z�p�G��}[E�,�(�
��=�l�s��a��^��7	��(��i۳�j��lӜi�鲎��6lߧ�`㼉�g�凞<�r������?q����ןW�;�[�aY+�K�e�OC�$�OX.���?�iS�A��*��l�~�����*���I�}˕��������%��Å:
�*HnɠCn�h܉'jM�k�����(����3���|�\J��<V������G����w>�����&~�i������H�*{e���iG@L뎧�Y�h���x�
9��"V>�-tɪ�l\���px��,�!j�TMǲ�Ơ= �;l��z��	3Z���F4�ɧ������/���ˊp?��ĽB��X�B�q&�V�Yt�,��V�
��2!(`�)�xg��+"�d>�!��p�]���%Z��^�@�˔<��(�*�0dllO>�$���b��7T�����g$�L	�#��b�?֊L�הu���4j�Afe#U�f��|O�R�r���{s����7���"�E�i�茹܁�Ūz`�E�Ip6�D�&]�QK�|a�D���amm��_ɗ�\�¿#��"����:�Fc7��x<�_:}O�Z�s�������N����kw;�QɌz�$�8x@��xqj�� l.l���O3w`g/�c� p�{�w���3�f���X̠	b�A�8W�o��֮!�J�Ib�H�ZƠ��5�(�̥�E��S���l�g8�߭`/��6�|��d���f��ѽ0	��q���:�CG��w�"��l���$>��7�[�*x�ܩS����XtE����w!���/�O��	���Z=C�4e�z�k5��)ֲ������/*�׬�5�E�vE<�C��ү/�m�Mk��9����^.�]9�i����e��2.�a`���8q��Um5'�X^�vc��P���^�����p���R���:�u�>��x�A����O�|����g�����ދ���!\;����T�Φ��/�;k߱���wY�	�V�l�-[�~���r,")j�M�G�)��%m�-�^߾[1.1Q�Rޭ!.3E�y��e/����-��i�)��K��g��aUL�n$>W�����
���C����~��������R�jOp9�u|P:W�Bmif}j��U�3
�ejVu��A�y���`���̌	����W^��-������֓�����z����hTU�l�^M�+���_�\�`��;-aH�UE-4%z'#�80��#�6Q�d2�6.o��i��Qw;�9�ŝq��`}W���G�F�r|�_f�ͬ\�����!�� �e8�	E)�iA@�P@WK��ݶY�!s����?>�����RY�޿��)l���	:@�Dz�KD�(�Y���2�bA�5�D"��%|v���8�Mn�4s�&�e����o���!_(*)�Ő�{���g��F&�G]���t��;�sZ��^��H �Ŗ2>�)��P���Z>sE�`}�1�3͘C#��k3�)WI=���|A����JD����?�V�}�U�UG��������'.�L�F�.�Pr�ן0�vp>ݡ ����� �^J�"ªc��1��*C.�R��iZ%��!k�@7�@[q�./�|	T9hb��*H>�["���R.�q�P�9�����?	Glo=,w�р�n�3�cj�sY�����Oͮt�����ߌ��Q4�R���P�i�l�g�@ӷȸ���,��n�3zf������>/̯��@�*h��sp^��*zge&�Fs�_����@ȋd#��kߡ�n^�7H-��m��2 ��~���l���%ĮW�۴��R�M�f��SG���G�M�$����6������"Y5�2��d�N��Qo)���{���\n�� �K5�UjUo��+_���b&�2���2����!���Z�xĤi�EE1�>�ݒ1\n���[����u�� �Ί)��Z���|�ӥ>`iv��[�0��i�����pE����E6�K�^��>������b�!Lm�y2mCΟ?����TK��F(,��N��-��@��xI�d��a���I��l�Z����	Ֆ�@1�pf��a���W�^�k!A4ׄG��2�9�� �Q�Ii�H�G斻Ԅ?:�b OE���\!%�Z�ѱO��,6�����iҷ�x1+?�8�X�9J_f�4�A���~8�W]z�2琚??���!v��=5g�O�
2g/��K�e}�7�˹ϊ��va-:��gu��_�tB��#�|��E���.��O&oz�1��M�px|ΫL��|f�2�7��0��d���:*'����U5Aoo/f��q��AL�̨�y���%�>	�A��%�k)~�x%�N~�`P!��TJ}{�� �HR�U�.!/.-�o���%����f2j�nwaf]�	��>�^a�駠W+���o�\m~s�F�5?.��7X&ϟC�����BW|�G,j|H��5�i��!���hU;�E��q���Y�Fe��ڧ�j�����.xD]}bj��F4��H`�Ѹ��.�E��:؆�;{P	��:D�ꞁ,9<*�l�_��v�3�v�D�ކ�;��u�HBAvB���!��{M��?6`�+d��!�)S��B��M�}EM�����[�78��pWe9�u�ǅ�D:�"��v����v2-�ɦ��M)g������+��&�׬"���� ��ˑk�/����U;������}��b"Ygu�v�m����Ik=���l���s0�04�Lz������u�o˷�L�õ��(�dĄl�Bf��_  ���rF�    IEND�B`�PK
     t$v[��Н�� �� /   images/0657d52a-d145-430e-bb7e-5d1be0618b5b.png�PNG

   IHDR  �  $U   �:�P   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���y���}�����=��13<��!�")Q�$R�D��,q�X�ۢ���bi��.��n�E6�i�x�,�6i⦎%Yr,K�NR�(R�I��y�������?H9�E�:�|��y���C�������~�O28sV           ��B�            ��          ��0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\(�:   �h(|�kQ���Y�    �1)=x0�oۚu   0p  Ɖ���b1�    06UTd�    ""��u            �0p           '�          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\(�:   �D��~%��=� \F�icD��u�K�����Y� ��ͷD��e����/�l�����!��6�   �k�   W�ȿ�w�>�T�1 ����]MMYǸ�t߾��ײ�0���Q]�u�KJ_{�� Ƹ�'��dɒ�c   @��            �           䄁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�g    �zk����&�j���"�/\�U1PS��1XUI�IC��&Iz��(�D�p)""��CQ�ʾ����������ʾ��=���=Q{�/
�RF�b������i�����Kv�Pe1Ҥ���_62eC����Q�7��Q�{��u>@�z�*�gRmt7�D_MEVUDM��ί����u~MW_�w�F]g��   ���  �e��<:�M�s͓���!�ꢫ�:�jc�|4W�Hߝ�i�t�G]gO�w�F�ٮ�r�#��>�����`��(����q��!ڧM��ƺ�x#SV�_�����Q���g�b�鎘r�|��|�Od�X�S룽�!ڧ5D���8�F���Q�>F��D}GO�w�DÙ�1�􅫦�o�    �w�   ���������:-ζ4F{��j��H�N��$����詯�����ZU�`L>�SNuF��s�|�l��@\�p�,�̘m���ٖ�8���5�&�)�4I���:z뫣�u�{~�:�|4;-�κ�	���ř�qj��8�29ε��몢���}�_�?SN���m��|�\�=�F'   �q��   ���89�)�fM�S��ƹ�IQ*��	��诮�s��Ĝ�x}݅��u�D˱c�G�D�ٮlCdd��"NΝm��ũ�)q��1J��?��v������c��ع�~�L4�9�qJ�lT/��o��fN���'��������ŉ��⍸�������:�t4��:   `�3p  �	(M�8����N�����1=t�0�k���6���Ə����??3�E��p�	���i�qx�������P�_���q�T��B���D�����8�P�_x�SuO�<x�B�:C'   �2p  �	�T(ı��qh�8:�%�k*������ػ�6���e#�h9z&��=s�>սY��DJ�B�w��-h��	���u����ؿrvJ�h9z6���=�Y��DJ�$��k�C�̊�Z���*�H�ꫭ���O/���D�}�h�t{�   0�  �8��85sJ�fVX�:�G�d����6��ͱ����|�\��{,�y��3t��S*�Ĝ�81�)��q�/:�[�����˝pY넿�郔
�/:���W�|   �1��   ơ��I�w��8�|vTUdgLI�$�fM��YScǭ+c��S�dϡh���R)�x ���4)޾�B��W����}��t,�s0Z���B)�:��tL�������������U:�Ճ1��:    g�  `�)/đ�3b�yq|ns�qƅR�GN�#�GM�@,z�p,y�`�w�d�����s�#���}�B!�,h�#Zt>�+:���$�.h�����(�u,����O��:    a�   c^Wcm�~âؿ|vV��3n��Uƞ�����b�S�|�h=x*�a��U��Xo\�8�����޽R���=���çb��}1�`�������x���:���+f��{�̋���Ō#�cŎ��z�d$��   ȊO@   `�:;}r�~��8��5҂c��4I����86�%&�wǲ]b��CQ><�u4`{��.��B!�8Gq|ns���=����:��ζ4���/��W[qbNS������ʡ(��    W��;   �%I���3b��%qz攬�Lx�'��[��W7,�e;���]�b`(�X�x�D^4#^[�8�fM�:̈́��X{���_K_��^���Y�Ƌ$�Ȃ��E��:-�4޻����kb��b�������|   ����   ƈ�s��-�����YG�W��V���+���c����������'r|ns�ܲ"�Lo�:
����2^޼<^�qq,�u(Vm{���D��m���Wę:?o�j*cצe���E:�^��   �w   ȹ�s���-��a{�TUĮ�����Ɗߎ�/�򡑬ccH[��xy��89��y7TQ�=���΍e/�;�Gq�����Z�Ʈ[�ǉ�:?������纡   �*0p  ��:3�1^ܺ*�Z^ƚ��عee�q�����7c�?�$M����ٖ�x�U��cP������^k�{�B�t>���57ċ[Wŉ9MYG�#z��ַ�.�5Ͼ��9��   � w   ș�ڪؽqY�}��HI�q����{��[k���'���#g���LuE�r��xs��?���U�sw����-�O�YOe	��?~��Tƶ����/��O��ڲ�   0��  @N�
�x���k��,f�Qt��1}`s��2n||O�u�d	�X���[�-���P�����7���'c��D}Go֑�����7-��
͍'�S��t�����^�   �
�  @���߽6�k���td��81�)V?�f�ܱ?
�R֑���=-��gm��\�u��#���ͱ���bՋoG��f	����S����F����pY8=��k�k��k���u>   �'d�   �,�K[V����"���p5����-+���9���;cډ��#W�`Ey�ey�y݂H�?���������������t�=�H�U2XY�]����	d���6-�C�̊��+����:   ��e�   9�pF<��譫�:
ho�?��X��`\��Q�:pY8#��ku��Wg��O�?�ږX���㆟���a�;�`zl�{M���	��iR<��-q�+�↟�����#   �9�   p��WWĶ��ġ%���B�J�B�q��8�pzlyh��}a�*ƶ������YG!ci���5���������hv�/�;���q`�Ο𒈽k�ű�M��G;���٬   �)��   �DrbNS��[[��y����x䫛c�ƥ���� ����)��7���]�5��W6��-+���a�8=sJ<�����GwCm<��-����F��cY   ��	�   p�
I���}��Hc6ޯT(Į���������KQ�ѓu$�c*
��%��&7�pii!�=ǉ��b˃;t>�a:��I�$޸~a��95�<�#&�wg	    �    W���u��7n�]��sY��y����X��Xm��7t�2NO�~�8�lv�Q�����6��|Hgf4ƃ߼-����    �c�   WБ��������2XQO~v}<��(K��qtAK<�qv�䬣0�V���]�|o��Xqb��x��[���#�(�����    �S�u    ���=��˛W8���m�y�1�.n}�Ũ��:�At>��B��ǭ?|1jz���|�w;��Nm�cۻf^���[�=ߛu   ��q4    ����b<���c疕��|bm��⡯��gN�:
p	�����oܤ�m�S��o�m��f����b<��:߸�O����x�k�F[봬�    䎁;   ���ƚ��W���-YGa魯�G�%,��u��t7���_�GN�:
�H_]U���M��·<魫�G�%/��uƑ޺���7����   �+�Y   �����)��o�}5�YGa)+�S����kc�soe&���'��_�1�j����8T*��O�����X��[i։`b;���}�譯�:
�P�P���^��c��F�*}    w   ?�ff<}ߺ./�:
�Y�k��T7���(��_ ��̈��!��:�+�b�w5����B��u"���.h��}f}U���8������*6��(��   ��f�   ��k��K[VD�$YGa�xg��譫��~�#��CYǁ	��uc�m�t>W;�s�gRul��Q1���jzs�x��k#-�|��C�̊��ʸ��u>   0��    cٞ�cǭ+���o�yS�WWd&�=ǋ[���\u'�4�|���lX��\m��Uwrδ�_S�u   ���  �ǑD��uU�ܲ2�$L`g�7ƣ���UYG��-��q�J�O�ζ4�#_�}u:�����|2u��1y�����   �e�   U���k��u��N�1mR���M�[_�u���n�6^[�8�$�S���l���ڬ���t�&�]�e��sj}�諛�K�   ��;   |i!���]o^�0�(��S��6GOCM�Q`\I�$���xc��'?�k���d��-�xnb%W�j��n1r   &w   ����mw���+fg�ާ��&��M�WW�u���w��wV��:	�OOCM<��Mnl�Q��U���yYǀ�驯�G�%���  ����   >�����k�e>PWcm<��M�Wk���K[V�[k�g>PϤ���6Fo]e�Q`�۹yE���vr���:~�����|   `�0p  �a���������9�>~�śc���u�vݲ,^]�$�pY�'��O��)�*��c�ƞu>���X?~�ͬ   ��`�   ��ʍ��0��kn��~�.�eƜW7,��7-�:|h��&�c_�9�*ʳ�c���ŮM˲�Z��x�7�`��Y  ����   ~��f�˷,�:|d�fM��}v}��$�(0f\�/m^�u��NO�?���(��֡kfŎ�Vf>��:   � ��   ������E�3FY0=^�uU�1`Lhk���w��g�:��%�ݹ:�0&�����{}���gl:6�9�ݥ�  ����   .�sj}<���b�̏Όmo�[o\�0��k]�������|Ƽ�Wϋ�nX�uȵ�ƚ��n��bY�Q�y��y���%Y�    �"|b   ����2~�n���b�Q`T�x۪8�xF�1 ��k*�￴1�k*����[W�ϯ��uȥ����7F��g��yˊ8��5�    ���   ~I����>�>�j���&-$��}�cZ}�Q WJ�B<����ը�?��B�mi�:
�JZH��O��'�eFO�̽���铳N   0��  ���x����:-�0�*�������YG��x�֕qr��g�./�'>�>��+����s��86�9�0�F���gu>   0��D`|H#�#�h�4:"�#I�#M���Rw�WH��H��4��HJ�i�tEDJIW$����iIRJK��$I�w�KR(T��imDD�&����[QJ��$
�i]Ic����Dc�{. ��:�|v��vA�1��9?�.�������/���e�����Yǀ+���6������l�$U�Ll�όWoX�u�bzj���w}��HJ:  �z���4Ҏ��#��H"�(t�Q�.�Ig$�p�:����eIғ�J���}��kʓ$��.��")�'i�!��L"jJ��&5Ic���i�Ic$��H��ph. �3pȷSq4�8��q"M��$J��$9Y(��JIr����dr�PG�A?�t��i��Rs!ʛJ�Ҍ$
�i�6%I2#��%���1%� ����4)��{m�1��;�hF�ٰ$���v�Q 3��&ų��|ƿ#��+7]k�+�(���)��̽�E$Y'�+����ؽqi�}�ͬ�  L�$�dq8I�h��Ǔ$9���RĩB��I��U������1Nχ4"��������P6�\J�IMi!mNҘ�F2+�h�H�FDm�y��2�Fz2��;��$��i��$��H��,/?�:ԟu�і?~&"�\��ҙ3k�tn!IZӈ�4
s�(-�HFĢ��y `�V�����Ų���;Ł�RM�`oq`��|h��0Rj/+���ᑡ4���~_!-U��k"��Ჲ��Ų�����ʚ���b�X$���7-����1��鬣�U7TQ��d    IDATO|~C�5:�*�K�}}��C=�C���FF:
��y_�GZ5R^V{����e�F���j*k�t��۽qi4�h�Y۲�W�p�<����,fe�)��.���Hi8��|�����4��Hy��b٤�bY�@uEm_ue1-��Ѵ�ƥ1�ع�}@� ��4�8���/�d��q����iz�j����ΝCY�mIDmm�������M�̙<X*�����RDk�&
QZ�F�(.�:��Ff �'�� \y=雑&o$I�F)�}I!�Wܟ�>ݝu��J�7/^�Λ�840�0M�E�$Y���2"�FĲ����Q�q`�����&�cZmw�`mg_[U�������#Qz���l�o���~�?�o��튩�^[W6��`Uq�@U����Yݍ5���'�~i!��?�.>��Ge����#/�~m��\�u�1�����|頻�����������ݕ�F���r})�q�X�8X]\�W_5�|C]]����H�$������_<U�Yǁ����VE����c�i���Cu]�mU��oWm+o�o�����W�=��r��O����m�%##7V7TW�꭫j���_�ܽ��g�≨�w��  \)ݑě���I�o�"ގ��}�t��=y�ĉ�1��Ç�#�="^�ԯ����*Ǣ�PZ�F�HҕI�"bnx� ��Μ�f`���7"bw��I�����ЛUmm��]{��e���RiE!M��I�*"]K"� �X�ߌ����Y��@�_�j�O=�u.�������벎1�L:��]���jU��c�e߻�?|�������ņ©ޯUW��S_u�����R���G1w��������+�ݻ"����qI�]1�����1�Z2+�����c�9�==�=�V��4)O�wǟ������I��ů�?�;�zݹi�ZF����Q��w"��۳�1&��Q��C��g���/?�u�1������o�:Ƙ3�������������J���?{譫����3�_�,�LϤ�ڛ'5�Y������O&r���'"Y�$���:�7e ����p�ޮ$�גR���~���ɟ�t\]iSS�PYղ(+�H�dYD�I"]�|c�L8���鉈=�+"��Ȯbm�kɾ}���X1G���D�߽�����v����4bM��ڈ�u��p�; Lh=5���Y��FJ锓�k��TL��������Yg�������O���kLϏ�����/�mnX�_[e�x?�ff�}�X��P�Q��뭯���Y�u�1�l��Nm�<Rs��G�������}ɧ�]M�~����.^�ȿ����������K�W��V���8�hF��f~,�}0�(p���V�s�\�u�1�0R��mG���=R*+|�?��׳���?�+"�{������G���U�f{��սu�>߼�#Z������ ���xwӑ&�"F^��ȏ�����q����Y�Zi��,bmDamza�>7�� d�@ �W�HފH_�4^�Bl/;�Z1�u0>����'"�]�"""]��b��sM�bCDiCD�!"e ���BO߻.+�YGɭB�S�:��w�����)���幬3�:����uD��E�����X6���?묮��ggNY5PUt��xq몘~�LLj��:
\1i����]UYGɭ����S�:{��������ÿ:�u�_������������[w��O�&U���3����l�m�bƑ3�p�+�(p�$��{]�W����Ҙ��q����o�$�����Ne��׹8x������o6���������̩k�+t�xi˪�q�LL>}>�(  WZoG/D��ۋǏ�I"���GSs��ш8������e��|C�$�4n��uQ�UF ��dp�,�Xx���؞D�tDl+��z19p�3�P\���M#eeF"nJ���#§a c@�ߌ����Y��@�_�j�O=�u~�k�Ŏ�����KU�CSN���ߺ��*�?�'���J}���h���3-��F�u��i:~.���OG�z���{WDS>�����ß�?�c��/�n�ĎK���r��g�I�����ￚu�O���9ߔ~�����i�<M�_�����<II���w"����qI�3����:F���f~l��;.��w`h��O���o��~%�<��K��_�3%��;���Ӷ�M3҂��USNu�����(��\)�H�,�:�%�����MY� ���H_L#y��&ϗ/$��g��#�(lm]��čQHo�4�DĜ�s0������H�+D���g<�j�JN�<_�"��������&I��H7%�l�H'e� ���jc��eY�ȝ�s]��:�����߾�����yb�m��������O}�S[�����ZV���e-7NϜo���v�:
���I5��-˳��;�v��k��7�����D�u=�����WsJ����:=}r�q݂X�������뫫��[Vd#w�����Ϳ��?�롬󌖋����O�S[�O��ö9M���Y�_t��!^_�8V��v�Q  >�ވؕF�l!���&��g�l$#q���jD|7"�g�����$�H�M��
�Xf�LD�|��OӴ�X�䑗��q3�at%;wE�΋��+VT����w$I��Sr K����^C~$~״�G�ۻ~�?{������|��'"b����S˻k����o./�FwD�ܲ<��;�]}YG�Q��51TQ�:FnL;�~��l׿�����_��l]A����5�������=9o�ơ�Ώ�x���1���Q�ٓuU�߹&+u�����8>�\׿��g?�ˬ�\i����S�n��>�����'�6m*u~D�޸4�},�;t> 0f�DĎ4�BZz�|���?��K�=r�xD|����f�����;#��#�9Ӏ |,>�&�W#���䱲t�餭�;�|,��F�S��M�̙<8TښDzg$�]���# ��o��86�{�S�:O6���_���C�u��m�_<�FDܼ���-ko�����6�)/d+SC��vך��o�eF́��Ȃ��c�´�ζIg��֝`���n��z+"ny��.97��{�浬��'��c۝k��������}��Y����y�����lz'		�"E�����+`A��9^_�=���z<�
R�J��&A��FZB	)��y��^�}����9v��ٽ�~���|��~�\ܙ����N��y�<iY>G;�$4��w4t������w�v�T;�^���𴥻k�n
��<��ot�z�S�S�xJ�j�   �E�E�ak�#~"��in����'�֫���� %"׋��V�d��}�YkŬ�cD$�[ �,���QyJ�y g�wW�a�v�ɴ��ȝ�����Z�O,�?K�=SD��� ���T'���PW�742'��?k���r�mG߼�ey�����ƾ�����5--���.�-;WΗ%���S���V��˓��PW�?42;��������-ڎ����"r��qXOS����7-+癟�g�l_�@�ni�N
6����|���t���k���v���7�h���~�g�{Z���M+�y懋f�k,��/��N  ����yΊ<`l�~?�ޤ�h2"V��YyVD�b�ϯ����YF�۬�<�F ��ǂ;�Ȱ"i#v�y����vhH�����E�r;~�x>���Y"v��4(� P�~s�~2���3�xc�����w�f\��k�㕮������,{�}�_ܶ`���k����<s⁲`{��3Y�� ����V����ع;�n�=+vщ��7��SJ��q�&Y�ąg|�m�����ꪵ�����e�km�s,�۞[���T��|�x��kf�k�����{�|w�f��O��m��o�5��h7i���d��P�1f>  P�'b~d%��=dR�� ��J��ȣ"��xf���m̞iĞ)"�*� ~� \�"b�1"�{a�ш��������."�[���ܹG[�s��s��K `�uϪ��\����)ݛj�>m�w�ެ�Rʎ����?���O��yŜ�d���q�&)/�\y�e�`���je�A�;�g�{�u݃�N���[J��7n���'�pcӲ��w����W�3?!/�B{����?�V^9d�v�f��9���tǹ�޺���]+�;�ye7�G�����Ɵ���  �K�ِ�v}���!�ed�d+m���_���G��]Xacoc���E$�[ �w .�j��i��;yM\aDr�O��SV䟳��k��s��sx�  S�k�n�A�㹹�:�x�UwQ��k6n��r���<��pɬ�{fN��n�j�߸\�}a�T�k� ��|��~J�f��[ڿ|����v�+�lܘ��r�O߹���ų��U_��4ն�T�}~����2D��'$�X9��3�9��q�w���v�+�[�>'"�?�3��\P���F��ҡ�ȊgwJ]�v
  �0#X1w���O��4"9	C�2௫��\D.Z�`��˝#b���D�B� �O����U�V�W���0X��ϲ�W���Jm����0X`l�8�JD���  ����m�t�)���߶0ݻ����Y}��?Y��KM+^l~0��k�L�l�B�9� �`BZ��#�3�3�\S{���m��>1����o�vKӾ�w=Pn3?W�gN8P;��֥�%X2S;c��n��>1�߲�goK�:c�K��T��k��c1y�Df>  �=b�jcc���`��>�R�g�pLukk���08��f托���/�� ��p�;�R�#V���O�>eD��f�#b%�~RD�����\[�)yk�%b�,"��}  DA.�_�J;cJ�rV�oOߺ��w�o�X���iSF6�O^p��w-�w�Pm�l�Ki^1O��7ɬT�v
����[ԍ��`{��S�u�;���1�%'r�YO����w��󽡺ʲ���{0dNK�v
���1#�ZS^�1��\*y�{������uٜ���<����!�d��v�  �a�//��DC�Cf˖q� `2���v�BD�]�`iE>�Nk�]"��r D7�(5���]y�g{�s�t�a/��S��Q̦M�xl����^.;�Z�yT�� � ��a�N+�����%���v�]�a�x���G�[�y�Aw�v˔1"���_��+[^,�e4��2�E[�����og�����y�o�/���ݡ�2�~}�"F��s�\$����S��?9���G?�����٭]m�-Si�q�3� �DY��Q�\�e�g�a��d��r;�E��u�_��`{��\D�% &� J�b�^>7���� �;��>�H�n��`m���1b?/Fvhw ���W!/�B;c�4t��[��y��W��]�(:��m]��E���h�L��y�%X2S;�#�xL�?�|f����K��r�w�Z�%��gc�[�/���\�H�f�K�>��3�=����s�|���u�%7���2�g�K��9�  �-���/�s��t����Lg�v���g� ���P?�Z�6+�d��  *Xp��W�|Kl�p?���7L[�A�He:���/zA����1r���hw ���Y*�5	�)1#�i���\t��w���e��o_w�]G�x���X�<�_~s�*nw�^y��IjgL��aO�����_s��-Qv��M�uW���/��^,_/W{�����p�փ�P]�vƔ`�O��֯ϝz�]'����oVd�c��f��bC  �Uc"�6#v��$����-\���e�x"��+gy^|��yU� \ǂ;��g�W"�����~����No�N\`D��Jm��/^1O�|BD^�� �Te��l>r�vƔ�������]z�7�[��\�p��|��s^&�-��o��vG���W!/��vƔ�������}�^��_��\�p���i�g��l�g~��zٵ|�v�We�e�Ǝ��?�j�%���s�M>�ߋ�K�E���;�N�W���   �i����w:�w{a��)�� ��]��^~��������z�hw���� �ƨ�_�^����1��LKK��|CD�1>g�a�}H�\ "�q]!  {�Ö�h���1���~`ݷ�<���H1���y×��Ӄ����x�Շ��R�H�D~��z���2R�-����Ӿ�����%�g��}�iY�v�ƒQ�������b,C���7,��2xcǢm���֝�kw���7>x�O�sz�c��;�*�H_��ꕲxk �L�N  �����������HN;p��?��ؙ3ge��{����b�4 pF���P����y��l/��B�ہb���M~\�e�%�ȿZ��v  �r�|�>��ˊ,ږ����vh9�o�����K�E���Y��Z2K;��r1y�K�3&ݼ�w������Q�V���[���s*��=�{��$�t�v�g�cF��1�oi�"���?`�]�q�<x�gw�U54�Ů��Ҳ��5 P�:��/ecf�kA���v��LGG��.��`Y^�E�1�& p� &�cy�g{a��SW�;x�*0�Lgs�_��[k����n @˶U�"����}��wkw@����p�]oK��E����/��Y;�_(���^��������w<vϊ�Z�NG{�}33%j���e��R;cR-|-�uݕw�C�"���ȃK6���e� �(zQ�^����D:�תT*��Έ�ax�'ۘ9H�|WDF�� �T��������6f����d�o^��)d�lO�S��a�F������"��� `��-�G�&�E[������;𿎼��{�m�����xd���E3�{V�v�����7.Ӯ�T������z�v�ב�ڰ�]oO�Fw�-�.�s�3�?���h/�.��v�iW�����cn��}6������Ms�}�t�  05�"��o/+<����f�k�T�E?L]������"Ҫ� ��w ��m�|����ApA"�zA;���tz����"��"2�� �dk]:G���jgL��;�]w�o����:�և������D��Q_$�{RKfI_S�g��s����S�����?����xt�'�|83�%\4SzfN�Θ4�w�?~ڷ~�f���co��˷�^�e2�}��[� ��1{m>fV�a����F�l��47�����^C�21�>yY�	 J� &̊m�b��%Ka�󦭭S�	��W�����G=����/�H�v  ���#���53�y���ן�݁�l��_�����|4j^9O�ꪴ3������.c�l����U'jw�/[����]�e�c�h^�k߹2P_����(��Y���_��$��e�o��-K7��[Tg~��ّ~P �26 b��Y�ᇒ��k�A �<�e˸7xa�*/�l��v hc��Dlk>����D�����ѯ`Ϙ0�J��K�\v�o_sբ� @1�̜&��3&����Y͙C��f�Rw�-]�lK��ɐ���Ճkg ""��T'�3�3&ECGoUG�A�^zi4��"���e�[���6f��7,�� DDdwC��gjgL���������9痾�o|�K��ܬ�1�1���K�3  @�tX1_����0�XU��� �#b�ax����c��� �)���5o��`_?���47�j���>�S�{sf/11;��  (��]����1�7�_?�݂=s�w�?s���Hވ��A�$�+%��z�b�IQ98��vz��i�`Ϭ����ߖ~E�c2l;���Ұ��E"F����F���a��k�`������a����3� p�	D�G=�[�S����^�& ��S�08K�f��#,�(3|K`O�(F.����D:u���D�ٴ)㇩�9�V��E$�KX ��WȎ�hg]E.og��8o�uwqˎc�6�k����(��ꤤ����@��U�d�����X6/��߽�7k�`�,mi;bz{o�f�HUBZ����@���b��E�E��eގ�w���~ް蘪��GMo�ܛmG+}ٵ|�v  ��v#�x�,���7���?����[m.v��YDx�#����;���7V�[��    IDAT�08���$ �̦M?n���^%b�/"۵�  �[�+��X���(�����^{���jw`ﭼ�遹���K��E�!ᨾ-�صb��V��E���o�pÆ���{+�{z`������X�?�zp��ᖖ�sd�*��Qt_����~�݁��f������C��|  ��U���WU��S��T�7��ho���b�Pc�.�R ǂ;�?üd�9���ax/7�������0X)b>hD�) ���oX��PtsZ�^>��{�E�w�]�<����3j��J-�%CuU�(c[^��Pt3���\}�?iw`⎺k�/�oi�R�f~�x��Wkg��E���9���O���Ohw`⎼��oi������3dwC�v  ��:D�Ǽ���~^i�m�0u� x�����C��� �,,��}�b��^�:(�N��b;P��H�S��ꗊ5�H�v  Mc��ϛ��QT5#�U���hw�po����.����vG1Yc�U�3P��%=�I;���G3��Ǝ��@��t�C�_�-ܢ�QTFd��|��V%��EU50����o���-|�m�vGQ���w  Jؠ{�7:��SW���7?�K���b�hy\� ��w ""�"�^C�2?��ƈ䴃 ��e˸�N]㍎�k�|AD��  �sv����PT�Z����'_w�E��W��j��2�����ܱs�<�]Q<�Z�����]sWZ�ű(L_�;8��QLQ;k�;W�k�3�2oW�E�󣣾��i���Ŵs��H��  ��+�k��ŉ0������P:� ��'�b�yN� ��w�����2���0�M�eK�~xP<��gw"L]��sKE�7E$R�Y  �Em�jNs�/�^w�M�(���Yǲ�Z>ilt^��;�N��j�3P�v�@;���tn:�{���@��w�3݋_	?n�љ�����3s�v�Ў����5w��D���rԭ?ڽx[��X>��R4�U�5�^;  �./"�gcfy"L}�A�v��O����0+�]"�K� 
ł;P��b�fϋ/������sP;�L[[���9����� @D���N���3��jp4S32z�v��;�b���W�;�i����	(3����;#:3�rh,[��8C��w��j����bb�c��WI��팢��T����݁�;��GnY��}�vG11� (	?���a���T*Ў�#�O���^C��b��E�_�	 &�w��X1ۘ9��̮]����$�`�發9A�D�� �{�#v���]�]s��]���[��U�F�zǝ+���C��;Z;.=���۵;09�{�UFh�G��ҷs�|�]Q<��mfg�i��Y�bٹb^�>  �ż3r�'�a��v 7�-[��t�r/�[."W�Hd���|�����D�:5�J��] ���^�:B�\`D�9  �"J�VMm�����5�L�C��ؼ������?=Z�i��5G衊��}k�s;0y�kcj���F�b�����ѹM�/J3F�'�m���s���U��24�J:�4jg  Pn����{a��xlЎ������b�V������;}CV���i�x�ԏ�c D�������}��/�Șv �|�7�Jc�vFQ��y���{�v&_��m�޹{X��Xv-����21X_�*L�Jc[���|ǎ<����}���Ҳl�v��pm�tϪ��(�X�J]��{�;0��ܰ�c�����;��e��  �E^����s��A��-� &A"_I��3�ص"�v �	܁�b�&/�-K��K͖-��A �̈́�p"L]�7r�5�#� @yH�3S;�h�t���|D����M�2s��]��Q,A�>�(m�Kfi'֮͜�O�~�C��|f���mO�_�bI-a�S�uitf�ܖ�_��������3"vNk�'�j�Gj��| (aO���� ����uj� �>/�|�Pc�s"2�� �@4=g�秃Mgs�v����� 8=/�l1�C� mAD�cټ$GF������uf�ӫ�Q�se,�kg�Yv��奦w���:G������n�b�=MF��(����㹜��d8痑շ<t��;���̘&#5I�  "Ɋ��ȅ^��s�= ʋin����٘Y!Fn��c� ��w R�n�Q/���)� �-��{��ʊ����	 @�e�Ҿ�I;�(���|���}I�Sk�Ύ����m�Hz��D\�"&m�1�g��|f���u������H�|c$��7w`r�cF�E��lvs�S�_y7�~/3M����oD���x� ���W��#+� �ɰT
@QU*�Ap�{��l���?Ƃ;��3f??L}ӈ�{ @��'a�o��� b�� ������Whg,��ٺ���;0��X��U����bh݇�L���3$�ǵ3
��2�=_�S����}wNkW$^7���dk��$����l�Vr�/C����g���b`� PT�;�Ï�����1 �;^>���A�ʗ�������Z�6/�[��j� ���H�_���1r��D�} ��pI4nu���y���mء�M����n(�p	�/�\aD�0;�~��o߽U�:f�v��vC1��g��
DY���Hu?��7kw@GC���j7Cz���� @����K�08�O��Z; ��J�$����1s��<�� ",�.�Z1_���7�Nݥ ��~���s�����=  ��-h�N(��V������?;�G�;
5\����j�DX��,�[���3���������?��Q�Ѫ��7�jg ��L�N(��V���>��=������}���:���o:3 ��2"�eŮ���eF$�� K2�z���"�"���P�Xp\dd���щ0�i���(�����N?.���F$�� pS�����N;�`M���)W���v�;���V�bh���2JS֫��YӴ3
��ޛ>��{����;3�u�vG1��k�N@D�*b�=�A;�`3֓���g��5���;���9 �	�b�����°U; ���~~7S;��ܧ��|���%k�^�UVΫ� �.�J=Y%F��� pK���1�_�^�;p�v�-�����Ș���y,�`rt�n�|f~]�෵�o��ݟ��kw�eGL��������Um��7��/�:��ʡQ�oj��� �^�"d*b'��m�- P������7[#�H�v������@�xQl��D^b�mӎ�b0==�� �����"�M� ����Z98���c�"~��٭�[�;
���%JS����c����W�;�o��O�Ju���Q�(|.Q�:"��D��X�b���зf��љA�3���  �1ra"Ϊnm�c �XA���eW���- ��@����zsf�ӛ�c `2x���^f����6w �����3�z[s�ƬvJCc{���n(T��:K����������'λt��vJCS��E��廻�FF�������	�vs��������3��ZFj��  �4#�������[ `2���/���m���= ��@i{El�M^~�lڔю��d:;�t��F�:#h�  J����{|<�%���7������~[��S�]�����u�!�a�>qwC��펂��9�/"��tE�����]�����?����@��PQ8� 0I�Ś��08τa�v L�D����UF�~� �ǂ;P�����e�ӭ�֎�����q�;@�ު� (M�u�2��3
R�38�������@i����s�B��`��5\���J��P�74|���<�݁�2����s@��i�	��Ѫ�W�}Kt}���I���3���Ʈ�Οzf�i'  P�ˊ=�O�����d::ڽ08[�\("��= ��w��X�m��9���M{��v h0��}~�緯���� �����>�{�'�(=�}_�]Q��&�?�(-QX�m����vJOc������P��g����G�Pzj3_0y��~�Lf>  �gԈ���S�°U; ��ApS.�=H�<�� �XpJ����O���R���9���" �����KE.������{rôށq�B���b��m������(=�ܳqcC���vG!���!JKf~,o��݀�s�m>W�=����Qx  �"y����^��̈�c @[e{�N/L�h�^*"9� �;PFĚ��a�v��ܧ ��2[�0�ƈ�DD2�=  }�/SU�����=�;P�;��h7���V�1�nB��:�LU94�Y�kw�4�w����P�ݍ5��3�Q<�?(W502~�w�zZ����{`�vC!�%�ŵ3  �e�fO�����) PJ�H��/H̬1;�{ D�>��K6f���)n������0u�9� \_p��=��3&Wm������b�?�F;�;�����ݯ#V����g��B�c1����������v��݀�U58|�vC!�1���9 P������Ap�	�a� (U~*�K/�""?�n,��̷=?~X"��o �~���F�=�-  6fd���ի�F��n@��<pU<��[<w7��E	1"����{�y@���>�:>���ʘ�(�ݮ��G���n@�J��ucb,��Co����	  L=#Od���P��bv�����"�EdT���Xpt�[k����?��f�c {��R=^�z������k�  ��pm��cF;c�H6oo��@�Z���4thwb`Z�v"b�:)���__�<����h��O4v�kwb`Z�v"b�*!?��1qV$f>���7m�L����(�| @��[1_�प Hi� �k�0���̑"�U������p�s��9<�Nq� �S����٩� �:���^��=����o�����W�
1Ȳ#�d��KTU#�~�N�?Ϙ|���[�
1X����c��s~�S���U���z��s���V��  �T��͙�0�y#���@Q"�z�;\Dx�	a��R滞��L��i� @���&��7Z�?�n L�!�gk��Yn��T�?��vC!_JF�r|���ox�vJ_��ч�
1X������s~M����������� (�̉=4ޖ��v D������b�"����܁�1*�|�S���Q� ��~�n�\"ܢ  ����������(}�ãh7b���d���o�N�;}K+�F]��{�
1����c�����k��>/g��]1q��i ����5^C�q�aآ� QbD���!��ji���܁ɷ��̑~:u�v D��^��̈=MD��{  �g�����O�P��p�OQ92�����j�]�(t|ٱ"�yZ��o�G~�|��X^�c��U�5}��Y����ێ��G���Ѭv�D�UJ>�O� �H�b����f˖q� �*���W^>w��<���|L&#Ox��щT�� (^>�{��٤� �#�	턂�T�N�̍�aD�=����*d���3#5n�|�{�k'��[�?ԯ�1Q�XL�*}�D����|+���ޠ�7��r�r�|,&��| @�������k� @90mm�^��b/�nP�Xp&��5/N2mm��- PN�°��e�7"�[  ���鉑��Y��>����#�vC!XvD1�&��;��2����s�vܐq�|��G1��wT9<�=���۵;����x�vC!\�� �g��{��n��v �#�K��%b�"2���t��ߨyo"L}ʈ�c �����x�݈�D�� )�����X986�� w$F�wi7��QP:F�ܝ�U��C�pGb,Ӭ�Pf>���s~rh��7�`�Ud2N? �� D��k�9�י0��N�r���"�M"���! &�@q���կ� �ɈX/L]���E��׽ ��X��?�'��y��X"�}U��./��t�|Chrt�[��H�����P�1f>��噟�p����m�n(3 cb�~\l6m�h� @����Y/�%"Ok� (=,��b�/���o�S  �+�J=h�7��oG ��*b�����e���{^��./��4�c1�=�	��2�v��d��n(���`Fd<������V��Ì��Z���� ��4bO��B (-���ͫ�<I�ܢ��������C��5���M� �mm/y"G��'�[  ����\�eG�xF������+�%=�]1q�L>�� wxC#�h7���B�%<������d8�c�y�8�֎Q�ߪ ({���!7@	2۶��Ap�X�q�k� (�~c�{E<�݄�v	 �/3A��UV�*Vn�n LL��|ED$cYv���޹M�v��e|w߶�Ґ�+�
�	3{l�kۍuw�g=�?����[�DD�9˂;����5�wwW���+ �l=���� ت ���t�rk��"� ܁����0����1 p�ٶm�O��/ �)s�*_�I6�n�;f�rs�?��Θ0[�����n/̚\�eG��;�cg7�]��B_��ퟪ*�6�� ��#g���s� ���5ޜ�g���>� ��I���j#¿��2������^cc��A�-� � ?��܊9_DƵ[  {.w{y�X�m��cF$�:���s|Q�\��ۦ� �0�Q�\_p�Z�Ԅ��gs�>��� 8$o�|���ͦM��� ʕ�em�yY���� ��	��/��S� ��%��m��:��n ��H�V����x޺��s�����ݞ��|~H�n�����|n�E�\?�W�<�|���9;��� n�b���࿴C  W�N����E,;z@�r�[C`�ٜ{��k�  
���6_�ZDZ�[  [���|��a����rV�a��/'C��I+�|�
��]�}�r1���Ɠ��|�X�ݙ��C� ��0`Ğ�S�i�  
gZZz���SD��- ��B {�q/�8�*Y��I��l�TĎ^���������fG�X��&���X����Y�`�c���+�>�A���UX���^1�f�&�s> ��Y��9�Ç�[  �c�m����V�W�[ L-�� ����k�_gv���. _ukk��+ֈ�'�[  ѕ7�_M�)����"�z=P(s��#��`���*,3e�0� %˼�{��i�  �ψ�D���s��mP6�q�[�|�S�1[��k�  &�믶J�5b��n �y����Y��H>���n�[l�8{%nE��Q�X��ˬ_7���N�[l���*�n�Ѡ/�u{�g�1f>��5&��0Q1�� ��d6y��	Uaت] �\^��L��WD�}3�=����T�b/������a ��m�X<���[  �"���6^��;����p�6P�ՠ���Yk������pw���R��"��ߐ?:���^ɻ�P�| @�1�7:|�ik��N L?n�b�NDF�[ L.g�@&�5F>��K�C  Sˈd�0���\�� �C�/O�s���%3�~o��r2���<�q�/�N��w�ځB�~�ϙ�|��pv��8� J�s��y�LO�n� ��J�����""C�- &��_� �('�\��i�  t���`�� ��X��ҭ���p��e����۸��}1���ab2G�nOx���G�\���<��e܏{��� �{k|άsMs3��@��ҭI>�FD��[ Lg(&I�y��N]� �煩�Xr����������pǮc�����f�����~�)�`�c����!�pw��y�>��%c�c��K%6�;� ��o� D�U^�o6m�h�  t�m��#'�H�v��s�`�[kޑ�;�C  ��S����� @�?����X�l�����v�vC!��v獻�0k���� w��Y��5F;c���?�����!_��c���<?_��̯p��j ���/��� �� xΊ=ֈ��- ��w�ucy��H��� �?���, U�ȸvBAr^|�v�1��Wh7"9:�� �%F��Xw��y�eG��@�G�    IDAT��J�B$��>�A�?��X��[���
���c#���
�� �c�|�O�r; ��%��ؓXr��w�����ax�v �t�a�m�!q�W p\E./�÷����y�pG&Yq�vC!,;�@&o�sw����cc��vC!XvD��H��Y3^|�vܑ�+�n(5 �X1_I��Oiw  JW"_��ǈ���- ��w��a#��dާ (}~��N�|@Dx/ (qy�e,�7i7��~���YvD�<��+���pG�����g��忣�Jo�vܑ�ܾ�=�9 ����b"L}F� P�*��w�s��Ed�v�±��r6jľ��G�C  ����1r�p�; �H��{��hM�F��Kz�
�p���ґtx�q�:Y�� w�'����H���YE�p��_���n�;2	o�vC!��~V n�"��S���  �#�޲#�ˮ�V� �a��j<f�\�� ��"��; L9�ovM��|�\���1uF���
��g��忣�D<��ߺ�v�0\����P��0���p��3�:����7�T%k7"9��g � +_O���ig  �S�޾33'�P��ı��r�ɋ=7h�  ����Ě���n�rR94��P�����(}V�b�����㙜�����U�j'�����(}V�4TM��\��|QU���k�����#��*�k7LT,o�~  �#�����hg  ܕL��匬�"i� Â;�MΊ=?��i�  ��S׊5��� �rR����K֫8N���7��Ѥo�;&���G Q5���
���c�P�^<�CG��������b,C�s�����݀���w��h���B�c��w�H,�- S�~��֮  �/[��5Vl�v��ǂ;�I�yW"� �?��܈�D� �EmߐvBAƪo�n@��N:}��n�?�(�}n/��Uyi7��Ψ=[�����P:\�[K��j7��zr�8�H�H�| �T�r��3\�  (�d�j�Y'"=�- ��(V�|8wh�  ��S�Y#��� �f��eǁ��%�(}�uU'k7���5��op�o�Y�݀�7T㟢�P��~�?�(5n����n@��L�� +�| ����y��Xn ��K̜&"��- ��(F�g�0u�v  �A�Y1r�v D����V&��m˵;P��Vh7��D;���#�I���@��������
���((5Ο�]t����<X��՜� �����}F$� �&?�z�y���j� �3,�#�/{a�U� @�yA��"�}� ������ݾ�'f3�k7�t�v�!3���j�;
Q���R2JG��ĳ9팂Č�[��k�ɇM�Q[��Q�>D�H���7��Θ8#Rab���m9w��7�v�vG!�8� &���3o6[��k�  ����Xk�-"n��	�uW%���#  ����9�/�"�[  �L�J]πvFAF�+��n@��7���
팂L���(+R����Pu��(]]3�>���������eZ��˳#5ɷh7�t�T-~���Bp� L��x�-&��U! �)�H��+��o�� �0s���] (/fӦ�/�<yJ� ���s�vBAz�j��n@�h�>G������(-n�����֊��l�<�uU�j7"��˴n�Q<�}�	�^�J��k�2��[]L�ʴ.��e �����eך��^� @y�����ȧ�; �u,�#����׈�C  �Ǆ��8[ļ�� Q��ٯ�P������<I���wƴ��
1�{@by�)��i�r|�W������(M�Muh7��gH*r�|O����T��|�-'hw�4�M�9L��u}���3  bŶ�r�u���C� P�� �/��u� �#�=��;�e˸v
 �|����lLN�V� ��op�'�n@����ǝ������(Dc����(=�?�$"���?�݀ҳ�'��^���(3���[;DDr�Oh7��<��uo�o����(D>� ��2`DΨloߩ (o^:���Y���ǂ;"ň��֞n���~�)  �R���b���]�"r�fG��uk�Pzzf5~R��PQx �%
�T=3��n@��^�)1��ip�(=Qx���iډ�(=�Չ�Y���� (����s�0��v  F�z���ȣ�- ��|̜^�ܔ (����&f�*"c�- ջ�%1���(�@}u��:�%w���9ӎ�n(TC�/(���QI�}��V�����8U���{V�j�BE����ȸT�jg�����ы�|�vJK��|h�& @qX{��n}H; ��1[��{�#o��[ �!�����J�R/j�  �ǼTj���"��- M�^턂e|��(�:����k}�Bk�)ݣ�����?ZS��P:�}���ΨMhwĊ�hs����3#t��*��N���g�X{RoS]�vG�8� ���7?���  ������Y�g�@���b�Q`�5���'�C  �K��-V��;  *f��	��x�㗞��@i�3��B�w8�v��H����<����^hF�t̞���봞�߮��4+
3v㉜��;���_�]Q�ھ!�d� 
d�&/��� �_R��V�Y"2���u,��yV̿'ҩ[�;  �[�0�{�v D�����/#Չx>5�����Y�5�-���vG���Di��r�����DEb�s�An�1�4�-l:P��PQXBFi����HM"nS5���O8!�9����� (�����iG  ��a�l���E$���w��~��T; �=aD�����ϵ[ �uMm���3
�?��#���6}������:��Y|������X����ײ��?G+����W;5��O*����k?�� }fq�G����� (�vO�[Ͷm� ��xl0b��v ��4���~#b�K  �S��y�{��l�n �y�Yi����(X��ƹ_����;�Ǌ����x�vG1D�m��x6'����3
�5�a֣<�L��"�m^����0+ե������������s��y�]t։���9������9 0qf����b@  ���W����@�c��j�2�3Mk�  ��Lv�\�-"f�v �lv~d7"�U��kg@���qʿ�6�%�;
U58*5}C����Y����L�z�yש��9�R��P�C�R�7������ۢ��pm%��2��g|�gf]�vG��#�2�{@; ব���%�[7k�  0���+�;�rƂ;\4,b�b:�۴C  ��D{����#"�w �̍�?	��M?��|����1�����0og4>�(]swvh'EǼ����g�����Oi7�ܝ��S�jns�vBQt̟~��m�vttϨ�T���6���} �D�����
  &�lڔ�b�w"f�vP�Xp�s�؋�0|V� �B%��~c�R� p��n�gr���c2�n�������O�x���z�b��=��(]�[���jg,��pM%3����k/j�;}�vG1����c���A����ي
3��1��Г�=���y��hw3 0!Fn����  �A���[D�W�
Xp�S���$��v�  �%_�;�; �E�lNf�vkgE����?���;0�R���;��������T��]�t�;�=�=�� q�} 7@Ddqt�.��uf�q�]Y�MP��=@���=�����}߫�����Ȗ��?U���s�'O�鼽}��~���nH�pT��f;.�I$T�莟���)�W�r�i�;0�"Ӌ�%c����Q�A^j���$*�w��Y���\�g�����f�׹�� 0������v  ���;�����!0�XpG�p�<폄�l� �d2��Eo��]�[  U�5�NH��ף��=�;0~�����QV�g�#�#�
Gmg L�q�	�	�G�99��݁���/�|kya��d��ܭ���� Sk]2��g�L���Kol�(,�ݑ�-���� H#����\nB�!�-  $S�)��#�[�;�LÂ;҄��K�i�v	  �f���G��$��n�t3��';JRS�E����R�{�_h�U���RQ�4���u.��ӧ���+�o�c�j�b_Ü���vG�T�d��oj]�k�Ek�Vt�.��vƞs�<MS�k�#Y*�� �����P0
� `,�#�/;����dܑ��0�K  ��in��$��$%l� @:���פ�^�I�x���~e�c/\깧�(/�vG�L;��/) �M�Pak�팤p�Q[q��mw`���X��������x	�iJK�팤p<F]%�8�=�i����E���J�$U2� GĹ��Ը�v  c�H	�/�Z���n2�H}F�B��3  k���r��7mw @���/b;!i�K&�<s��j�cg�eg�=8�|��d��ޫ�6w�d��0c�{��,ʟ���+]s�7^o�g�h�W�Q�ɒ�կ�.Y8Fz���=3����d��W|�v��9��qv�;�eb���43� ����?���
  ƚih�3�LҰ� ������g�p��  �S����
� �Nf�	�NH����V~�#%�;06�g�,�	��2�E�gH��4�NH���)_~���*lw`l4WNyj(7�5���vͅ�7kO��خH���⯭���\�T��IO�fg��H��{C��� S�|Ѩk^� �����6�ѝ�;�L����p��}Y泶#  OFJ�Gc��� 8L��}*hw�	�C��I<n����G.��3Kf��H��.:M�ab���N�fg��>a���Ͽ�qV�q�;��M_P@z��RQs�팤�x�'f3�]h�G/�xxV�B��4s/�& ���I�^e���l�  0��M�I��v�v,�#Uu%F��2�А�  ƛiii��K��n�t1c���"ӧ���Ko�݁��}ՅeuǕC�9�]*h�U~�/1�f�l�*2��5���6�H��/xWq��S������>���B��.�r@dZ��go\�I�H����ˏ�-�?�㞙��կ��� �4�ȹ9�ܼ�v  6�F��h����XpG*rr>���Pk;  [|��Fc�E� �.f����1j�Q��n���v���b⺾I�^��4kO��d�Y{#���2RÌ����USm� 9�s���M����H�Y.[2F���/,�g�;�(2��'\�Gk`�Ꞃ	ٶ;��� 8L?	D"�ێ  ���2�p�H����H=F?̎D�� �m�p�{F���0�u��4�a;#�'d�:&������p���k�]:�vG2y	���`;jBπ��lg$�Є���0{�����\���9e���H&�8����;�}C��s���:�=�]ɗg�.�ݑT�4��| ��1������  ���Hd������H5[}99_� @*0��M�~�H�- ��m����t��g��������{�s�w������H�������@��r�턤k-/���������M���ꓦY�vIrUԵ*�g�v2�[�������[w텧�W�u����M��� Hm�N"�A
�  ���et����XpG*p�|�80b; �Ta��۔0�4j� R݌}a���3���ܒ�W}�����۷t�ʟ	�]��"���b����#�t�-����7�����lw��m���Ig�>5�����b����
��ź�9�����������yi�eZ��`�u�Y�|�v  �9�hj�c� �T�Fo���v�6���4ftG �k; �T�k�u���v ���xB�w5��H��ף���V���[p��TϜ�bWQ~��d�����v2�'�М]�3�.�e�<��׫o�|���p唗��&mw$[�DS4��@��$���}34ˣМ�{���Y�[pd��:���lw$[����h�� Hm�#�_َ   ՘��~9�k%��$.�"ܑ*�ÿ� @���_���� Hu�\z����l_[yі՟:{���U����𬒙�;�¼��$�3 ��~PrlW$�Є���tR�37/˷݂ó�ƥ��g���9��I��/�μ�������پ���*����37_���ғlw���;�� ��F���f; �T�oj�2r��v�&,�#��d; �Tf���h�ZI}�[  �������vƘ�*�/��m�뮻�]>ŭ����,�<�v�X�$��Vo;�$�w�����vƘ�,�������O}���[L��v�X�$:~[��@�4�{@�u���@WQ~Awn����Է��|�������&���mu�3  �k����	�:m�  �ʼ���HZi�pn����񘏛��^�!  �����:ɹ�v ��/��0fZ�N�}z׮ն;���ȅwV�2�ӎ1�S�Ĭ=������jAU��1�R1e��={�����{�o߻p��8w��������������g�޵{������\z}͂i_Mx��hu���&v��  �(Gη}��F�  �:#9q�$u�n���wa�N����؎   ]�#�_G�� ����Y����mhf�YO~z�c�;�z/}����/��ݸ7�vʘY�{ː�*�ZT��c;c̄���ۯZa����G/�f���4�s��?����HOem*j1fB3�߽�����݁�[s��K�N������7�$��R�� @���/(���  �E092��� ܀w�c����}�v  �ƛ��.��v �,GZP���%K���������l����v-�y�H��ڥ�/#}�}��[~��ۯz�v�f�G.�r�I��	�];���4�����z�|�7�)��������͆k/9���������jiC������ ���8�1�kW�v  �$	�^���ȵ7c��bJxn0��öC  H7���5!�&� ��f�jTp�ݿn�S��'�iٟlw@�pͅݳp�#��]t�8��k��F����Ss�?���z�v�M8g���=2�p����|��f�(�g�vƘ:8��O~�O����]Z{B��`���S9� �f�ѿB��;  HG>��VI��;�t��2H]��]���*�  ���H�1���v ���ф�W���s�Y%W<��e�mwd���\���Sf�7��w�=�)�ݪ8�d��<	'#^��(:���,[i�#�m����>����lW����Uֵ�� ސ'��I0�g�^��?-��&��^{�5�g?6���e�e,������v  %9����lW  ��L}}�q<7Irl� ���7⑪�*oS�[�+  Hw�l���� ��-��q�)��]r�_>��M��:�k�%Ӭ���سp��F�>W��+I�6��,R�q�������Yr�_>���?��f��L��c}u��?	�柺a3)m��u��r�$�f�����~�������K?_{�{G�}���� �����s���C  Hg��Ƨ%������3H9Q������C  Hw���Grn�� �ycq��)3>��^|F����u7,+�ݒ)�|����.��Q�������Z�I�Hm���Nya��q�^t�ƕ����vK�Xu��ݻp�]1����'7w����v�F:�}�3�Ed��ŝ���o}��L���W�d��3��	/�Nn�Ҵ� �T�/g�B��l  ��7<�9I��;�tĂ;ƕ1�z �a�  ��E"+%�c� RU���+I��J��kV}�Sl���s˖�,���m���p�Um�c;8,�^�Sn��q�^ZP�^^p`��KO���f��	,����S�]��~�Q�t*_�@����^�lg���҂���f�ت�y�o��Wo��?��DVf��E�� xc}M�َ  �-Lgg���6�@:ʌ'�H/{KK��v  n��|�Ha� ����Q��|f��(Iݓ'N<8�b�37-���7����7���e�K%��l����фNy!sf~O��	���_Z}�埱��F�>t�'�i8�l���r������K    IDAT3���I8Z�A���������8Xp|�anٻm����H�*�J ��F����FJ� �M���r8�8R,�c��d�q�ys�v  ncjk{r�� �j��zM̐�%)���ԝ0��o���w�u��'Ɇk/�cω�w���n7�tښ��+�#2w�A�w���7#�>O�	�����{�eY�{�b�u�ܺ�䙻��m����� �ٻ5���vƸa揍��������eŶ[���u�l'  R���o��f~1  `���g9Ͷ;�tn��ѷ���6�  �U ����lw @*�M�ՙ���x�斾A��y��W�d�'��>���o�r��Sg�h07�Q�D�w7�8�i;8"����We��o�]�T;��O�veƜ6>�/�Xy����Y4��s�3j���RI��vpD<���<��vƸ���w�紭����l����g��]�ɥ��_8뷃���{�ӌ}a�60� ���%o$�]�  ��	�:�x8�8,�c<�g�o؎  ��|>�mw @*�VQYC��q�Y�_T;�t��ۮ���t���_���ʶ����x��q��u�:"MU�6����vƸ�<�02���gny��m����:��m���V�`�y�L���Q������T~�M�5�w�Y����Ь�M+n��;�[��s�]���wW��?q�҄'��f��| ����j�Q�!  �Y�)�#=n�H�u�V9�2�А�  ��<�$9�j� R�;Vn�'���1���温_z��D��x�"�=����7_���S�>�U�?�v�'m�V��_呾���.O±�1�������?�k�����?��>;�ٛ�xt�i���,Οh�ǆ_�VnϠ��-yv��F3�:?�zꎟ��G�pmӺ���j�'<�l�ŭW>���;��'��ᤗ�kB��� @�q�$��v  � !�vI��;�t��;Ƙ�;_$��
  2�/���lw @*��ޫy��ΰ���������O}�V��ٶ{R���]����S:��O�xԛ��Mr{u�ն3�c��ѧ���ΰ��lRi�����?�����on����S�Y3�,�|���k;Ǌ`��N���Gz��=����ΰ��lR遹UO�~����=�j�KoI���Uw��ƽ���T�+r��u"3 �z��x���#  �9�H���5�@:��'�/]�x�s�#  �$FJ8s���� HE���V����kb>�98��C�Y��goZ��=�d�'���O��у�O��?��r�{lz������"5�������5�J?��ս��+�l�'�l��e��ӿ|�~��Y?�-���/ ,Y�]�X�vp�NٰG��a���|^spn�ձ��ݫn\�C��������>R����?�)���cӒ�;�2� �����ik�Y  Ƒ7�����;�Tǂ;Ǝc�`Z[[lg  �i��G���;  eE�d�v����L������]�I�=6U-;�����f~�����i�{l��/�i��lg I�iɳ/�ΰ�bN�f~�7���:W�z�-�{lڲ���+>u�K{�O{��b�t�=�Uֶh�ް� )�Ѹ��4υ���ꓦ���_�X�[.��v�M�>to����'Tnj��<Kyf��L�m��=!� �cd��D�l� �Lc��<�6I	�-@*c�c�_S藶#  �T����$5�� �T4kwH����+I]S�
�+��#_���ٛ�������K/��������^w\��Q/�H�#1�c%��p��V�K��=%����ʟ��K׵����m���?z���_��3��W~3���gnSYӬ�yiCze�0����u���t�M�{����.=q�W=����{��-�f�N��e� ��`\��؎   S�C�Mr��@*���+%�1�1�c; �LeZZF�����<`� R�;WlS�'�Q�ﳝ��K'���N�̓�~���[z~y�)�����1�]ca��\֓7�?�UN9���:}�N�mg I����<m��f�$u��w�������Z{~������-������0�_k��
��� �n�ʗ�4�X#��|I�,�/�,���������t�z毽��s��s��gF�),����u{��� �c��9�H��  2�/�|9�p��4�v��XpG���
�h; �L�D��W�"�}�[  ����������Sl�����'����O]�&g$������������]Z0���G���kv�M�ݓ�J�5o{��`L��x�.=�B�))�g��ܞ�����c��W���~�_�i��c�����=�z��kv���.J=%����v0&��#:m�Nm�h�픔�[8!��p���;��qպ�X����cU����ӟ� W��_�-�x�ޢ�"f��G:u��Z� �TcT����c; �LgB��hy�W%�[�TĂ;����8�j;  �z��d%���> x��ԩqN�"Ӌl����	��y�������m��=���Ĭo\�퇛m�����z�e������~�.o�?әOm�;lp��_�S��r�g�NI9Cކ�e�ǩ�×�m��5�����~����n;\U7/��EK>�?)������1f���E�:��2C�5oG�斩qv�픔3��6�)?�8�K�|��	��z��q�O�n;\��:��i�pK_^�-����S�DǛ�Ƙ� �7�p�;M}=��  �"����+n��	-�?0��
�j ��;��o �B�ߓ�;mw c�s�����7lg���G���v�����	����j8�o;%�y	���'t<�Q֏���#)w�����_<��181���҂Fr�,������읍�3R�o�V�(5_|q�nU����3��`n��|�9l��<O"��-=�	݃Ogy͏���G��n�G�n��(��}07pug��sY����{�o����3R��@���c;�9��+����HyC���|�9�Ͷ���<��&��4M�X!g�������ݸ�pD#��������������h����3���W�̛g;�9�����=�3 �!�ѓ���;  �������Ȭ��6��XpG2m�E§i�v  �g֬����>I%�[��Ă;���y�Zu��igb��P^W���Pt�|�{����;ƻa�ˊf躡�����&�&���w$f�i�{��r;LV���n�sʴ�w��H;z��v�FW{��s~�Ǘǻa�ˊ��6���??waWQ�䄇���Č�a��O/��H,��ChV����]<>Bz���GV�u��[���B����`�e�����f1������M�3�&Xp`�H�cN���m�  �׊VT�+G��� R��v ���3��  �S[�-��o2��m� @*��?�y�����S�J_~nN_~�i�N���{�qS<�o�-8���U9�����_�"���z�S�&Ƣ�0r��f-f���.�;1��x�X:Z�=�z���lg ��@���V��g�NI+��������J:U�����M�	}Cmك#�ޑX��FJ'=��������Ч�M�4[�u���Y���N�.ߛ���?��!��)f>2�����R�݋g�NI+�y�����"I�$��=߼)�j����D7{b���r����'��r��`N�,�8zG��}�H���Ĝ�Ƽ�`b:�4�`����T�}p �~�r;  �)n���s���� U����0�c�px��  ��|M�_��+>-�$�- ���X�C-S'��p�픴5����$�Iz�_���߾�����マ�h�7��&�nGRV|t !3�qF}	o��x<�qr�ެIq�wb�����]�@V��3w�$z�U�G�S�qw��j�:Y�S�l�����g����:����7���G��F�INV,>�0����|o��7+/�g��pt��U
Gm� �;�4}����Gm(��R��3%�)I��έN�?:��y����X�ǛP��a�z��2&�g�H�?'x5�꿞�0� o����}�v  xc�P(<R^�?F�7�-@�`��O$F�d;  �9#�ƌ�t=k� R�/׹�n��׽Wр�v���|^+�u�ĉ)�{p�ikv�$�a;��չܤ�\�>E��M����%M��I���VYc�����xB�>����}\�'Y��5��^3�N]�Kem�3  )�|���wۮ   o��~+���:X�x�p��@s�n�  ����U���mw @����әOn��%�ؚ�7�Ulg V�u��ǫ��p�i�M:����3 �&v�ǫd�>�mZu�N~��v  5��
�f;  �5���od��v�*XpǱ��ţ|�
 �t�8���� �jZuD'V� ����ӻ��f;H	��t�&�^y]�:�	^� $���Y�<��v0f�� ������ٵ+j�  �=_$�kI[mw ��w#����b�  �@S����� He��ݥ��V�@���1���M��l� )����5�����E�:��/���f�nܫ�Zg�}�� ���D"�]  ��F�mw ��w5#E���v  82>�㮝mw @�2	Gg��%�u��N��$������賝��8:�������q���fMj���{�9t�_��k;Hf> ��cX�  ��"������Ƃ;��#�U
��   G�<������ He�CQ]��s���$Œg���@�� %�����+���8c�vM���� R�$��yA9öS��`� ފ���/~�v  8
�狒��M,��hU�"��ڎ   G������N� ��&v�?mRV<a;8&'mگ���� Rڄ����s��Fm� �dA������ʄ�������S�c�� ���c��ڎ   G���Xe��h���w��+F��/  i���wG�c� R]I�Cg=Y%�p@�ӌ�a-^��v��4u��'63�*k�u����3��0��Kg��%�3鉙 x[����/��   Go�q�,v4��Xp������`;  o"�GN�� Hu3��u��]�3�#V�Ю3gY83��u���3�#V��ُ�Ȳ.p*k���g��� �3 pb�D��lG  �c���t����q�<	�E#%lw  �ccZZ��� �N|�Z��k;8lE�]:��䍏�N����-ڰ�vp�
[{t�#��c�G����:cK�H�| ��1?�ni��]  ��hb�k�Flw 6���#���9��v  H_A��%�� �`ц=:i�~���*h��y?'_4f;H[�۫�_`�#��w�邇�S`���U5Z�</�"�1� �i8��ڎ   ɑ��\/�׶; Xp�1r��   ������o�� �tqں]:~[���M�u�낇6({(j;H{���҉Ulg ojb��.~`�r�m� io��=:�E^lB�b� ��`(�]  �'.�?�)��@,��H���DV؎   ��e��� H��g^��|��'��_?�A�~�q�r����r���u&v��7(��EG YN[�K�o����3 pF��p�  .�D��7�;��Ƃ;�q��l7  ��3�8r��v ��8z�S[����v
���>]r�z��l� ��H�^���ܑR��u������#�s��:��j�%���� �#c~�9�  �盒�|/2
�8Lf��)���
  06|��/��'+�p9���k�s{m� ��ҭK~�����H��ڡ�kw�.�|^hƎ#��f'3)�� 8B�Qg�;�#  ��F"�2���`<�������ߍ���   c��)�|� �Ԣ{X~�U%�]t�zeqh0�N�T�̇US��u�C�=8b;p��7U�+��T�0� G�9MMmG  ��3�8���#����ñ�
=i;  �-���sI-�;  ݜ��ZK�}Y&���Wem�.x�9��q�)@�8yS�޹b3�njm�.z����t�{�Vy	�)�0�| �Q��:	1 ��r"���g�/,��m9F�m�  �=S_?l��v ����kuޣ����NA������yt��1�ہ�v��:�����0�1>��׹�>'/4�n���:���y�㆙ 8*����v  2CB�oI�m|d��֌j���#�3  �����XR�� HGSk[u���+�7d;n�H�6�ѻ���i��Eu-�������Xze�g�Vy�j `M��V]�����7c� ���$<߶  �Gv$���<f�,��%�-#���   ��tv�:2?�� 骰�GK�]��V�B�e�:��p�^�) $��j�k4���v
\(k4��>��REA[�.�w�&7w�N�1� ��H�Zw��   ����?m7 �w��_���v  _������mw @�
��߯��}�)p�ܾ!]��u��'d;��������׌}a�)p�`ߐ.��f�f��$80��ؠ�{����a� ���߶  ���B/�h��`����7ed�oB!�� @�1m�͒s�� Hg�hL�<�I������8FemZz�jqb(��|Ѹ��؋Z�j�<�|�҆v]~�E:m� x�h\g?��޵b+3ǌ� H�|��F�  `�yF/���XpǛ����?�  �HHߑēZ 8�t�j]����خA:����C�R�#ͯ�х�W� C�Qp���k�|~���wܶz]����F�Q`� �đ�_�  �Y͡�$���%��&�_���n�  ���Hd��h�� p���v-�w���8}�/{(��}��  i���CK�Y��p�����pL���-yv�<��� ��$Ԯ���RI��v
�3 �<���<n�  �a$Gr~`�K,��8	�'�#  �]�|�v �EnϠ.��:-ڸ�ee����6]�gUY�d;�Q���%����;�a��m�5����<�i���@:
����7h�*������ �$���FmG   {|��}�Zlw c�w���ώD���   v�"�g$m�� n�I$�p�^]��u��=`;)ȓp�h�]��F��m� 8&���Mպ侵�|�!O"qh�?�Q��!�9 ��qͯ�ѥ�[���~�9HA�| ���e��  �2�82?�����zF|�  ����v �MQ�S��v�f�n�����ѧ��]����8���EQs�.�{���j�����٧K�[{h�s�?�S��u�ݫ5wG���f> `L8�����  ����W�&��Xp�k��ëlg  ���f�+>i I����ǫt��Wn��X�I$t�j]q�*Mn鶝`�Gb:��:��)�����<���o���w�єff>�F�h\�Y�Uݿ���33 0�	��mG  ��`ZZZ��!��X`���0?4GH   I�|���/mw �[U�6�_=��7Usjw��ҭ��]��kw*+���`�M�m�U�^yh�s�k�)l�ѥ��Ւg�����0���u�oW1�33 0���_�klw  �b��N Ƃ�v RJ�/���  �ZF��3��%e�n 7���Z�v���4iㅋ�3y��$�1_4�S7��	[jYx2�76��kw��:�����)�|����Z�~�l�a��3���6^|�����N�c� �G�'�  @j�G"[���$-��$��;�ݦ�e�v  H-�H�1V^�#-�� nV�Е�yV�'Oז3h8�o;	��H3��u�����]���H����*U�<M[�3_����$$�_g�����a�����K��v53�͘� ��S�DVڎ   )��rXp�����W9	��m7  ��d<�N�a� Ƙ'��m���7�m�>^{�T�㱝�$��ԭ%���8�a;@��$�|���ܥ%��P	3�+�6��ڹ�8�<}63�%�� ��d���H	�   ���y0�8�#��v�,,��Gk��lg  �Ԕ
=�(�Z'93m� @&G���횷�^/�s�"Ӌm'�(���u�5kO��خ���~�t��
�,�������u�5gw3�
Ǵx�N��ՠ��>Q�Y��t�� X0���v  HM&�VT�#Gw�n��w�Z#�    IDATH����v  H]FJ����7m� @&)h�ՅnTK�dm=�5M+���Ô38��/Uk��e�9X��+h��?�֊�������Oك#Z�R��o��7>j;@��ޫ���Z����ǩqv��$&f> ���MKK��  ����S��g$�-@2��Ij��Q���  �¼���bY޻$�-� @�)	w�6�e�dm9s��+'�N��j���YxpԊ����C3���T9�v�ī3K��1f>�#W��y�<h濇ZS3 `�q8�  ���Hd_��b��sl� ���;���mv���   �ʹ����*s�>`� 2UI�C߿N��J��j���c�������r����� .P��E��WhV�v�1����҂�5:n[�|Qf>�cW:�Bkxf�v�1G��Ŷ���`ߐ�o����j��  ���"���#  @�sd~e��W`��3�[�	   =�,�'�� �U�6���Y%��k��ͯP�㱝��
[{�����Q��c;�M�m���Vu�k�isU7��0kCA[�N�Z�9;�O���Bu-��kQgq��.��'NӨ��|�� �Tb���v  H~���X4�%��vp�Xp����=�#  @z�
��N�W4J��� �&�t�'�t��=ڽx��O��h�g;��L�����������!
[{t֓UZ�a�v�6[�'N�H63��QE]��WPE}�� ���G�Z�U�<���u���5���z�| @��{}��lG  ��`�뇣�H��vp�Xp�t����  �>�4:"�wF拶[  3�g@g�ڮ�kw�qN��-��ȴb�~�*�?�9�uܶ:M��� C����U;t��]��1��?���u��u����`GnߐN_�S�����C�| @*3�rs�`��  �F��ȓ`�i���6�x�  ҋc�o��/�ǩ �r�F��/����<Q�O������Ͷ����F�ZӬy��UQ�*�8�� @�kg~o��?e�j�O������I�2�_>���-2	f>����3����^P��	\�-f>  ]$8�  !s�K���N���3��#����v  H/����hy�s��m� ���;�t��:m�.�V���
�_���a0	G�M���/�Y��=�� o)��_��٥�kw�:�돛ʲ�ax���R����$ xKy]�Z�v�N]������+4�u��b� �P��0�	5�lw  �4c��q}�vp,Xp�`�q��   ҕ�ɰ� i�8�JB*	u���;�4�H��U(4��%��㍏���]��G4}D�a�������g�ޡȴ���Rr�﫼�Q�6th����U7�"���3��r�ꏛ���%��c;/e�:�Ú�?�� ���̮]��  8b�x��X���Ď0�?�ʑ�|��j�   =����e��X[2 �F<��*�ZTQ�"I�T�25�.Us�%<˅�kb����[U~�Uu-�E㶓  iL�QE}�*�[%1�_;�[��l'@Ҙ���m*?�&�3�e��f1� HK����N   �ɴ������42�n���8��H��;  @z2���������m�  ����Aͯ����E�^�L+RKE�Z�NV{i��a�;�T�PI�S��m��=h;	 ��kf~����S�:u�Z*
�|��f~g��Ý7�l'��������\9Y���2�P����y]�*w���� p�_sc��  ���1���H[,�g,���  @zKs�qĂ; ��?W�&Uh�$�fy�^Zphٽd�����W��6'������G�[{U�PQ�Sك#��  %�Gb��iRe��f~Gi�Z+
�^:I]S��[8!mf~p`X�=*l�Qq�SE�N�0�@���TYӬʚfIR��Q{�$�VLV{Y��������[��.�;��  Wrd�3�c�  �/���c���I
�n��逿�7} ����|�Ec=��m�  �/k4��p�J���٨ף��y�*�WW�D�LP~���s��ƽѓH(�wH{4�{P�*h�UA[������ �*k4��p���~�gy�=%O]Ey��&�??�����3�Qn�&�jB��&u����W���| 8�DBőNG:_��Wg�+s�� ��u��\E���(����:�gP��{���^^Z dG	-  �Ĵ��E�+��A�-��`�=9��n   ����G�+�$�z�- ��OhrK�&�t����??�����r�5���H�_#9��'�W�E~IҨϣѬ�W���q�����UV<.4��PT�CQe�(0U`(�ʂ㐂�C2	����5��3$ۯ�I����`0[��@�g�(������Af> ������A����9Es��>4��n�K�����qe�G反*04���7��=�
�1� �ΩʎD�ٮ   �ϑs��a�i��4����v  p�x�wL�w �+�QMi~�R �]�Q����l� 0��Q��o��  Ɔ1��� @R������.I�[�#��q�5;��  �������v�         .����#  �;�F$��vp4Xp�0���  �=���c�;         \�ŜH��v  p;�HS,�g�D"��  �.�        +#�g.   ��rr��L���H���Q��@S��  �]�JJ���e�         ��feqh!  H*s����'lw G����/  f���<i�         �m�nl��  ��q��(����  ���:        �(��  Ɗ�$�K��	�3�Q�?~�v  p'���        ��h�m7   w2�Ƞ1z�vp$Xp���   �eB�!#��v        @�1�47첝  �ˑ�b�8,�g#=n�  ����	�         i��3  0�|��OHJ�� ���z'MZo�  ��ϟ��$�v        @:1�á�  `L���6I/�� ���y�����  ��<�$�-�;         ҇����]  ��=a�8\,�g ǈ7} ��p�u        ����B  0^��@:a����x�)�   3���        �ar8I  �8�M�A���`���^2--��#  @f�55n��b�         8�X�C ��1z�vp8Xpw9��3�  @�0�#9���         H�Mk+ �q�H+m7 ��w���Â;  _�p�        �6�L  �/V�JI��;��Â��xs�lG  ���xVHrlw         �2�,� �qe�d��v�vXpw1GZc��  2KnccD2{lw         ��a���v  �<NB+l7 o�w3��  ���        �7��D"��#  @��[�4����9�g��  ��<��/     ���ޝG]v�u����95�2��*U�y��"��!L����� A$�p	��(.Q�Ah�����A�!	AW_n�Ƶ����W��4��#d"&��U�<�9�w�(��J�s�{��z�O��Z�:ٻ�g� �}(aX ��r�E�]�p0��u�����rv 0��KK��     �6���� ��T�����?gw����T��|��� �|*��vW��Bv     @ݵ��|� ����p0�=U��Iv 0�j�     ���?���^��  �X��t�j�=U��g7  �F��/     �=j1( R��=�/"b_v��~�}�7|); �o��?��&�     �UJ5p R�k�Y��%�{�(Z�� �d�n�����     �"�G����� �Z���e��G�� Z��     �?����k_۟� 0�5���{�F��  5�ϲ      ڢl: �v--�EDL�;������u뾘 Q��?�n      h�Z��n  ��(��枈�Rv�����E?e ���[��6"n��      h����; �%\H+��M�>l �V)��      �ߗ[ou0 �~]��2p�6 @�Tw     �2 �]j�8T�V2p�:,� �v�9+      � m��替wdw�=���?l���k�#  �n���_#���      �TJ��� ��+5"�[vܓ�{��(W�� �5�7��'"���     �h:��bv �=�(_�n�{2p�Ƈ �V�S     �9V�g�馽�  �����1p�2 @+�(N$     �� �N���2p�Z�L �V��     �_Ŧ h�7��Ո�+�����?��p��dG  ܛQ��n      Hd� �R�h"⯲;�����/��! �:妛�Y"n��      �0*��  �ͯ��.��A h�&��
     0��+7�p{v �}���	pw�}Qꗲ  ��_     �N��?�  ��Ʀ�V1p�2-_�n  8�R��     `�� ��F7��*�=1���! �ݚ��!     `�hl: �V+�^{g��)����{?�Zn���� ��YW�_��&�     `�w ��j��i�>��A h�r�M{#��     ���֯��� ��UlQi�>(�[3 @'T/�     ���r�wfG  ܯ��t���x� ��a     �5�M �	�46���{�:�jv ��(�^��      0+%�o�  �he�M�a���Q�P :�ܷ      s�ֿ�N  8嶯�{�; ���&�l�.; �PL���     ���  �rmv D���ߗ��^Ɏ  8���#b)�     `��� �Q���h���>L �)MD�}v     �4�7m� ����h	��+>L ����=     `.\W���/� �Q��� ����j�6; �p��     �y`� tJ8t�v0p����  ��D\��      06 @�L�Z����J��  Gc�     ́j� t̆n������n��a �R�c.     �%�w" @��k�Y��[�;���ۖ��[oˎ  8�C'�     �W�C �*a�A:�.+qC�h�3  �׿~KD,gg      ����� ��Whh�n�! t΁�ʍ�      ki����  �����g��e�z :��     �c����ۿ�] p�J�m*��;�ܜ]  pd��      }V} tR��t�����J�[�  ���     �ϊ�B �N����0p�Z< �TJ�0     �V�� ���ǐ����J�C ���     ���B ���/�l:Hg��a�L}�  �TK�u    ��*��t  �t��n��&;��f��a+áa �I��w     ��ju�; �M%b����|3p﮺i˖۲#  ��t�E=     ��j8� ��^�T�U����^ɮ  8�ܞ�      �V5| t�]��;�~+�  ��}�kߎ�&;     `-4��#� �H���eHe��]>< ��*�����      XM�8� �Zý�ܻ���  ��xa     襍���u  �5p3��;���A ��~     �i�~��� �#UmTIf��Q�  �>o�     }tg���  G�TUr�wV�3�  �h��     �*6 @�l:�e��Q�?e tZm��     ��Wm: �N�a�A.��b_v �Qڛ      �| tڰ�3�2p��a �>�3     @� �4U��wU�� �6C     @Ո}�  Gæ�l�]5�0 t��?�     =40 :�{d3p�(o�  ]�~     �#߁  ]WKq?C*����  :��     �K� :m�`�~�T�Uk]�n  8*��?;     `ՕX�N  8*զ�\�]5-�� ��Q�2�n      Xu5l: �n��.�R�wՠ�� t[q?     �O��  �q��He��U�� �q�/�      =T�M �m�6��!��{GUw ���3     @5�; �ۮ����ܻj:�� tZ-��     �Z t��R�w�`�� ��`0�n      Xm�Rm: �N+5"��旁{w��  ��Q��     �^� �^�#��{w��  ��Q��E    �^� ��� ��j @�M�f��      �ښZl: �N�a�1&��|]5z :�ԁ�     �j� �u�gHe��Q�� �u�3     @� ��۵���ܻ�� �ZG�	      ��� ����� ��{W5C @�U�3     @��ph! �q++�gHe��UC'� �V�q     �6 @�w�M��;�Dl�n  8*Mq?     �O�  ���Z��n`��w�4bSv �ѩ�g     �>� �i�j�A.��*� ��s?     ���@ ��s?C6���� @�5�g     �j� ��+6$3p�(o�  ]�~     �R� �n+��t�����|x  ]�~     �#߁  ���B��wT�� ��sz	     �Oa @�M�ϐl���)����  p4J�j����r��QO=5;��3h�y�a��� ̷�:�- ��0� �� ��J�ǇM�ܻ��d'  ���se����ח �r�9��/���@�r���  �| tZ)�Z�+�g->������ �y'e      ��j8� 讦�Q%��{Go� ��~     �;v�� p�J)6�2p�b t��    �^ڿ�d� tW��eHe��Q�� �U܇��     ��á] �Y�:��\�U�� �;N��     @O�R�: ��*6�$3*���]�#  ��Ғ7}    ��j�rrv �Qp/C*�۷w�� �#1N�f7      ��R�Ӳ  ��{R�wب}�  ��DxQ     �� ���箋���;�o�6x� �R��     ��J�� :i�-�l�����|3p��� �Qe�w     ��J�� :i�46�3p��� ����x     z��_� ��T�T��wX��/ �Q%��      �� ���:��t�]Vckv ����     @��t  �T�M�ܻm{v  ��);�      �бuǎ��#  W��M�ܻ�� �z�t��     ����Ʈ ����t��6��� �ñw����>�     `-k5p :�:|�0p�Ѿ�ŭ�  �c]�x�     ��8 �&���w��۾ @�x�     �� ���Ǜ"��0p�8C @���     ́b� t̒�Z��������  p8��     �	��  �2t�BK�w\��3� �p��n      Xk�w" @��Rve7@��{�0 :��     �@�X���� �C�=Z����- tG=p����     �(����� �CU���
�Ww�ݻ�gW  ��۶m���      31�:� �Z�{Z�����Kw��T �F��!     `n"|7 tB�(Qï��
�=0*�� �	��     ����<(� �P�[XX��M�a��M�n  8��G\     `�� ��9l�1p�A���  ph�ò      f�F�n ��4�[h�>�� �n(��      f�Dl���'gw  ܿ�-*�a���b @���xSD���      ��IӜ��  p���;�a��'��gl͎  8��:|X��     �L�NC :�a˴��QOL֯�` �mи_     ���i� @�Յ�S"bKv�����x Z����7    ��S��
 �ۤ�_�U���ԇg'  \�0     ̝a� �Z46���{<*;  �`��n      ����n>ckv �}��n    IDAT���V1p�g�s�]�� po�֭�k�8�      �d4ydv �A��*���q��[� po&��!     `�9 h�1�(�3p�2h< -e�     ̱�TT ���ϊ���pw�� Vգ"�c�  �T�JQ����~��� �����Ell��~��|+ zop�F����I�����gg p�?+���3�5��v*զ��i��r�|�  m�>��7��߉���gg p?O{jk����c��7gg ���y?�ځ{|���[ �q屏�b���Au��˵�ޙ �]�xd���n�� VQ�GU�� -SO=���ؕ�     ��L�.?2; �^8���1����m{Hv ��M6lx\��     �ݠy|v ��Ոa�xLvܓ�QϔR���  p�O      J1p Zee<>'"���{2p��a h��O     ����8/� �8T��2p�b@ �K�x\v     @��m�x�=� ��9���2p���~. h��۷?("N��      h�a)Fd @�8��V2p��d���� ���2��      �I5p ڡ�q�"����7�}4��  ""J�/     �?)Q�/�  "b:�|_D���7�=Ԕ��� �ܗ      ��c�x�); `�46���{�O��� `��;N���gw      �ȺI)~ HW���Z��t�ʶ�̎  ���d���&     �wi�1 ��;�(snv����*? �x�     �{�Z�?� �o�R΋���p_���۾ @��G      ���gl��  �_����{�F�W��� @��y�qQ�Q�      -�q����� `~�Z�i5��:ye<~dv 0��6<)"F�      -���  `>���c���;�`�{�D�`v 0��Z���      �V5��R ��iyRDl�1p�1C @�Z���      �bO�'�|Bv 0jilKi=�~{b]\<&; �/{"�Y�      -6Zڸ���# ��d�N�����I�<1; �/�Z�%�     ���e ���-[N����;����\C �l�     pP�w* �L-�;��N0p��i� ���%�<%�     ��o<ޑ ̏-����� �|XY\|lD���     ��R���  ̇1�O��Ca��e�ĳ�# ��P�w      �Z��� `>L-�#��@-� ��(Q�w      ���:o��  ��qh!b�>J�S< k��oGģ�;      :䘥��dG  �W�L�����c��<9">� �׺I=?J���^:�\tQ����kj��|&�-�d�    0'���Gv �_{���qNv*�9�4q~� k������G'��O~2�#�]2?~��1������%    ́Z��5��%�W- ���r~T���� f��8��' `m���c���X}'��O}ʸ}�N9%FW^�q��.   `��m+۶=:� �z��d��9Q#V�� ���4~("��� �N��'>�~)0�������x��    ��:</� 觺s牥8��n1p�#��� �~*�q���N8!F����۳sL�~��^2    `͕��n  �iy��#bCv�9R�>�F�� �_�]"ʳ�; z㤓b��+������c���Eپ=�   �~;si��� @�J8���1p�/g��Ǐʎ  �e�o�S#����^8��]qy�ݾ�j�SN��G?q�q�%    ��`0q�; ���x��F}Zv.�9SK�& ����M_�Uq�)��{Xv	��<��1�ЯD?�   �ڨa� ���RΏ�M�p���L��m_ `��s�]�:���N=�������K8��ӟ�K.��    ����??$; ���B:��}�����xNv ��o���89���N=5F�_��.��-Q�{Bv    =5,��� �����vlD<3�����<j�e'  ���� :���e��(F��Q�n�.   ��j��� �~X�{nD��G��}�(/��� �R=㌍Q�s�; :k��]q�q{m����pĺu�%    ��Y��̎  z�8���2r�O�'۶�/� @�-//?'�����I[����WFyș�%�r�1���dg    �C�c4 ���œK�S�;�H�ϩZ� ��2� Gd��]��(�ve�p��xE����    z�D}a�� ��J�?�;�H��_�ݻ}x G���qR������ٲ9FW\�L'��B)1���<�A�%    ���ɶ�O̎  :�V��i����;�xzv �M+�悈ؐ��%e۶��Dy���SXM��_�qcv	    =R�E� @7��wD/��i�slX�K� ���/�. �2���WF9���@9�^ziv    }R��:o��  �gt`jL��<�j�g׭[7gw  ݲa�̈8/��+�������G~$;   ��8q�~8; �Qj��y��m�J�(; �R��"�dw tAYX80n?���f`���Dy�ò3    �R��. px&����e�>�J�߲ ���A���; ��,,��J����qc?|Y���g�    �O�ڎ�� @wԩ��w�^�� t�ta�5b1���ʎ1��UQNߑ���;c���dg    �e8��8; 膺y�qQ�y��܉��7v �CR�xiv@ە��^��(���W��>7_��   @�����  �`eݺ#��Xn���zq�7eW  �V�n�\K<;������1���Qv8�}�/�4����   @��N��dW  P�+�`��񀕈�# �v���+"bCv@[�>0��(۷g��6��×E|v	    ���� @�-/,<"J<.�V��;���� ��jĠ�rIv@[�>����۶e��"�3b��_��    ��j�g�]\\��  Z�'�`5��h��[޶��������) @�L�M}`v@��;cx�Q�n�N���~v��������g� ����@���Y�?���G"��Y�?  �cF���� �}ꩧ�R��������*"^�� �Om�_{�e׮]yEĖ-����Gs�g����E�f��o��s8�yO�θO�K/��߿��_�NX5��?=/~��������  ��&ʫ�羻\}�Jv �.+�׿8"����d��ݔ��?[���� �=����k�3�; ڦ<��1�⊈-�g{���h~�7b����o�l��R�U���G?�O�N�w6��×�䇞q�]�5    tP�ض��o<+"�0� h�rIv��Av ��ieҬݱK @'kyUD�; ڤ�y�wNn��^sML����������n߾���Q��O�K�Sٹ3��~wv    V��&� h��������Xm��C}]�� ���k׆R� wS�q��َۛ�~6&�|Vԯ|e�����c�җE�?�]r�</Ͽ ;   �������s�# �)��	����]K���� @;������-� mQ��}��SO��u���w1������u;gi)&/}i4�G�%�i��wGٹ3;   ��*M��� ��m�vz���X�|�A��g7  -Q�$��r�Y1���[fxr��JL��Ƙ���M3��v��JL_��h>���{w�1��_�X�.�   �N*?VO;��D @c���fw�Z0p��<yya�� @����i�g."�<�a1���SN��E���_�W��}���W���'��sΉ�O�tv    ݴa2]� 䪧�z|�xyv�w�]-?��  �jJ����6(�w���OE�|��.z�1y���ٟ��}���K^����K�����Dlq�    G��O�ݻ�gg  yV�m|yD���k����P_�'� `~-��-5����-e�~�m1���Q����]��&��������f�|���c���fW    �A5b�|��?�� ��(�u���ܹ/�#����*1���(� ��9����+"N:if׬7���]�+_��5{o:���*��~6��{^�N��    ��J�o��������pAD<(�֒�;���xmݹ�OX ��ٻ��Q/�� �TqN�>�Ɉg�HTo�1�ϻ ����sc2��k^Ϳ���%���c��WeW    �M�L�->=; ��R˛�`��s0'N��^� �֨�o���� Y��g�����=n�-�/�(������f2��k_ͧ��.�.�K.�ؼ9;   ��Q6� ���������Xk�\�7�ݻ� `N|��[��̭r�wNn�fw��o�ɅF���]s^M�1}�������iS_��
    ����,,��� �N��7悁;U#V���� `6&KK���Y��я����v�~�1y���Ͽ��5��t�7�t�F�X��8;   �.��g� ��X^XxdD<9�f���CP~��� �W��5^����<�11���#�?~vݻ7&]�K_��59`:�����g��~}^���
    :�Fy��x��� `�o�����`�̡x����� ��Z��+#���Y+�yL�~�c��7ML_��Q����]���4Nr����.����.�r���    �gPJyKv ����m;�F�q27�9$�ַ9� ���q��R��%0�c����l��1}�ۢ���q���^�ӟ��h>��쒈��)�    �/�??$; X;�1l8�#��s���充�eW  kceyrI�X�� �����w�L����oF��>2�kr���~1�����\pA��۳3    �� ��eG  kc���#�fw�,�s�J�ow�; �OݵkC�����Y*�=!F�Xı�������b��w����Zc�����#�/�F1x�s    誋�/,�� ��AӼ="��0K����{y��s�+ �յ�w�%5b1�`Vʣ�����M�fz���/���~*�ifz]Q�1�ŷF�ۿ��1x�"F��    :i8��w �����3w�9,�Էֈ�� �������� ������|���VL_񊈽{g{]O�1}�ۢ����kز%���w}    ����۷?(; X=�Z�NGb��s������� `u����*���������egp��oG4�]�v��eKڵ   �Ѡiޖ �����C���; ��;���xW�F t^=�c#�[�; ����'����38L�w�+�_��9s�   @�ոhya�� ��F�'l5�S��3W��dG  Gg2�!"N�� ��n��;.ͮ�M���h>���    p8��wdG  Ggy����(���,���uq�� ���;N�5ޘ��w���7bϞ����}��9;    Y�������; ��P��FD�΀,����R뫳; �#�<i~."N�� �z��\uUv�`�����|pvܿ4�k   �K���f7  Gfe��'E�S�; ��;G��[��'��� �z���J��dw �]�ꪈ�$;�U�|��1�����u���M4����_   ��+OZ���] �z��v�k��S�7�3� ��YYY�4"6ew �]��W�Xeͯ�JL����������/�سg�   �ܨQ�Wm� �S���ew@67��R�M���� ��YZ\<'��,�`ԯ�mvk��Я����^�?��;c򢋢~�����   �W�ZYXxqv ph����K��dw@�s������ �5���fg ��t�ￖ]�i~������Z�?pϞ�������3    "J����vڱ� ���|�[���]����/o���� ��&���,Q���0�7F,/gg����.����Q���A��1���~�    wS#&���; ���;v�Tk�%������0�A�� �ՈaS���; �ƭ�d0�o�VL���#��o��Ϗ�W��a    p7�ƛ��o��  ���d���89������Q������:; �w+�^5��0/ꭷe'0#�o�NL�g#n����Gw�ͧ>��?#�W��vq    p�q+++�fG  �n���#ʏgw@����A�Sw��\�暥� �_ԓO>a�Է�(�) ��p��t^��OD��ODl�e불㎋ش)�ƍQ��1�F|��K����={��   �;���[���������% �w+M�`D���61pg5������xov �/V6n|W��5�`��a�>�n��N﯉)    p�4�\#�X�� ���x��q~v�� ;�~�Qq�x�#� 8`i����� ����    �{���m�eG  �ݻ��(���md��j�4����%J��Z�+�����;    �>��ԝ;O��  "&��#���h#w�@}����dW ��[�_%~ �`.�    �t����_Ȏ �y�waa�����h+w�Dm�j�(� �Uݼ��A��gw ̫����	     ��D}�Ҷmgew �<��@D��me��Z9{����� �W+�ֿ�F,fw ̭}��     �˺R�e5�d� �<Z��fw@���fj�K��v��; `�,-.�?��0��   �V+OZYXxIv ̛�k׆�C��vM���׳# `�ԈAi�#b]v�\ۿ?�     ��j|�nݺ9; ���}o���dw@����J�Zڶ��� �+��OD�y� so2�.     �?����ˎ �y�<~H����w�^��Vw�<1; ��n>ckDygv ���w�Qr�u��?�[��YYH�]ϭ�4!(A$�(*�Q#��
q�N��0�Gp �2�+�����QA	*"!�&.$]�V���e��]O-��9z8F�9�J�s����       �9���t��  t:�,�}NR_��0pǘ3����0� `�����$M�� �4n\�       �����0��	 ��+��%��h��$�Ƽ2�w�
  :�H����;  �0p      �>��eْ�  t���O����h�ĭ8ӫ��C  �4��;��,v �L��        6��N��� �N����J��h'��LO�
} v  �&�N3�@� �Cl���       `K�����9}�C  �$Y%=��/����h*��=a��  t�z��b�^� �O�L�]        [�I����Ď  �S����>�hG��l������q�C  hw>m��E៏� xSy�       ��c��d�ʼ�  t�z��9I3bw 툁;b�%˲�bG  ���q>!i0v �_�dnp      Жʲ�L�;�7v  �¡�zy��]1pG&{g>P�'v  ��K$?.v �Qp�;      ����lݺ%�#  hW�}6v���#��}ѧO�; �v�3L�,v ��Y���	       ������2�w�  ڍKV.��$M���3��w�{{�;v  ��� �?v �1�i�       �����Ņ  l�<T�d�cw 펁;"��k���cW  �.�J���� xlB�       �F�c��wj�
  �E-�]$_������f��  �Ս�$s�~ �`��I\l      �͹��t~�  Z�ϛ�cҗ%M��t�h�Y�t�K; �V�R9i_��]� �汔[�      ���u�ϚU�� @+�V���dO��t
�h	�:0�T��  �Ue!�,�ٱ;  ��v�)v       ��yV���R�  ZQ^�>�d��t�h�d!�; �V��Љ�;  [h�α       `t��_U�_ �?�E����Q����O�����'� �U�A �Wr�aRoo�       YM��    IDAT.?9OS�8 �&.Y=)}��J���0pG�����}2v  ��B ��lpPɫ_;       FK�]�����!  ��z��ݥ�cw ���;Z�1Y%=2v  ��Cx� �����Vi/�      �1��z��#  �-|��>��T�њL˲4�#v  ��i�l��A ��;���Ǯ       ����,TŎ   ����GRo��S1pG�/�E>m���C  h6��)�Œzb�  �]�7�v�=v       �"?5a��  4�KI�h�/���[�N���l�|��3cG  �L.%y�|�Ki� �()�U���R�-      �=�]�3b�  �L�4}����t:�hu��
 �U�>$�� ����7Iy��3m�]Uzm       t��yR��K��-  4C����kI��0pG��ei���  ��z��7��� ���'׫���K�zS�M��f�Svo�       0�����bG  0�֧i�]����`��v���___���C  +#i����eI� �A��q�;%��Z.����H�&5�L       c.[R�T_� ������ʅ�*if��[0pG[0�@���}Μ��-  �6�>}R��5ISb� @7).�X�����gڎ;�t�i��<      ��af�������!  ��<�Z�g�� �	w��g��7,� �hr��=}gK�o�@��_T�O4���/Tr�	M=       ��$K_��a.t t�,T�,�kbw ݆�;���Y��.v  �%�%nzE� �f�S?�bYs��-��=�g=��g      �{B�e�T� �h�C�K�Scw ݈�;ڏ��@u��  l��1���  H���⢋�w`����>'͜ټ3      `���Y%=)v  �jCC.�����-@7b��v��_�a``8v  [�V����_�@kpW��w�����9s��_:W�8�yg      �3�{k!� ���3flW�}C�U�0�B��YJʗ����!  l)�1<`�_*iR� �?h4�x�"����iG�n�����K�r��      �1f&;'O�g� `K���{�Γ���-@7c��6�fYv�K,A  mÇ���=��%͊� xy����oڑ�߾*-�H��      �&�o��͎ ���C�Q��$v�������y�� ��p��,���g�n <�T?���~մ#��W�4�<       h��I���gϞ; �͑�p��w�� ���e!�1v  �'����� ���׿���#��}ӎ,��D%�ڴ�       `�����ȅ.�c�  �X���ޒ}.v����C�i�4=(v  �&Kӣ���� �-p��jz�|Ŋ�g���>��/m�y       �&{Q���� ����u+�!�7v����S��Ey�>;v  �,O���:C��n l_�Z���9�J*�~����9�      @S���P]� ����`��q����[ <��;:�w}k$M�; �ժ����5�/ �-���?\Z��9��*��L�߾�9       ��������  <ȧM۾�Q\.iV� ���fz"}�g�� ����a��&�n l��oT?�hi����ӣ�gȞ���       c��:3�WX ��y�z�q�/��G� ���;:�kv^._���c�  ���������n ���Տ9V�՚s���*�w����4�<       {=.�$KSƄ �h\�|՚�$��#c��eO�J���y�zb�  ����O�]ߒ�K� ���k�U��o����8~��眣��6�<       {��u����c�  �S���tT� ���;:�I�׬�ХR� @��y�z�r�bIω� �������.Es��Q��W�`As�      �1�R(��W��Y��- ��W������; <6��h�zY�O��  t�J��5_6��@�+��55޿�y�J*}�T%�Ӽ3      `l���Wx�:-v �;di�:7}(v��������Jzr� @gs��>'���- ��(��E5>���X*����U:��R�ܼs      `�����m�1c��) ��V�T_&קcw �<|G]�L��C�sϪUM\�  �I�KM~B� @s��.�~��׽�ig&�+{�S�xӛ�w�ٴs��٬!�3�;�c���c���Ųu��􌮱~���/�]    ��yO�7|Μ���j�c  �'� �_ ����a����S�J�Ͻ��>#v ���i�>w��� �8'H����WѴ3m�=U��﫸���~.5M;��5�*��=�=v	�QfO{�J�}"v6S�%�:��Y��   @;�����t�I��1 �ΑW���¿!�/v������d���R#w �h���m��`� @D�j��]�v���%�;��Oɱ�J�ۼ3��;NTqᅱ+      ��⮗���B_��0F� �ѐ�鳽�oI����Ib Mf2�\�R}u� @��Bu�\�� ��B�Eo�_}u�����O�>=v      �u���<��T�� hoY{��rI�b� �r�э3?���C  �+�5��� �B�u��V~�u�K���LQiɒ�      @�zeҳ�] `+ei��dWJ�����At��ɾ\���! �����1��!�b�  Z�Ȉ��'����.�6J^������      t�c�P=��~ `ժ���JҴ�- �wt��ɾT�T�=v �}d!'���Q �G�׿���W�o�5v	�Q��Ə��      t)?.���e� �\Y�>�
�Z��[ l�Y�v�f~q�R}u� @��*�$;S| x<���.���%�64����;      �^���z���9 ���B�S��%͈�`��� ����,M�� h]Y��N����O ����ܣ����'v
�A�p���O��      t1?.��.�c�  ZSV|�dW��ہ��@ب$��Y�� ��<����x�! `��w�q���ڵ�S���e�N9E*�b�       ��<����y=�C  �%�2�ZҴ�- FO6I$;3��=��W.� hy���]�� h_��[U?�0�/�X�~��9�
��S�y��sΉ�  �m`�>_6n\�`��-���yg�  ��+�k֔|��#l��,v  �<M�uץ�O��`t1p.��sy�{V��h� @<.Y�K��?b�  ڟ/_��q�Q��/Kj�R�]��W\!_�*v
   �R��Se�3�1�X�D~�bg  0����|����/����[� @<�4�_�.�4>v�ї� Z���ZK]��1 ��s�����ĸ 0z���T?�5R��N�֘4I�3�I=�      �l���{����C  q�B����51n:w�Q�lq^I?��:���s���!�@�b�  :���j��R�;[���T�����       L������`�� h�,�7��˒���`w��bz]��}�<�a ]�C���]�MI��� �\���V��wJ�S���W2~�       ��=�����N�K  ͑��b�>#��@��9���֬����O� ;^�N�eW��E�[  ����"5N:)v�R�?.�y��       �;��5�����K  cǥ$�t�/���9���\��5>sf� ���000�~����n t��/���bg`kL����?/M��      �z.U-i�8��� 0�|Μ�<��K�(v��a�l6{Z^�n$�'�. ��Z��[9)�X�.�[  ݧq�)*�<3v����D�>�I�,v
       i�'~E-��c�  F�M�ׯ�B�a�[ 4w`�������!<7v	 `��!�o�~�R� н��^;[!9�EJ^���       6�5���P=)v `ۭ�VӼ޸F��c� h>�����pH� ������}[��c�  �����X���.�V(��ݲ���c      �E�ɗdi�	g m+K�=z
����c� ��/䀭3!�}-�űC  [�%���Ir�-�'v  ��FC�7�I~�b�`K�J*�3����%       �zkVI/���'�N l��2�B��q)�nw`�\�4�L�7��$ ��3�/��&_"�b�  �0y��������%�RS��t֙���K       lb��}?��S @��*Յn�e�&�nW9v ����|��a^`wܱ.v ��y����.�sc�  �6lP���U��bٓ��[���U�S�X�(v
�G�׿��#vEǰv�&��%x�b��h����U�7v    Ĵ{"�IV<�w���ǎ <2�Jy��&��b� h܁ѱ��?I���V��5v ��j��O�U\*i8v  ��U�U�V�k_��S�l���/��x��sΉ��W\��+bgt��ҏ(9��1��/�|��1��    �ä����V�ٷ���� <�O�>)��������u$���s�6�V�; ��R��ĸ �N�_�#^%_�:v	�P�N�=��3       <�D3�$���v�b�  6I�'�}כĸ��0pF�t/��<T��n�塺8�}]Ҥ�=  l)��n5�R���)���g�!͜�      ��%n�p=���iӶ� ݮ>P=0q]/�I�[ ����+�|i�y^��� ��g�خ����|��z ���P��#�?�9v
���*��R��      �?q��|����͎� �����/�4%v��T� t.{U^��*��z���k �[�T�s���\sc�  0�׿V��cU:�$^��(l�,i���c�y�Jo�;5v
      ��[Rj�,��U��� ��g�خ^����_�@kc����&f?�+�W��^���1 ���i:�(�˒�/ ���O���_;�e���J_:W6���oK-R�ɯ�A�       �j�˾�����U��䱃 ���T�;��_��ɱ[ �>��3ـ�}���]u�L*b7@�q������))��  ��׬Q���U��b�.O���$Q���T��ҽ�Ʈ  �z�#��z{bg c��^; �vTr�G�!}��KG�]w�� �h$�C��ϕą� 6w�9�&_R�| ���3�t����  "�ӟT?�0���u��p욇찃ʧ}B�W)<�  ��rK�   �(���_d�z׬�Y� �.��N6�H��= �7�M���� :A^�<���n�ĸ  H�ݧ�GH����al�}�����3       <�YJ�f��[b� @'X_��yH�1�b1n����7KI�,����v��!��-��K!v  h~�]�{��aC씇)�k��)���       ������,�g{b� @�����ʅ�(i��- �w �񒝕��%>445v �����R�}TR9v  h=��_����I�z씇��*}���ĉ�K       <�cs�Y��; ډK�Z����I��@�b�D䮗���/�xR 6C���Փ�M&�  �6��j5����c��*��]�3       l�]�.�T��Ŏ�V�!��<�ט|��R� 퍁;�,�]SՓ�_� ����	�+]
�{  @{(�;_ŧ?;�a�c���_�       �g��O����=Mw� ��V���$�I��i��P6��<���Y�*�c ����W�k7=���.  `�4�.U��o��x��J�~L�:5v	      �����_���c� @+����Yg��W%�� ����Z����-�J�U�C �dizT�(n���[  @�rW���xc쒿��~�>���       �̠[qM��>gN_� �-�V����7Jv|� ���;�z���yyH/�juZ� ����g���Ε�]�  ��j5�_���U�K�.9�%/xA�       [�$[��_C�Sc� @.��P]��,�	�{ t&�@�riA^�/�4�/v 4S}�z`V*����n  ����8�8i���%���Ai���       ��͕��Z���R)v 4K-�]��s�RI=�{ t.�@krוY�~�C�; ƒϞ=9��E��6��  t��f5��v�=v�$��T���5v      ���c�%y���; ƒKI��Lv�dO����1pZ_"�[s�_q�;�NU����~%���-  ���]���bg�]r�����       ��흔7硺���t������^%���������5�]Wei�̧O�; F�O��tY���%��  ݡ���Vq��cgl�ӣ��cW       �6�]�4�j!�; F�KIV�.L�/%��@wa���ka���y�ǎ�m1���,�Y���[  @�qWc�"�M��]"IJ9X��      t�g�����������:�/�41v����hO�.�"ճ�Z�; ����!O�Kٷ\Jc�  �.52������.�J%%��?      �C�s��<M���t��1 �%|Μ�<�%�4n���{ t/�@�2�_����R]�����૫z�kw�<v  ��\���'Hy;Eɂ��ɱ3       �����Y��>}���9 �x�J�y���]v����= �w��M���<M���.�c ��di��<��n|u�o�  �A����q�ɱ3���,xE�
       ��,٢zo�oj�*��hI>445K�en�$�5v H܁����d����?}����9  I>c�vY%��\?����=   ��8�*.�j�%G-/�      :�K��/������4v H�K����y�q�\%�M
 -��;�Yƹ���u��izP� �m$���ޛez��r�  ���x׻俽5j�͞-{�s�6       ;�zY��[k�z�ϙ��@���t�<�?��I�c� �?c�t�9��ZH/��;@w���K-T��Ⱦ%iV�  �Ͳa����aCԌ���z>      �17��K��~U�V_;@w񡡩Y���sIܺ�e1p:�I�R��Y��������|xxJ��&���_�  `K�ooU���ڐ�"��'j      ��ع(�r./�.%Y�����l��R�& x,܁��+٢����Z��d�� t�JY%}m��n�T��  ����"��O�L�(M��|       M���k��\^`,��}��L�s%͈� ���;�=f��+y�^�W���3�!쟇�F�>/> ����H��η���       ��fz_�����R}�s��Q0R��"O�I{���-���6���?���ґjuN� �V�<��K]v���c�   �&��&�^/`;.i      ��t�����W�4];@{�juZ-��I�r��/Ж�]ʤ�I�˳J�qO�b� h�,�3͒_�4?v  �X)>�)��>��;      ��v1�E��[�V�p�f���qy'���d�%��n�����n�2�=w�Qa�O��}�  ����{{��$;^R)v  �X�+T�}v��m�       H&{�~SҋF�՝c� hM.%�4]�g�[\�1ISb7��b�@��3��|���硺؇������b������	��   ��q�'��k�����&      �Ve.-H
_���C�  ��%���<����"�w�� ���;�4��K�,�M���874]�����BuQ^*�����^  Ѝ��#�f�~r��      ��z�Z��(~Wa�W��b�'�T_������zb� m�<�Yr}1��e��B�ʱ� 4�ϝۛU���7�&��f�n  ���җ�{�m�k�y       ���-��3�t�9�?v���CxnVI��Ϳ#i��= 0V�x��̗�!e�t���׮��̗�T��  �j55�8��GڤIM=      @[�N�Ey��,��}��@�  c'a�,�׹�G2=?v �5� 6��W���    IDAT���o���y�zb^���BuQ}�?0l  xdŹ�J�S��8�yg      hw��=��j!|�C�;��W�/�B��])�Y�{ �Y��;Ivv�z��J�-����hS>}���R}K���$?ݥ�	  �e�_���_l�ye�)      �Ŷ3ٻr��Y�~i�Z�9v���R2��Y%��(�rIό� ����֘%���R��Z���i�C�  ��g�쯅�Iyo�]2?�a;  ���K.�ܛsX/w       [�O�#��S�Y�2/v���s��eizT�[ٷdzF�& ���;�m1��KrםY����R�;�#���K�g�垻L�DҔ�M   ��W���Z՜�z�      �f�I�e��j!�,�T�;�#󡡩y%}O�~�]r�+鉱�  6� F�D��R���ZH/�C�?v�������"��,�k$��n  hW���sP�ܜs       t3� ��YHo�*Յ><<.v idpp�,���zc��>$if�& h���Ĥ�.�2�Y����q� �d��*����G.-�T��  ���曛sP/�$      O���<�洞�I���A@7z�¤Q�V�E�&�n�V���X�S�s��ܞW�w{?Ocl}��Jzr�~�ݛ^Y�[�&  ���?6�+�0      �1�o�%��,�3�4}J� ��y�ĬR=��
`���k cʥ�L�K��~S�3ʫV]m��n:�KI=��$[�ҿ��g;  �X�?6g���      ��%;A��P�A�3z�8�V�Z;�#!<Ѥcs�	�O�� ��h�ލOڂ<��河��g�ʕMZ� ��g�쯗{�ɥ�J�c�  ��� ��      Щ|�L�r�G�4��'��g�ͱ��v�s��f�ֽ�\%��$�� 톁;������Y%����.������<6�J�4}�:&7"yo�&  ��R�]        cm�\�T�������c�Unu_�Z��܏�׮{�I�c� @;c� �	2��G�!]Q�_P4���s�b��d$M�`nG��c��s�   �Բ�       �,&i_��͕|:K�o���ʫV]���C|������P������ ���;�V1h�ťR���P�Jҹ����v�=�b𡡩y^�B����~   �d�      t#�^�#]vd�_��sr�&�\yw�2 �ʍ��E�G�#���4.v t� ZMb�HzA^*o���j���;e�7m�r�$�h><<��e$f�z��2M��  �P��.       �؞�Sʮ�d!�Nn��W�{����R�'��r١�����N��@+o�|���k��1�E��WʫW_kR;����Y��D6���  Z��y�       h���d�W^*4��
��ҷlժ����R�VwWQn��%͊� ݂�;�v���׻%��Czf�N�~q_��]��V&h+.��!<ۥ��Q;  @˳���	       Њz]:�d��H-�W��➾�o���9v��jCs�L�J�$�b'@�a��M���Dvd�z͟�4��p��o������Y�8�����Z���-�]�H��	   [��;       <�q&͗k~>R�e!���.�)��=��;x4�0j?\j<!v t;� �ݴ���׮[�����vYo�ߵ�+�;�����S���tP���'����  ����b       @;铴����K�S����L�7�Kǭ\yk�8t7aBM�?1;�\�i�& �C��$S$f��F�7�t�y�Ҟիo41-�ث�M�b��V�x�L���   :D7�      �V*K��]�&ҩY��.������S�g˗g���|������暟K&�vrE Њ��T%��4O�,�BX��~�nW�e�l��b�3x�̬\�Ǥ���bW��  ����       0*\�%-Ld���Bz�ɮro\ջz����<�	u�9���)�?��)�B h�t���@�z^d!��fW&ҕ垞��;Fb7�=���5J}�+J�����>�ɇ@   nҤ��|e	      ��L������%�Bz��W�ٕ��߷U�����R)�Ӭ8��r�9�z�� �� �Q"����4�ޝgy=�_���\�����Gv��bG�5���꽽�,�<��{��ޒ�n��c��   �D6cFs���       �i�dǛ��\�,Mo�t��kE��W�;���r^�<E*=���ʥ��b*Sv h�@*K>�d�L���{z��~$�������+V�����000�$ɳMz�d{��n��I^   Lߡ)�8w       x�k�����6��~�d?��k�(_߻�_�T�������)�Z�Y��Y&^.=K��Yu @�a� ��,�&�L�i�j!]-��nHT���$���wo��m�����SݓyJ|�\{K��  D6n�l��	�����?�.B���wo�A�      �̑|�d�Y�Pҿf��I~�����Ѹ�֬�/v$��K�l`h+5��}���g�SeJ,v `�1p��`RE�|��Ly��,To��涼��>�:[���حxd>{�����n��m�\���^��Gy ��J��v{��$�@���Տx�TpL���U����9+�7�       ��$�%�^�Z�'��]d(��j�n�]s�-�:�%��y=�����И������č�L������ �NY�]����Jd�%�Bz��~Q��"��2�u��ɿ��˳���«��yQ<�=y����溴G>R�L����  �̟�ҧ?%������Ȟ�<%G������쳏4iRs���        ��/2�K�x������~%�_���r_�-v�����-\*ժ��(�&n���\�=%_�fKT~h� �v�`����ܴ�iӈ�]��u�,���iyQ�7��w���r�{��wǚ����%ې�i��/��\�9���Үy�;J�ئ!;3v  �x�CU�c�J���,��������Ieh%v�!�;��      `,L�t�LH.w)�)��.�Z��r��I�5J����Xq�I���V𡡩y�s<i씘�q�]%R.�>N2�Iw� w {eI��k���$�)�ɕ��o�n3���ߛ��tgb��GZa+W�1r{4>sf^�tkTMɐ�g��Nn�S�Sv�swIƋ�  �VK�:J�H�͸d���8C��K���ǡeX���5����      �Y\�J��u�d�.|/��4Ϥ;\�{Sr���QH+���$�s��w�1��?�>}RV�0TR1T��.2��r�#Ӝ�ޘ�d��]b� �R� ��$��=6~D2%��R.)�zIwJ�[�5*t���q�{����XSO�{��Z[�j}Ŀ���3fl���gj9I*����}��x��r�!Y�����4N*����\�  FQr�a*}����ob;������C�ư�$Yx���ۼ����       x4=�v6�����q�`*�� ~���VI~������VܓH�5J�{�zz��o�sܿ���s������Y_}FR�'���w�7Y�K3L��M�SCŦ?������  ���; ��	��$�I����M�g*6�^^.\�LYH3I�$������L�V���}ĥ���䖻k�����Ö3I��E������Hz%��a���d���m�T��S2Q�rM�4U�)�ciJ.�˒T��9�^9��  �Y���T��}TJ�-�sm�=U����x��:o&�x�&)yի�z���oM=       �Uz$���/�����7�\�M7�7j�B��ɴVnk%_g�u�N�����Z"�wȓ�_��ٻ�(K������Vݪne��I�3�;�wΌ3�w&��(Q"q�F��hDp51nQ��ƨ��+₈��+Fc��(��ƨ	J#uouˢl�U�>�� *K/u�u��s��z��9�9�>�;O�6� �$7�Zo���a)�����a�/ex����z�R�\:90�Xk9����Cj�%9di�M��M�p�6����=�[�� �j�&�\�#v�u�0n���G?������x��an�$�S�s��5��{y_n�k�� �qS�s�̜��4n�E�aK^����L#�	�y�㓃^�K��;    ��)IM͡��)n�p��Uǭ���Ncx�1�s���3J���b�}�m ������ ��}�n>   �A��c�u�����#��3�p�Ϩax`fN>y��v�R-      ���  0Uʆ�]��:���7��t�+v&�s�����̪�[o��;      0��  �.7��q��?<�g�+9��=��=43�4x�=I�3p      ���;   S�̮�k��A��y�I�v�?�6f�������\�w      `��  0U�w�3�s��ϙ����=�1��Y=���N礓��pc��      3p  `�^���+�������.H9�ȑ���9�Iw�_��S�z/�      ���  ��r�5<���Gr|�W�*3~(�����V��SS~���\}ur���      h��  ��S��,����Fr~ٰa�K�~�H�g4:'<.3�M���T��      Z3p  `*կ}-�O|br�M��ࠃ2{�Y��������q��i������sZ'       4e�  �Ԫ��,�މɎ��`v63�~uf^��������2s���Lӎ��/����i�       К�  0����M�O>%YZ���N��k_�t�#��}S�s�̾���|�����	       ��  0��g>��S��,/��Σ����79�����)�7g�w'�:%���3�ԧ[g       4g�   I��(��>m�#��K�5���D������`|pf�>+eÆ�%I���ߐ�3       �3p  �݆�X����֑�Q6n������1�;���s�I��_h]�$��]��>�:      `,�  �m�����y#�g��̜��̜~z2;;�{�i��e�]�L��_l]r��g��'       �%�   ��睗��^6�{:'<.�g�����#��$�nf��?R���%�����?���       c��   n��mo����G~OyЃ2{�E)�����j��g��H9���%?Rk�'�pغ      `l�  �����v���)?�s�����y�s��?�����ޙr�Q�K~����~��3       Ɗ�  �����_��_4;��s������q�������?���.�1uq1����u      ��1p  ��08�5��_��]�L���I9�U�o�qDf?�����[����0�S��\}�      ��3�:    ւ�_���̤��g������ޙ�;ޙ���y�}���0��>3�=/��~�u�O��ͩ_�b���R���ԋ/��7�<��    ��f�   {hp���Z�yֳFY)�tbʯ����ן������kܾaC딟R���^��� �mx�Y�uV�     `uZ   �Z2xի3|��V�r䑙=��̼���ᇯڽkU���2{��rܞ��3x�3����%       c��   ����We��7�ꝝ�O�s��G&����kE9�̞����Z�ܮ��^�����       k�   ��<-�7�yu/=��̼����ȇS��Yݻ�\籏���ߖ�_�:�v�??����u      ��3p  �}4xşf�������?���~�̞~:���V�a,p@ʿ�w����f�5g$����nW����/l�      �&��w~  `���I��Γ���w���Rf��K�YZJ���d�����d��S��:��R��&��䚫S��&��U��c���a��zhr��~xr�a�����S��3�G��3��h]|�n�)�'?9پ�u	      ��`�   �i�?IJ'��?�M@��r�{'��w�]}�Ν�F�?�Ar�ɍ7�^}r�����v}|���u�'�oLv�L���}����7����KJI>x����ɺuI�rЁ����A'�r��'�xЮ�:h�����)���3&��E/N�ַ[g       ��   �/{YRJ:'��:���ͥlؐl�p�/��(�}2�������       kJ�u    L�Z3x�K3|�;[�0�w���=�u      ��c�   +��^��i�>�v����''7�к      `�1p  ��Tk���>�u	��������       k��;   ��Z3x�2<��%��������o�      �f�  �(Ԛ��^l�>E�7���K^�:      `M3p  �Q�e�~�٭K�����On��u	      ��f�   �Tk/|Q��~w�F�������/o]      ���  ��՚�^���i]����?~Q�      ��`�   ���^���9�u	+�^rI���u      ��0p  ��r�����[����2�'��,/�.      ��   ������\#��n0��3���m[�      ��b�   �m0�=r�`����?K��Zg       Lw   ha0��9�����.a/?�����       ��   Z2x��3��C�K�C���2x֩I��S       &��;   �4dp�F�k����tRr���K       &��;   �v�K��h��������n�      0��  `,/g�ԧexᅭK������      `�  ��2x֩~���%�F���^���       S��   ���rOyJ�}�u	Ir��<�����[�       Lw   7��<��~�Ƚ�n���NH���%       S��   ���r�<9�O~�u�t���,���ԯ�u	      �T1p  �q�{�^?��%�媫���Ǧ~�+�K       ��l�    �N,-e�I'��G%�3�k&_�~��ɕW�.      �J�   0�v����m]       #�i            ��;           c��          ��`�          �X0p          `,�          0�          �           �w           Ƃ�;           c��          ��`�          �X0p          `,�          0�          �           �w           Ƃ�;           c�Sk>�:          ��Vk>ޙ;�G��[�           0�j�Es��Gw�7��sv��>��\�:
          ��R��ͭ_�Ȳe�͝$)�\�4��=6��i          �t(5��m���r�;��s�H�~�	)9�]           Ӡ$�ݴ�w�%�,��k����A��{bj�^�<           ���f���'?1pOv��{'&y�j�          0-�y�~,�����{�{���#o          `J�wt��;nO�`��$%��~��I9stq           L���n�I%��g���=�e�����~��           ����~��;�'w1pOn�����׮\           S���{2nO�`������zϮ%��           S��/�������ɧ�����ދj͟�[           S䌹��s�tܞ���=I�{\S^��_          �t�)�����`o�n��I2�_xiIy��|-           ����>�_x޾|�>ܓ��_8��          �[�ԗ�����3��{r�Ƚ�Ӳ          ��QJ^����d�د�{�t��W�����9           �M����^��{�~ܓ���&%OIRW�<           ֆR��n��ʕ8kE�I2��9��          `J��rjw��g+u��ܓdn����rJ��J�         ����    IDAT �X�Iy����_��+:pO��Ņ�&���          L���g��^�����=I����ה�'��|           ��)y�\��(��=I��響'$Y�           ��AJN����4�F6pO��~����q1r          X�n��k���t��$���k�O�4�           Xq�Z��z��G}���I2���)yT��q           +bPS�0��p�j\�*�$���>��G%�y��          `��<v���պp��I2�������          `���5��p�j^���$�ݺpQ���Hr�j�          �]�9L}�|��j_���$�.^��2,�%����           ܮ���\�����M�I�ݺ��R;��;          �8�^R}]��?[4�'Iw�/���\߲          `�m/%�����n�t��$�~���F���-           S��Rr|���l���$����Z���[           �ȍ�S���z�k����=I���j���$״n          �ז�c��:�c3pO����K�zL��[�           L��S�����u�m���=I����O�1I�j�          0�~�Ny���[�����'�\�����nm�          0A~��9vna���=c9pO����o&9�&��[           &���S<�x�W[�ܑ��'�|����zTI��[           ְ��Ny�����Z�ܙ��'ɺ~�ۃ��J�k�          �m�Ù����:䮌��=I��z��<< ɖ�-           kEM�Z����~��[�Ě�'���[����I��u          �pE�t8�u�?��S��������oڴ��3)'�׭{   �T��S�<�u weݺ�w����9�� �ov��u�a�� �q�CZ'   0]�7����+��:do���b��MG���߻u  0:����9항3    `M�[�d���:  ��s�p0s��m��n됽�i�/����.u��5�T>          �*�2,�����'I�r����Σ����-           c�_�K�~۶�Z��5;pO����o�G��[�           4���N9�^o�u��X��$)۶}�����$_o�          ����f:G���k�����=�=r��yPR�ں          `}�۝=��+��Y	1pO�����;7wlJ�Һ          `���p�r�勭CV��ܓ�l���n���I�ܺ          `����zLٺ���!+i��������&�R�          ���ݒcJ�U됕6q�$)������1����-           +�\��cK�wu�Q�ȁ{��m�n���O��-           +���޼�貰pM�Q�؁{�{�z|�϶n          �۽����5�\�:d�&z��$����M}D�ϴn          �{�o�;wL��=���{�{�~���k���-           {�~������UW]ߺd5L��=Iʥ��;��G��#�[           �JM�T��yX���Z�����'I��7v�z�cJʅ�[           �HM��\'�Qnjݲ��j���2r��o���n          �I�䢹��GN۸=�{�{���?&��i�          p��|ln��G�-[nn���Tܓ�$�n�����Ӻ          �&�;`��˥��h����ܓ�#�^9�u          0�J򁹍5���d�����b��$�j�          L����{�S.�d�uHkS?pOv�������u          0U����W���!���}���n�����ٺ          ��=�~���1p��]#��g$���[          �IV����_�A�qb��v����J�_�n          &Q}k��prI��Kƍ���(I���N�%ֺ          � 5o������>�;1�뽰��i�          `Լ���{JIj�qe�~�{\S^޺          X�Θ3n�K�{`���Ғ���          ��SS^=���A뎵��}u���          {���>�_x^뎵��}/��W��          ���k�����^0p�K�~�եď           �PI}�q��3p��^<5Im�          ��R���~��;�"�}4��)5O��;          �[�yQ�����k���~�[�%���dغ          h�������i�C�2��4���֤�#w          �V5)��-�^�:d�3p_s���k��Z�           ��&��s��׵��+d���zB���-          ���I}�\����!���}����%���;          L�aJN�����:d����h��͏)5�&�n �iQ6oN����:    ֦��S����   k� %'��zg��4�#��y��Ú�̷n          V� 5�7��{w�Id�>B˛7?|X���         �$�Z~w~q���!���}Ė7��a�^�d]�          `�-�Z~{~q��!���},m<�?�d}�          `���5��_�:d������|P�ԏ%9�u          ��v������n2:��Ew���K��Z�Z�           {d�0�7��W��W�ҦM�)Orp�          ��TR�[���t�i��U����XR�K�u�[          �۵��>¸}��7����6�<$�Z�           ?��R���~�3�C�Qi0�vn���)�O%9�u          �K��]X���!�������6�Ǥ|:��[          `�][J���z�:d�uZL��~��SrL��Z�          ���6%3no��cb�ƍ�I)���[          `��0��й����:���cӦ_H��%�غ          ��2�<tn�_i�.����|����zTI��[          `�]Y;�������}̬���=(9�$��-          0��_;�!�_k+��}7m�p�����ܫu          L�mu�9f~���:����1�~��-�:|pR.k�          ���n�Ù���/�1�~q��A�N��-          ���d�v:�2��{�h��+��k�7m:r6��$�n�          k��N9z��¥�C�s�kD�ǽ6,u�?����n         �5�{Ù��뮸�;�C�k�kH=∟]���lR���-          �\>,�~۶�Z��g:��s�����]^~HJ��u          ��-������k���s��=�z�          S���)X�u��!��5�l�����̃����-          0f��4�9ꀅ�^��^i���?�s�.�L��Ӻ          �����٣��/�a���q�^�:di��'����-          ��7�Kݣ˕[��a�uZ�ʖ-?쮛h�/�n         �F����+��k��'D��=Z���hjԺ          V��wK�-��խC�^p���+o�./?<��Z�          ��(�t;����a�>Aʶm7vS�Orq�          ����l�ز�pM�VNi�ʫ�6����$Ǵn         �����7�Z���Z�����>�J���{���k���-          �¾�ݹ�8���d�>�ʥ��;��G��#�[          `e�/t�vW�����%����+�����CyLI�p�          �/%��.-=�\y��S�	�k�~�ǖ��n         �}QS?�-�8���WZ�:j2��i��I���-          ��j�'���Y�l��u���)Q�A��BJ�i�          {��|ܸ}��O�����Ssv�          �35��܁�e�>]ܧLI��މI�j�          ��Ԝ?�qãʥ��h���*�h�&ei��3�<�u          �������J��:����)U�������3[�          �n�3n�n�Sl��}�I}}�          �]9���`�>�ܧܮ�{�Y)���-          L��n��wv���z�Skɟ�n         `�Էu�O*ɰu	��s��^敭;          �%����b��-��1����;          �p5o��zO6n�J� ��Ҧ{�QM���          L����-���:���wnW��pzIy~�          &KM��v�ܹSK�6�aMyU�          ־�������`|�s��6o~n����          �]5���~���;o����n�wFJ����n         `�)�/3ngOx��=�s��SR��}         �*%/��z�h���`��^ٹ�OJ�o���         �����^;X;��k;7�������         p�jj�3��{m��w���M�NL�[c�         ���I9u����!�=���6�vIyw���-          ����g���oh��d��~ٱi�o��sb�         0�jR�>�￱uk��;�m��͏)5�&�n         ��aR��g��6wVĎ��|t)���         L�AJN����j��g�ΊY޼��Ú&�o�         ������{�n�d0pgE-o��q�N� ɺ�-          �Ԡ����ŅsZ�09:��,�[.*�<2�ͭ[          ����vV����M�~��\�d}�          V��Z�o�/.|�u�����Y�x��2�X��Z�          �"v������n�d2pg��6n|`-��%9�u          �e�0�1�����ar�3rK�6�rM��I�[�          �ɎN�o��zm�d3pgU,m����t.2r         Xs�������?�:��g�Ϊٹq�/�t>���-          ���׻��ŭC���L����K�zl��[�          p�n,%�����YUs���N�1I�j�         ���t���^�s�C�.�u �i����!5�Nr��-          ��kS�^�K�C�>�4�c����t>[���[          H��0�򰹅�/�a:���͛6�ۙ��k��u         ���a��_��z�WZ�0�:��n���oJ�*I�u   ���w�a������wU=U�=�g4A3��D��66�	�(la���8�����&�9��`��x��9�`���p c�<"h4���t��h���]]��+��骻���y�����5u���      ����f�Nn�d7�n�[K[S�D�         �!�������{?�;R� ���^����Q]��         `H쫺�[[�{��;"���2:9����#���-          C`���o1ng!�;ΉM���G�PD\��         `)����^�����ݹ[���΂3Z�{�Rl��{r�          ,A{�Z�&�v"/��`U���S�}(�zl�         �%bO�^�ed��{s������U��o������n         X�v���[F�����c�΂Wmذ�So|0"���         `������2:=}_�8�Z� 8�4=���uo����n         X��:��&�vw�45��h�o����         ��|�S�mk�'r���0pg�H{�<P��Q�'r�          ,_��k�,ۻ���*���U]uժ�ə?��o��         �@}�(��ݻ's���0pgQ������-          �g��nKey w�/w�jÆe�z��5w         ��"�m�ݾ?w\�Z� �Piz�X�#�ù[          �O��������<^DuGD|0w         @>i[QK��,z)w ̇��F;��O#��-          ����祃����w��41q��#E�7w         � }���y�q;K��;KFڱc�1��%)ҟ�n         ���bv�����#�K`�������g��JQ�I�         ��������������g�^�})Żs�          ̷*�_��s���Gs��|K��_��zg��ߍ*^��         `>TQ�y�V{q��8�����,Y)�[�ۯ���         �bU)>�l6�4ng)3pgI������{�[          .T�����i׮��[��R� �*��ٴ�7#���[       ��+�ĉ�?-w��FĞ�LT�ʝ�MQ�+����8p ��org  �0)�76n|yڶ������; !E�����Φ�'"�͹{       ��/zA̾�U�3.ء�?����G�3�;%""Fǖŋ��uqb�չS�{p��; ��"���q�+����QUe�-�M��"����      `p��c|ͺx��+z k�%�7�K_���j���  ,
�h��W��=�;��; )ETE9��H�˹[       ��7�k����q�e����1��7�ո �s�?����a��P1pg褈�h��)~)w       ��|Ūx����^�����ħ<#^��7E�52� Xl�oe����#w�R�����۪*~>w       �U4�q�]��g�����W����ϻ3�{�K�V3�  �l��,ʉ7��^����&�Zk��3UĿ��      �`���7?'���/�z�޷{��V��eo��~�M}� ������,и�af���k��UE�7�;       ����x�k�c˖��٫V���|���5�>v�� `	�����;DDD����)�O��       `�.���x��k/�0ogn�lK��M?���8og ����b���)��������/���e�       o|�%��������_�Y�?��׾9�-[1e  ���,�o6n�����e��)�?��      ��5���ޗ�!���g^�倫�۟yK��%��FQ�s  KQ��i�m�Exw�E���"�?�K(      ��S����8�{�K�V������x�_7?���R�c!  KE�/�ʉ��w8�f��_"ś��      `(=�)ψ����j���g�Ɩ��_���'<y e  ,��˟����;�F������FD/w       �w�5�ū��#�j����̺���~��eW\9�2  ��������4''~#��      `X�[i����o��߻���Uo��X�j<C  �QJ�3EY�������Y4ˉߌ��F�       CillY��5?��������x�+���H�2  �T�O������; �fY��̦M'R����      :�z#^�=/���blly<��ȝ ��QE��VLN�r�Xu�����3�6�R�?��      :)���gݖ; �ť�H?ڜ��s��bQ� �I�,�Q�xEDtr�          ZQ�H�4n��a���n���;         pU��'Ͳ��r��b�� �Q��~����'zU�qD�r�       �[�_�C����` Z���N  X캑�����������.P��~������ժwG�H�      �~JG�D����@q�P� �Ŭ)��l�?w,V����5�&>��tgD���         dխ��:�v�8�p��ɉ?OQ}wD_��    IDAT���         dѭ"��59�C`�3p�yP��_���܈���         `�t�*��*'�G�X
�a��{�.U��Gđ�-         �@�VQ�՚�xw�X*�a��IQ=/��        `���E��VY�'w,%�0ϊ����s#���-         @_���z�HY���!���Ce�����D���-         ��:���c�,ߛ;�"w���䶈궈�?w         0/��/*��r��Re�}�,�OG�gGā�-         �E9�R�Q���K��;�Y�����F��s�          �X�����s��Rg��l�?WU��"&s�          ��PJq[11�7�C`�À�&'�Qݒ"��-         �99��������!0,�a�Ze���C#�v�         ���Z��91���!0L�a�F��+�Zښ"&r�          ��@T�ۚ�����2���g�׽)"ݗ�         �&��Z��9��S�C`�C&�SS��Uwk�ؙ�         ���}U-�ښ��|�V������nUm��{s�         ������[[_����2-�=sQm���[         `UQMU��-��_���������[t��"�ݹ[         `��j��ZSS6|� �����*�fo���_         0{z��֑���C�������.��n��/�n        �%nw�[�:�wｹC�����4=���uo����n      ��R��F�; ��۝�:2�gg�����������͑⓹[       8�Z�W?��q��-j�z�  ��=s)n���/w�H�@�={(������[       x��يko��X9�.���+�J��rg pf_����c��D����aK�v=X��n����      ���Y���1�|�7��j͆���'d� �,�ҩ׶�ML�s� ��� �Yڹ�Pu�U�휜�@D<#w      ��[�bu\��o�F�|��.ٸ%fgN�Ԟ{�񵪊81�H[��E��y �S�RQ4nm��=�;83wX�Ν��n���7��      V+��ŕ�?5���O.6m�.:�3q�Ԟ���UU9>;��ڲfԛ��� ��|��uoK���s� gW� ��4=}��ͽ0">��      `��py\����q��uW\sC�^�q U  ��g��������a�0p�E$MO+��#">��      `�l���r�#�s�Z���Q�=9��\��2  ��3E�g��<�;8w�Ȥ�<^�ҋ"�r�       ,u)����'��+�?�߭��q�c�#c��P ���mE-=;����.Ώ�;,Bib�D16zG�xo�      ��*�j��<9�]��>�Q4�17<#FF��/ ���>U4j������K��g��Tڱc�1��%)ҟ�n      Xj�"��o��u�.��fk4���7EQ�P �Y�}q��iϞr� ����}�lc|�])�{r�       ,Es$���;b����v����O�Ψ�L5  ����������s� Χ&X����K7ܕR�;w      �b72�"��g�貕�~��K��O��H)���  TWtf��8���8����K۶u���:�6�^Dze�      ��h��5q�c��Fѷ;.�ty�Z#1;s�/��Z�j�gO���}w�� �%��s������N.��;,)�[��k;�7���W��      XLV��W^����}�k��u}�#"�ı�Ѿo W dSE��T�3MO���̏Z� `���n�n�>"~/w      �b�v�q��Oȸ ��S��@����41a�K��;,1)�[��7D���n      X�6\vMl���H)�N �<T�oŋӮ]'s� ������+��#��r�       ,D)����c���N �<U�k��~�q;,M�D���(�o�H���      `�_�)�n�"w  �)U��_�v����;,a��'�Q�J�      ����v�/�˝ ��ygc���m['w�?��=4r/,R�R�      ��db��x��d�  ���,��+S�\����a����n�����s�       ,UUŮ�|&�>�; �3��GQ�_e�����Hk��3UĿ��      �P�zݸw�'�ıùS  8��[EY�:Ets� �a�C�U��U����       X(�s���ŏ��̉�)  |��7�r�RD/w	08�0�Z�ĿN�~"w      �Bљ=;�����ur�  Q�+���a��Ð*ʉ_HQ���       ���G�޻?�� @VU�z1��a�vN�0Ċ����?��      �P=t��ʧ#�ʝ 0����͇���AC���\Q��1�����      ���x��d����  C���������e�D�n��H��0r      �����cj�=�3  �F�/�ʉ��������f���Q���^�      �s12���痻��O���  |}�^�D�`a0p��99��G�#w      `k���5�����ϊ��X_��s�������z �0KQ��q;�p��7i��Q�)��     �&��7_�?��X9�.j�z\q��zgUU��˟�c��� �a�R�lQ��6w�����,�߮�zUD��n      ��]�2��g�eW=.j��7��r|}����׻{�n�{�'���}� `��*~�h��}�`�1pN�U�o7r      r���q���uO�)Ɩ�>��\~��Q4��1י��?�ٓ}� `TQ�ۊ���,L��i���U�WFD'w      0|��Z�?����+���N?qh��|�c��3{�x���ǣ;���
 p����c���/�.w��Z��;��#w      `@�"�x�q����e��;k7\+����,�ıñ��OF����. �%�����,'~%w���g�j��UKqgD��n      ���K6�㞺5.ٸ���kn�Z�ч�ov����뫟����w ,UD��fY�j�`�3p�I��~��^'s�       KO���������D�h]�͑���k����_��_�]  �\/�zc�,-w�8��11�g�Jw��;      0�.ٸ%�ԭ�z�Ƌ>k��bl��y�:����bz�ށ� �Hu#��e�;�C�ţ��XR�ɉ?�l���U��D�h�      `�]�"�x�l�����R�-��_��G��z�v���;j��7�g��������Q�����)�7s��@  N�U��Y�� w����(˿�l��yU�z_D,��      ,.)�b��bӖ�D����]�2�o�*�'v��٧�w����>t�'g�r�ʱf���� �<t�*��59��s� ���J�B15��=?"��n      ��+���O~Vl�����ۿnӖ���X���f���h�~  N���]�����)�`���GRTF�      �Y�델���ǵ7~G�����}�V�+�����|��n�^5��j)E�n� ,(�UTw�&'ޝ;X�|�.JQ�MQ=7"��      ,L��l��>uk��teD��ݻ|��X���1����ZDfL p���{r� ���;pъ��XT�["�`�      `�i�(�#Y�������������c��KZe���C���'`^4''�ET�E���[      �����=q���Y�7������\o`w���� p'RTw���{s� K��;0o�e�鯍��n      ���|>z�n����m��k7��������{J)���@� 8��)�e�W�C�����WͲ�L�xv�      3{�xL��j��/��	Qo}�cv�U5��{��"y� ��xJqGQ��,-���k�۟��޳����-      �±�}o?z(��Es$6=꺾�1�̸="��0�  �:�R��h�?�;Xz|���59����Q�n      ���b�W?U��r��K���k�v�l�۷��U���v  �C)�mE��׹C�����VY~���Ƚ��      XN;���e�=����Z��A��^�v ����-���,]�@_���W���5EL�n      ���_���ǲ�=2�<6\��y?���EUf�^K)�5/� �`����v�s� K��;�w#����7E�\�0       H�׍=�|>��/�&F�V��ss�{��h�{  �@�j�7'&>�;X�|�btjjW��n�;s�       �y�@�?�7��)�b˵7FJ��
�L�;og���; 0`DU��9����C���00�����U�5"���      ��޹=:�3Y�^�b<.��Q�v�\�� �������jN��T�`x���hYjkD���      �57׉��۳ݿ�Q�E�5z��t{Ut{�y(:��Rus ` ��n�����r� ��'`���ro�)n�Hw�n      �z`;�?���z�W<��G|����ɓ'�СCq���q��ј��=�9}��^��v 0���^�����/��O#w 0���]S����t�E����      ��{�c��K�^��a���_�)�O�����w`|���u�"{kd$6��$֯��W}�띹���Q4��������^���T��@^p�I��M��-�O�      ���9������^��f"��������8p��S��#"fN��={'�S۶Ŷ�|6>�s݁�S ���V��M��)�v �z�������׽5">��      �g_�+�>8�;�?���?����#����݃��?��عsWt:�{��Q7�  �fO�^�:21�#w0�|��KSS��F���S�[      �\��s���f,~��}��w�^��7��h4���RUq�Νq�ί�����Z�] �������<�wｹC ܁!���@�l�U|"w      ����Gcj �?v,>��?��G�|��G���H�7 �UU�`_��}�|&�R�0�  �bW�׽ytz����8>� Fڵ��b�u{D|<w      ����{���#g������/���8z��#�W��cdt�y�W������jǁ����x:� @|u���9:5�+w����,(i��C�H�9��[      ���z��s��#����_��s1=]�����eQo�|^�a�{��nw�b�Ψ٨��l `(}�S�m��h�x8w`�I;w*�s�E��      ��������~n�Ӊm��Ynt���Hg��^Q=l�ߙ���������R4�f ���rQ4�.ۻ�?�x�>� R��>V��^��      ^yߗ�3sr^ϼ�ޯƱ�G��s�z#Z�cg��^��W��OOFu��_�F��z� :_*:�ִ{�d��S1p�4=}��ꎈ�P�      `��ݹس���z殝���϶F�G�^?�Ϝj�ޙ��ѣG�7�
�� ��ET�J�wM�8�~�-���"�E�_�n      ����x���<,ZUUL��u�?�R��e+��3�ީ_T?����I;'͆� p�>S�xv*��C �ħ`�Key��#E�7w      0X{��Bt�:}�ɓ'b�3s^��(ZQ�FO��S�����f�I)Ea� \�O����nߟ;�l|���c�Lc|�KR����      Ngv&���}��?z�~otlE��#�UDTq�������)�� �PIۊZ�-ML�����w`�H۷�6�W�4EzO�      `pL�#�.�ѹ|>�j12��_��N��{��]�]���z; p���8y��v`1�	XT���K7ܕR�;w      08{��\TՅ�ǖ-���m�F�Q���k����F�u��]�F��� ��h1;�t����! ���XtҶm�F�}WD��s�       �1s�X�8v�tlY�t�C���+#��gطG�l^�=��,��z 0�G����ҁ�(�L܁E)Et��|m����-      �`�2z�ш5k�]���j�}��^Q����/��GܛR�k^p �C��-:3�O��͝p!܁E+Et�v���{�[      ��]�2���E��+����o�.�z����oO�b��5u��� ��UQ�E���ہŬ�; �b��nU���ٴ������      �c՚}�Տ�.>������[�:�N'�4g�߰)��Ϻ��U�^�z��^p�=y"���=o- ��VE���f�δk���- ��X�RD�k#�����=      ��[9����X�v]\}�u��/]��Z=Z��i������K7_����ı�Ѿ/w 0U�l5�׸X
�+`IHUQ���~5w      0���F,[�z^�z�3n�z�?�^yգ̸ U����F_l�,������}�կ�n      �ϊ�u���LV��gm�}^�z��+VƳny p&��w5/�xgڱc&w�|1p���F��E�_��      ̏Uk���y���	q㓞>o�5��x��7FG���L �s���d��i۶N���d�,9)�j��o�R���-      ��[9>����g<sk|�M�F�tQ�,_�2��e����o 8�we��)b.w�|k� �V���3�n�?��      �0��VF����Ox�Sc�������U9|�~7�W]����cdd�/}  ���^��1n�*w`IkM�vf��z��'s�       �o՚�����QW�e�o�/~�3���o;�нV��e�o��>�;c��M}m 8��)ʉ�O��! �b�,y�v��f6o�R?��      8?+��;p����q㓞7>�iq��}�g׽q�Ѓq���9˖��e˖Ǻ�����*Z���( p�(����ہ���
�v��g6m��H?��      87�z#���k/Yk/��� �<��(ۯJ��! �V� 0(����*�/��       �͊�u��i 0�R�*��+S�\��A�)*�r�'"ү��       �nո����R��1�~�q;0L܁��"���xkD�Z�      ��V�1p �W��O7�̸6���yh��~KT��[      �S]�2��H� �,�h���<m����0h��PJU1��'Q���n      i����!U��@s���I;v��n���Z)�WL�����      |���� �P�Xsn�i����! ��C-Et��կ�R| w      �z��V���  ����iz�X���܁���o�mV�K"����      D�_)�4  C�+Ew�9i׮s� ��� @D��<^�<yGDږ�      �ݪ���  ��N�vK��ޗ;`!0p��t���"zύHw�n     �a�b|]� ��H�nw�e{���[ 
w��Iey`��G��r�      �0]�2����  �p����>:=m��0� �blb�ݫ�۪��r�      ��Y9�>w � ���sZSSw�.Xh�Nad��{�V�="��      �d�w `ɛM�{i�,?�;`!2p8����R-�3�[      `��X�r<w @?���.��/s� ,T� gPLL�M�k#���      ����"%S `	���[��;sg ,d>�E�,�)ޒ�      �����s'  �MU��7'ۿ��`�k� X����ټ��T�O�n     ��j�����5י�ٙ�/��Gs'  _���e�gsg ,� ��n�tg�e�#�7�n     ��ft��h�Fv��{��/v 0����5��ק�*w�bP� �X���('~����r�      �R�r|��*�<�`� C��Q}_����X���1ל�����L�      XJV����ؑbn�3�� �a��+�:ߓ��x������<�����+    IDAT�E��'w      ,�z#���}���] ��:؋��Ҿ}ӹC w��vz��Gă�[      `�[1�.R܄��� @_uR�����Wr� ,F� �5�g{�j/����-      ���_?��:�3q�衁� �*�xc�n8w�be�p�ɽQ�P�      X�V���]^o �)����d�rw ,f� �Y��UE���      ��ht��h�Fv��; �?��v��� X���A�,*"ޙ�      ����vWUUq��� *]\��)�����̃Q������[      `19v䁸zOtfO����G���l�� �M���ꮴm['w	�R�� �T���Ֆ-�3י�DqY�      X��?��?""Z#c�j��X�f},_�6R��w�=�o^� ��#U7�(M��L�<1p�Gi����M��;"}$"�r�      �b2s�x�k�}�Q��cŪKb���r|}4[�}��� ����R��1����C �w�y�,�O�l���T�;""��     �Ũ��ơ��q��tD\���s��8~�p?R�a��5����� Xj����n�����OLU�T�      X
.�u�C�ED��P `X�n���/�# �"w�>i��?�ٴ����+w      ,%����: X������ K��;@�����̾�S4���r�      �Ru��ݫ��#ȝ	 ,��^�δc�L����������GOl����Z��qI�      X��u��e+cl�����f. ���Q�^�����X��7� �W�SS�RT/��n�      6'�������  ��?ܜ�ܖ;`�3p��,?���W�;        ��◛����� � Ҙl�_)�rw         ��c����"w��0p�Q5:�o����n        ή����k/M۷��n� ���?�K��q(w     �o��>�����sf���B����=��@�`K����_k�K��իz�Zl����K�բ�zY*
?�FE�&��$ �$�	�YB 7{sΙ��fI6�ݝ9s�������������y<��u%����k�Ȝ����  �1ZQ�������! ���`�m���<������-        ������~��� ��� ��~��5�+�;        �GR�>��}cv�42pH2��,">��        <D�[�/�� �V� IJİ�:�����        DD��:]X��c�! ��� Q9p`�U�'#b��        S����/.ޖ�0����{�������        S��s��˲# ���;����_^�^��        S�v��4; w��P"Fs��OF���        �2���3?Z����! �����.u���f�        ���Q_�ei�]� |��;�i/.�X��<�        �B�����wfg �����\������        h���v���]�73p3%b�Z�qov        4�r����?��73pC�z�n���        �L���z�[�+ x8w�15��}oD�Qv        4I���v���� ��;�kϵ)"<)
        �D��J��Q�[ xd� c���s�[?'�[        `���K�(;�Gg�0����ZJ�,�        &Y��{�^�� <6w�	0��&"���        ��T�877�� <>w�	P"F����jv        L��(�'ʞ='�C x|� b[�۫��Bv        L�R�es��-� �w�	2��}[D�3�        &C�q��{Mv '��`´��/��}�        0�����K�0;��g�0aʞ=���/����        c��K�..��� ���L�v����zqv        ��q�\�wiv ���`B�O�xiD���        �1s߰ċ�# Xw�	U>RJ�����-        06j�d[���� `m�&X�׻>�^��        �F\5�ػ,���3p�p�'^��;         �}�/ʎ ���L�r��R�?ED�n       �45^����fg pz����]Q/��        �5⪹��e� �>w��h�8�����        �M��0��eG �>��>|dT�/fw        �檿���ߟ]��0ph�������        �M��v��G� �w���m�_�ew        �[����)�� ֏�;@Ô�{�įew        �F�Q^1Ͼ�� �/w�j�zo�(7fw        ��}nn���# X� T"F5F�%"��[        `��Jԟ){���`��4�|������        XW%.n����� `c�4�\��""���        �uro�֗eG �qf� �8��=>�q�k]��     �d=��x���eg�	Jݚ�  ���J��eW �q���������{j��n     `r�3ό�mO��`�f' ���d��Kv �� �����"�hv        ��j���Q�C �X� S`[���D���      �t'��Ǐgg ����^�s� l<w�)1��:"n��      �I��Ç�7�..y����s `jԈ���y�;L	w�)Q"VKԟ�i     �S��ww\���Ž���6t����oϝ�Y 0%�/���?���a�0E���'"�]�      0I>��O�;.y}{��7���������8���$��T��\�yv ���`ʬ���x0�      �]�5>qõ���]���a�|8Ɵ]������F�^� `u�%��h���;�����uK�Wfw      �8[YY��\�����>�����1���V6� ��Es����# �\� Sh��zUD�;�      ��G���+_�������>���u����6� ��W�Q�Wv ���`
�n�x��߳;      `���{�o��XZ������^��5}- ��o�~�Pv ���`J�/v��F�Pv      ���v.�~��������8����?� �Vuw�߿(��� Ӭ/��av      d���M��>����bu08�뭬,�{/k���ס �O)�K�jv 9���|�������      Ȳ��W��mq�uWE�uݮ;��뮊�?pE�F�u�. 4]��@���Hv y��\{8���r$�      6�ѣG�mo������7���)���7���v h���h�ײ# �e�0���ҁRꫲ;      `3�����5��۷�������7�&:�����V.��g���
 r����nDl���     ���+�ş�������m�=�{0.{�����wn�=`�<�^]�?� �3p J�{<J�Fv      l�������_+�˛~����w^zQ�z�_n��`ܕ�//,ew ������h�zQ�I      �4�Ϯ|g\w͕QkM�X�?��q�uW�v ���?�j�~v �a6; ��P"F�R~�ָ>�     ��Ӻ�p����X�Q�Go�P�gl߾#;'""��q[l��������Ny�r�� �L���J�{<���P� /˝��%�ew        0>�����D��C ��  �L��?�        6A��_1n���&����#���        4]�x{q��� �w f8�,"V�;        h�Rʯf7 0~�x��KKwG�7fw        �L��{ڽާ�; ?%; ��T�o?{К�3"��n       �Q�u4���{��bv ��	� <�r�=k��fw        �4��v ��; �jn���_��        �1����� �/w U���K��dw        �o]Z�;;��U� o�쳟8h��gg�        0�V�u���..��`|9���T<Zj�:�       �IW/2n��8���U�9�	��ٻ"�of�        0�N���3�u��� ƛ�x\ei���U�        L�d���p�; '�v:�V"�,Q�g�        0Q��W�(,e� 0����I)���Vī�;        �0%�h���r�; '�>��g���Fę�-        L������uqqov ��	� ��r��5��;        ��R�v N��; �d��k#�hv        co8*��� Lw NI���gw        0�޽���rv ����S�����       �8sz; ����S����F�K�;        O�������; �<� ��hf�#b5�       ���*�� L&w �d���wFğfw        0n�����'�+ �L� �]�WDD��        `|��rz; kf�����z�Ԉfw        06>7�ؽ6;��e��i)%^��        �x�%�o��� L�� ��[�t>Q�?�       �T�����]"F�! L.'�p�J����        ���1n�t9���V#�`a��Q��- �T�_��/G-�G��m�z_D<Xk]����2=iT[O*Q���Q�������xzD̦�W      4@�X�;�)�ݻW�[ �l~��i+ueT^��!� h�k�[�����`wYZz�t/Z/�����=�����@D�ӈ8�k     �L+��������;wn������- @3���(��ZW�����k�`��Y#��9������k��������     h������ʁK�! L>w ��r���W�; ��v�D\5�z�|�u�X͌Y޾�oGk����#��     �1v�\���# hw �ͱN���(wE�lv 0Yj�b+��ͮ�\Tz ��[Ո����+5�gD|gv     �x����7gW �� ��Ag��� `b�Z^ݞ�7�n�xv��t:��F�͈���-      �ʍs���gW ���  ���.�  ��G�_l�������k'e����������U�#���     �L����n �Y����[YX����=� �x�W��ܶ~v��睷eee�WK��[�{      6S��������k� ���p�; �� ��tg)�����i¸="���sb���ߣV����>�     `s�?0n`�9��uW�����c���(۳[ ��P��wvv�gʾ}_�n�(5�v�|I����hg�      l����^��� ��	� ��r���7dw  ca9j�o�~�G�<n��(un���R[��D��{      6T�ˌ��� l����G�Jv �j_��Gs���f�l������W�+J|,�     `��R� ��f2p`C��{#껲; �4��F�'s���C2����[�D�y     h���w�_Ȏ ����8��:; HP�3�߿��ߟ����q��l����g�      ��Q��e7 �\%; �f[�t>Q�~v �9j�k��+KKf����//%^��     ��������av ��w 6V)o�N  6�M��l~���Q���;      NW��f�v 6��; �}���#�� ��ĭ�V�7�폮��{iD\��     pF�:|Kv �f���*���wew  j�j���t���C�Y����_XK\��     �5ꇶ..��� ����p%��� ��9Z�������C&Aٵk0��raD�bv     �)�- 6��; ���҈ �ċ�o�Θ$����uԺ0"�e�      �����9�ώ ������7g7  뭼y�׻4�b�߳owD���     ��U�\Rv�dw �|� l�و�F�rv �^��v��O�\����     `2��[� �� l�������  ��0"^P��c�!���|�JD?�     �Տ�/.ޖ]�t0p`Ӕ�o�n  �C}�\�svE�Ç����rv     �c���� �G� `zԈ2�,|%"��n �l�=�~Nٳ��&Y�,\�<�     ��ߎ��v_ 6���4%���dw  kWk�e���7j�E�rv     �Õˌ��L� l�A�["b�� �A���-vߞ��D[�ݯDԋ�;      ��7e' 0]��T�z�n��&� 8u���*5���VKyUD�dw      ����s���+ �.� l��f'  �춹~���M����F�K�;      �Z���Mg����k���gw  '�Fyy�ew4�h8�����     ��Օ+�# �>� l��gω��2� 8i{��]x�	�,�+"ޝ�     P�~�8�����1p E��wd7  '�F\Z�*�iJm�5�     ���� �S� `:Ո��N�[�l�n �(�s����gwL��Z�,�;�[     ��u�}��9���#�! L'���DK�� ����q��*�Q�wfw      S�}�� d1p O���� �q��,;a*�Zo�N      ��(�M i�H3��~:"���  Um��^�1���ٷ;��     �8<��dG 0��HU�x� �V���ݻ�]1��G�     �)T��e��� ���; �j+�$� xT�gL�a�     l�2tX! ��H����JDٕ� <\�֙�ÏDD��      �G����ӽ1���f�@�R�'`�ԹV�Xv�4+KK"��;     ��1��1�� `���nvv�1��  �����ݛAܒ      L�0�HW��]�'��x�=;����      l���z��eG ��; c��'�  x�bX=F�     �&���n �w ��j�ueD�� ��F��c�      ��D}ov D�0&�u������ �kJ��Jv�Z���      L���~�s� a��)Q<	 c�����"J�,"�gw      W�=%�fg @��; cd؊�d7  _3j��n�|/     �Ub�PB Ɔ�; ccK�����;� ����9���7�      �����gG ���0Vj-��qp�S�Ǉ�     ����J�0� �����RJ5p�|5<���Uw     `ôZ�+� ��+s������ �r%.�`&;��+��     ������>; ����S��� `�<����J�3�     ��*W�={NdW �C�0vʨ��� �v'VW���E5p     6F-�F��c��ؙ]������ �f���	���I�     @#-�-/_� �����S"F%�� �fefƨz|x�      Xw5���С�; �[�0���; ��;���g��="��     @�Z>��  �����47^�� 0�Z��n buf��     ��^��  �����T����?�� �iU��B-�9�     @��[�fW �#1p`l��Wg7 ����	�     `�k� ���0�F�w �R��5�dgL�Z�oe7      �S��0��[�K�o��}� 0����}��gGL��*�0�     h�g�m�1; ��; c�~(�  �Ui�~ �a�:��fw      �R"�/wܱ�� �����Vk�+�  I)�e7L�R�     �uWK\��  �����6�|��1�� �iTk���sc�Q      �n�:smv <C �Z9|�HD�Tv L��;����iT�������     @�ܾei�]� �X�{��k� `j�яg'L��O�pD���     4L��� ���0�jˇ+ H�S5b6;bڴJ<?�     h�2j9d��g���k�z���~v L�s��w���iRw�<�Fa�a�    IDAT���     �q���ԏgG ��1p`안ZK\�� �j�r��f�F�!"�;     �f�Qn,���� x<� L�Z?��  ӫ��z�y۳+�A�(�fw      �Ӫ��� 8� L��p��� �b[Vګ��1V:�7�     h��
�0��[���{�; `Z��?W;��fw4])�f7      �t��}��� 8� L��N �)��ՈgG4�`ǹ?5�'�     h��e׮Av �w &�We@��%u�γ�;��F�ZF�+�     h�V�n�n ��e����z}v L�����#�h������     @3U�
0AJv  ������q^v L�Q���z���C��>�igV�_�����     4��~��� '�	� LO@�V���1�����¸     � �ƍ�� Lw &K�� ������?��+�(J���     ��Z�ސ�  ������Z��`��;+��wggL�z�yO�Z�>�     ��[ &�_�0Q������]� @�G���Yg=);dՈ��������     ���o/��lv �
w &O-�,�������eGL����/�Q�]v     �l5��1�� �Sa���yv �?������I2ر����Wfw      �תac��1p`��Z?��  <T}�r���+&��9�>����"b.�     �3����S� �TՈ2�,����[ �o�������k�C�ձ����_;%���     `*ۃ�����f� ��p�; �D��/�; �oҮe���;.�Gu���gk\��     ����q; �����Ԋ�)� x�3������}�!���s��Z3�Eĳ�[     ����  Xw &�a 0��RK���;v�Xv�8Xޱ����ѧ"�;�[     �)Sm+ �L� L��'n��Qv ���K��������L+;w��RZ���e�      �g4Sn�n ��0p`"�Ç�D�۲; �G5�^�����z���Ͷ���L�����     `*�;��ޑ ka��$�*- o�D}�`q��O��gd�l��s�֕N���ؚ�     L��Q�; `-��d� 0��o�o^^Xx^v�FZޱ����ED���     `��Jܔ�  ke��Ī��c 09�\j\��Y���N����Tw�ܺ����Ki}6j<7�      �+� �V5�:�Fę�- �)y�D�?������q����V�^Q���     �WF���,����p�; �DԈؕ� ��'Ԩ�=�,|fu����+߹�Y�@+����    ��R�d��$3p`��(��n  ���Z��+��[V^P#f���J��]���Q�%⇳{      �ԛ� �t�0�F� 0��#j\2�tnY�t�s=�'e=T�����N�GV:�(7׈�ED��     x$%���� L��N�9%�m� ��:Q">0�z���ה]��۟�w�����?F�9      ����?kw�7dw �Z�0�jDk�Y�?"��� ���������l�#Oؿ��a�z�3��|����*���Eĳ7�^      ����g�={����2p`�t>ߛ� l�ۣ�Ǣ�/���Wk����}%���E���g���Zf�Q�5�/J\3�     ��J�5�띟� �c6;  N_�9���txv�xvD�3�Ġ�p|%⎈��Z��R�h��/j<%ΈZ�X�<�~�/gEķ"�����j��o     �J�g� �t�� ��Z��T�7�D�����-�v�;     ��Ů� 8]��  X�>       �bC��3p`��<swD,gw        d���0���xe��bv       @��+,ew ��2p�!�b       �^��	 ���f���	        iJ�N �� 4B)���        iF�v�F�� ��0h�vώjv    0�f?���'<1;cz:�?��f�  ��+e�;� �C� ����Y�jD<%�    �\�/�q��S��yg�waԥ��  �d�v�3J�,; NW+;  ��m�     ��r��1�+��sNv
  L����h
w �z�    �2r ��S"���  �����(Ň5    �	e�  k7r(  b�@c�Q��    `�� �ڔ�P@ ������F�F    �pF�  �#w �������u#���     N��;  ��Q{4�Rv �w ���      N��;  ��{��҃� �^�hw    ��0r ��WG��v ���F)%��n     `�� �c+��Jv �'w eT��     �/#w  x�8�F1p�Q��;    @#� �#k��V�F1p�Q���^�    �PF�  �p��� 4��; �R>��;     �F�  �M��O~��� XO� 4�'�    ��  �aOٽ{%; ֓�; �S�    ���  "jT	 ���Ʃ�ܙ�     ��3r `ڕh��8�� ��j�%;    �j�E���+�Ny�3"�������������/�8pp]�  c�T� �8� 4Ni�;�fW     �l����#;c��>7f/g�S����}ֳb�����.������ �q6��	� 4N+;  �[{u���     ��zk������u�v9���y�Q�9gݯ  �g��n ��f�@�,-����     <��;  ������� `���8%�FD7�    �Gf�  ��r��� Xo� 4�'�    Ƙ�;  �6� ����ڟ     �c3r ���� 4��; �T�xJ    `� ��'��P� 4R�2    ��0r �SW�m �d�@#�yJ    `�� ��E1p���h���p    L#w  8y�(� 4��; �4g�    0��� �䬎V��@#��H��?��;     8uF�  �ꖧ>�� ���+�d     �6F�  ��-�w�dG �F0p����;    �����?�G�����������x����  ��J�D �X� 4��;    ����|>V�w�Ɯ���gE9�����  �����ޝ��Q�y~�����8�	
�#��h�O���(a�M��OQt$�(�
�H�	�� 2���8"�BP6���	T���q�k�Tw�r��奞������C���iw ���; �+e�    ��~�(&�ܖ�{��G @�%� ���; }+��    �E[K�  �s2��[
� ���%O�     �H[J��
w  zOf�; }L�����6�    �����D���  �J�w ���; }+5lp    �Ks�U7�,��  �yU{ ���; }k�s�<�    `�R�;  ,����� �-w ��#�4"�f    ��Sp �o6�; ���; }+�("��s     ��� �E+��X� �]��s��u'     ��)� �s�e���\�! �]��w
�     ,��  �] ���; }.yR    ��� �{t! �k
� �;O�     X<� �=� �5w ��'u       @�Ȓ. �M����<�    `Ilp �Ǥ�. �M����h�ug     ��)� �cRJ� �5w ��'u     ,��;  =��'��  ��@_KY6��     t1w  zL�rn� ����kMw     �D� �^�@�Sp���V�]�     ,��;  =&��. }M����ܵ    �)� �[Y�@_Sp�������    X<�v  zMf�; �-�;  �ӈ���=_w     �U�p�f�ZkE��J�1:���#=�@�)�.Wz5{ ���; ���~�    �X
� ]+�l|䧟1bD�Q:�O�b��n���$@+��w �Z��  �V?<?"ʺc     Х���@��#"F����3#�tӺ� ]ld�3ug �vRp��e)"��;      �t�ܾ��;�bR�_w h���  �"bt�!     �B6�t��/�/�Bɽ��G��n�;�4|xd����؈Q�#VZ)���{䈈|XĘ��uw�"�>����̋��ܡ�?�HO?��EQ��Cg<����# @;)���RĳY�!     �NRp�^��ȶ�.b� �����Q~�{�5�~���w�䞭�nd��6�׾6�ш��H���"�����6�8[�'����+׌Xu���X#bܸ�{�H�=���{4��G#=�x��n����U�Vf�b ����^ 0����     ������e��m�h~�3+�Tw��k�|s�94ҽ���s��hL��V��z�E1gN�;fFy޹�~u[�	Y���4�'Gc��#�pÈ#"����}��x\�_���m�ܾRroL��/�ȯc��E��^s�Ԑ�ÆE�c���G��j��jd����G�#�����]t  �{�� @����     �Ej���>����gG�������F~�5�x�uG錱c#��������rˡm���O������m��g̈|���fú��׆�Ɓư��$�Gٛ�1fLD�}����"���h�O�I�F��E�Pr�6ݴ�$m��g�h~���go|c�ӯ�l�;�l�e��UWF��C;Wn_�aâ���F�C�Nс ��)�0ܽ    ��E�	�"�t�ȿwmd[l^w����o~3�'�8T�W��2T^�ۗ��l�M#���h��g"F��P8'{��#�������|#J��c���c#�l��A��K�OK�	�y�1/�}���f�_�&�t&X�l��鑽�uuG�[Y�#��9@OJ�t  �{
� w/    �h�Vp��h~X��=?�5֨;MWiL�1�gt_Ѱ
��ox��=>ϣ��~�Ϙ�F�7�6fL4����"[����1y�PɽO(�/�>+�g�ͯ|y�o�;6��΍쵯mo�5rd4���h~��+�\w��j�_4?�ɺc�����{
�  w/    �eYw��d�|e�]���h�U�d���WD���s�<�����e�.�p�ȯ�<��7nC*�$?�;ј<y���7v�=[nنT��ܾ�����˿D���]4fL4�߿=�*��3��Zw�����A�G��e�\� ����; ,N���#     Х�d�{���=���&����ͣ����S#ƍ�;M%�M����g�F)��`�?�k�]I��(���>*�/�쟗��*:�ϯ�1h���C C�      \�V�	VL�G�������)�-��)�Mo�;
���p�=[o���V�;�_���}.�'�1fL�i  ���;      0�z������_ta4;,"��ӓ�W�2�K.��>{��r{����ht͖�l��#�~U4�ޫ�(  }E�      L�VDJu�X.٦�F~���6٤�(�o��h~���<��c�N}K��M�䞽��uG���;G~�Ց��5uGY~�VDY֝ �(�      ����7���������W�;M_il��ȯ�2�6�;
���6��{���GG��_��W�1jT}9*���g#�}��  �@�      L�Vp;6��};�XDïz�![�ȯ�2�n[w���2`%����g���WDc��r~�Z_:>ʩ�� `���      0����K-�h�ȯ�6[mUw��7fL4�uJ4�:ʍ����;l�J�٫_�lv��ƶ�D~������)�h}�(O<��$  ���8      0�zd�{c�"����^�V�QG�E�#?묈q��N=I��&�Rr1"�����Yy���L4�����c;sf�̟������NIu �v��       P�n/�gY4?�h|䠺��l��#���h}h�H��}�q�gd�o�ԩ������7��w��tn���l̓�Xu�ꆎ��gD���H?�ius�L��#͞��CV_=�SN��mom�9m�~8�-��t�-���6ҽ��	 �E)�      ����F4��}��$/[w�ȯ�<��{D��/�]/�l|[��匫�u�O>Y�ܺ��(�K/���'F6~|u�G�����������v�_1}F��go|c4O�vd�xE�ΨTJ��?�oq�o#͜��_Ez���� ,3w      ` ���;¢5�����ј8��$,�ꪑ_8-�=����ם�V[6�E�>�Q�}vu3�ͣ�F�ݣ��OD�����ܳ�lضٍ]v��c#�o�+�("����~u[��o�t��fΌ�7��d  �Pp      S7np6,�'��m��;	oaQt��#�xc�i��es�3�Dq��������ݪՊ�珍��C�<昈F���}��=�`���y4?��ht`���W�i��H��:үo���n�x�ٺ� ���; �/�,"�;     ݦ�
�#GF>ujd���7GQDz챈G�x�HO=�ԓO?�ɧ"��7T��;/�x>��s#,z[Q��iV+�q���W��GD�5T�;6bĈ�F��Xi��a�"V�ؕ#ƭ��ʑ�<.b�q��E��C����>�F�����]����CE�C�G���f��r��O=ͯ|%"���ӧ�ܳu�ڰ��s�|�ꑟzjd�lRͼ�U�n�5�O~�O��?��ӟ��D�Q� ��)���R6��;     �AQԝ�/ƌ���3#{��k�P^ye�_�b���H���驧���e6rd4v�)���T=e�#"?}j�8 ʫ�����eڱ�==�@�&N�tｕ��%�EGzxN�SO�3������=�#[w�H3g������N���� �r*�(O:)Z�uJ�ܹ��T�R Н*z=# �bY��;     ]�U֝`�ر�������G��#���CeҊ��{��(�9'�wo�'?�'ða�<�h�C=�C��6��W[n�=;Z;�`����(���"����F�L���ͬY��W���Ƅ#��Z������S��t�r;KC����� ��    ����+���߉�-o���4kV��.��~���WD���(&N���G׳�?ϣ�����Ν?�@��f՗��+�'Dz��f��t�QL���#�5*�3Ϩ�C*����m�ͣ���'V�}��ʫ��b��D���k�@��t  �{
� ��,bd�     �B�{���F~�E���M�_�~[oi��ZίDJQ�65��w���Ý?�ٌ��_��?����F�f�#�:��r��~��w����ҝC���3����GG~��}��=[��p�U"?��ht`���ł�:��h�OēO֗����{
� ��d�;     ��?�w���F>��6ڨ�g?�L�>8ZGY��B�?���[F��:x��/~!{������f������Ѫ�F��fώb��s*��~֙=_r�^��e��5F>czd�zW-�4��(��:�Ӧ֖��6,E�u� �vRp`(�    ���ϯ�܅��׼��G��o��=[Gyɥ?��<�ɓ���/FEg�βh~�?mr��e�oV}����֎"=�@e3�Q���(v�5�駫:jT�g����^����]7���������WD��W�1Ւ��Ŷ�F���2�V[M����� Yw      �O�c{y���򢋣�~�H����;�,���7�>������Yf�;}-�l|�S�VZn��s����H��_��>��#�=��X�����GG~�ٽ��}Ԩ�^��\�ͣ����1fL�s-��Gk�����OF<�l=�ͦ�; }M�����_D�y    ��t��>vl��=�������־�F�c���\�t�Ql��H�_�كnr�4���B�e���|s{<�|�/��W7s ���Y�>�����n�Q��uf��_����H0��    IDAT�ꪑ��ht`D�u&��I?�q��2�k���|�ϳ���; }M���V��    �h�,{7������6ڨsgFD�����߷�r��=�+<�x����~>�(:wn�E�K�E6~|�΄6�6߬�r{J�:��H7�X��R^uU���R��Q�"?�����j�v@��z���9�k�����`���R�_�F������@_jd�. }M���6��]w     *����fγ�V3g)d��G��wu�H)ʓO�������;�ۤ�)�t�������;w�I��G>uj����(O:9�K/�t�)O9%�+��v��ё�}V�ȑ��m��U�Z��v���#[s�'z��y��o�hw\D�UO�V�Ҙ�3 @;)������ug     �:�;���������٨.�|ꩡ���N����.������=������cQX�1c*/����/}�ҙ��uđ�ڡ�GGV��6��^�o�0bD4�?>�'�X۟�鮻����QN�^����,�^Rw h'w �Z�QxR    �'���#?�̈��⩃�NI��m[o�����}�|2��'Gk��t�&����V�g���~�a�+������kG~���u���W\�{���k�@�+��s
� ���'u     }����"?���ͲU�B`y�eQl�C�{�;J�J)ʓN�b�]"y��40p�O&b�ܺc��4kV�>l�1j���ZDD4��*��#�x�z�E��L��F<�L=Y�@Sp��5�    z[�G���G��"����Rp/�h}�3���G"�ϯ;MOH?�I۾7ҭ��;
���+��c���"�xc�1��J����9���q���0gN;M���9���e�@_Sp�����    ���V���s������'��b�ݢ<㌺������QL��7��_YF����NѿR�ַ�Uw��dY4��+"�j9>��7Q��}�n����Le�� �5w �Z��    �'e�xG���"{�;�w�3=��|Μ(vx��n�;I��ӟ��s�(����$�����{���ҏo�x�Ѻc��ˢ�~�H>XwL�Һ3 @;)��ײ,���     ,�,��>{G~�w"V_��G�9s�:����Ŏ"͚Uw����s��o�(/���$з�k�Ww��W>ϝ�jEkʔh���g��;(�L����@_�Rj�o?     ��*�D~����g#������G��.�چ\����!�Dy�u'���~���#���;7Z{��I'ם��R�Qw h'w �\ց߀     ���׿>�gD��ww���zv�{�яE�뮺c��V+ZG�;�N}%����j�P���EQw����'�m����� �B����      Ԫ1aB�^�Zku��t׬����y��ﾺ����t��u����~�È��1�΍��_֝�o��o�b��{ �Pp      �1bD4�||4O�ZĨQ�;7�(O�ڹ� X��GuG(�7��/��9?��&F<�X�Q  ��*      :.[s�h~��������R��>:�s��� �(�(��S��?�Sw���jE��<�亓  w      ���w�;����*�=xa�}��=`@�;���ү~Q�J�
�7/Z98�뮫;	 ��i�       y�����ӕ�@�я�0x�������/��Sn ���;      �v��kG~��8찈F�M�R�>��v�+��#��_����[n��}�E�󮺣  ,w      ���n��3"{�:xYF�ȏGy晝?`��_�Vw���n�u�zVy�Q�41��G� 0��       }bذ�V[-b��E��zd��w�+���ד�(�u�aQ^|I=��y�"{��)�yg�zOJQ~�����	u'  �     �zcW��Uk-�c�Q�/���կ���Ǝ��ǌ1r�߾m��Ϳ:�ٌl���G�1jTĈ�Co�G�1|DĨQ��1lXĸq+�1T�(�u�AQN�^w�����Y���Tk������u��Q^zY�I  x��;      T�1a�hLر��k��h���]Ww�����n�?�I�1`��<Ş{F��ֺ�  �W�     ��1~{����N t�4sf�&��� �ߩ�      ��SOE��.�� �����Wn �R
�      @��H;N��_ԝ �b��E1yr�ܹuG `1�       ��t�=��탑�( @�*�h���Q�uV�I  x
�      @�J��jh룏� �V��Eq�G"��ם ����      ��t�Q���y�� t�t�}��c�Hw�Uw  �R��        ˪��(>��r; �X�[��n;�v ���      ����߈�!�FE�Q �.U^~y'E<�h�Q  XFy�       �JJ����G��o՝ �V�?���ԝ ���      t�矏�!�Fy�eu' �QJQ^|I�>�����;  +@�      �n��G��G���N t�t�]���'#��guG �
�      @�z��(v����;	 �m�"�o��/9���N @E�     ���x Z��i�캣  ]&=�`�&��w��;
  k�       ����6Z��� ,�(� �)w      ���n��;F���   @�)�      ]�<��(v�1wn�Q    �A^w       �h��u�qQ�tr�I    ���;      P���������ں�    P3w      �>s�D1y�H��Vw    ���;      T$�zk�ܹu��i�3Q~�3�z��( tX�㎈矯;��j՝  ���      i}�(����E[o��  ,R��         ��_(�  ���       @ǔ�__w  ��)�       �1����  �b
�        tD�93��w�  �b
�        tD9}F�  �.��       @G���   t9w        �.�sO��w�  �r
�        �]��ں#   =@�       ��+����  @Pp       ���y&��o�;  ��        ,��##{�#[m��g���裑~��矯;K�n�%�(�  � w       �'d[l�	_�X}��y{��(��7b�#5%�Ŕ?���  @�h�        `��,�Yg�C�=""{�["�������gc��}w�	  ���       t���$�sΉ�QGE4_s��X#�K.��ĉ��J=Tw  �G(�      ��,�;A���*�����D��fKw������	�<�?"��XF/}i�	  ���      �C���\Ĉu��K��Gc���ct���u'X�Ƅ#����^��e�����;�ug�z��f������#   =B�      ��d[l�ԩJ����u��t\��C"[��c�E�G󳟍�'���y�馑_=#�׿��p+(ϣ��"��;I�eo[4��c   =@�      ��d�o��^�A.�GD�j�E~��6ؠ�$/}i��'��]ɸ��)��.�Ƅ+��B����W4��޺�Ԧ��O�s  xQ
�       =Hɽ_n_�e/���K#{�[k��m�Q�ӯ���v�ȑ�<��hw\D�W;{i��r���N4�ٺ��D��:��ԧ�  t9w      �6K��}Ă���6�,�o�����[n�駷���m7n\������э����#[k������"�pZ��Vo������_|Qdo[GϭBz��9�T:��מ�m�E�3 ����      �f��ۣ�cψg��|v��o�g�a��2ʶ�<��~+bذ�g���C�|���9?�,�6|x4���h�o5�^L��O*�'�1jTۏ���_#�>=�׿��gEDdo��#�h��f���4cFe��'��8�ڒ{�E~�W"V��  @�Pp      �t�Q�W{J�D��T�-6�|���ln��Q�W[6�/Ny��:���J�F4�9:���lV3sQƎ���3�q��;c�5׌��K���v�=g���/�8�5֨lf���hM�)҃V6�EϜ5+�	"=�puCW_}��'򼺙  @�Pp      �%���[�}�rڴh}���V����}����#V^���ek���G����^*�FE�䓢y�Q���]w���"VZ�����5iRG��>{��h�4�Ғ{��&���Q��  ���;      @���~�����k�}���ˣu�G+-�g���|����_����_�����\� Y4:0�Ό;���������W��<�������l�2ghCɽ��Gc��*�  �w      �kk�}�%��#+�����ܾP[J����E��w���w�l>n\ɪ�m�E�ӯ�l��Vl���ќzZ4;��`/H��]����Z���2{v�&�1��f6���^W�<  ��)�      Ԡ�%�ӧ*��`P��������y�F�����ãy�W�y�q�n6�J��z�_q�r���5ֈ�⋢��V��J��������t�H�fE1aBu��G����gE����  z��;      @M���o�����_�#��(��6��<�h��e����\3�K/�ƤI�ei�UV���s����tY���D~�Ց����I��3Tn��+�[�4{v�v�XY�=[c�h�qzĘ1��  z��;      @����gP���ӦE�#W��="�&�7��E���O���Xi����hst4O>)b��}x・E~х/{Y�1�=�Ȼ�ܾP�=;Z�v���H%�׽.�'}3�٬d  л�      j�����\�}����e�{Dd�~u�W^�ɓ#�lȢ����_pA��V���Nhl�}�W]��_����������y�qÆUzv�=�k7���4kV&T�ɽ�����*�  �.w      �.�֒���5P%w���UN��Ï���c�Dsʱ�_��������W�l�5"{�y���̧#��3;(�p�ȯ�2����G���"�h�h|��1���Gc��*?3�}wv��0�	i��m�U��w�5�?��Y  @o��g�       }faɽe��]�����Ї"�ϯtv7Qn_�rڴ�����G4����6�4�gT:�k�y4;,�������њ8)bΜ��U�4{v�&���i�l�o|�c�y4�3Ψ   �klp      �"m�����F~�9�GW>�(�/Yy���:���V�Q�;UoA�C�5+�	*�����h�O%�  �ޢ�      �e:Rr3���uRn_:��G�##ʲ�(� �}wv��r�B���,���C]�Y  @O��       �?J7��^{G~��#FT:;{�[#?��H7��ҹ�1"�w�6�����?�b�#�{���u)�M����W���ѽx��G����1�#[m���#�N�\ҝwE1iR�#���2i��hM�9�i�"^��
�kqxd�FE�_tc  w      �.�n�!�=�*�W\��6�$�M6�tf�I?�!�}��r�B�ZrO����<ҝw���&D�/�T�=ͼs����uG�\�5+�	�y���Xc��5:0�׾6���x��
  �L�      ���o�bϽ�Rrg��o�b��",�;J��Tɽ,��կE���-r�wy�E�fΌ�O�l��j�l�̙QL���cuGi��7�g[l���Q~�C����OD����S  @��      ���{gB�}��(�ϝ�C��k������D��6��tRd���P�e�f͊b�]��ܾP�5+���+���N4O=��d]�(��s�H��~�I  �6]��      ������>[w��6H����iӢu��܌^�4sf[m����?{��(v�=�o|3"���[�;����s�;JǤY���0!����7�y���Fd�|e�I  �6
�       =Bɽ��ܾP7�����G���#�{߲]�jE�_���D̟ߞp�!���QL����uG�4{v�&�<P��2n�Ы*  ��Rp      �!J��1�������R�'��{F̝��cʫ��b��#ݷ��6H��Ť��ܾ�M��&{�;�����  j��      �c�ܫ�������Ϗ�~�EkʔJ2�;�b�m#�tS�3�r���ٳ���D%���8��ѣ�  ��      Ѓ�ܫ�����*����b�	QN�Q��'��b�ݢ<��j�.�?�۟x��gw+%������<���c  @�)�      �(%��ܾx�.����<����t�m�9�(�5eJ�>�ю}��o~�ܾi��hM�9b�#uG�z����/�;  t��;      @Sr_>��/��6-ZG���{y�9QL�)����ˋ/*����t�mQL��ܾi֬(&L���Ō��u�  ��Rp      �qJ��F�}�\о�{QD�GE���(���/F��ϣ�f�H��u{����(v�%⩧�2���ٳ���D%w  �o(�      �%���ܾ��.���GT[r�(v�-ʳϮn�2H�C���EW;�W�E��n���@�  �{
�       }B�}ɔۗ_9mZe%�4s����n� �
X� Z��)S���n�9��#�|��p�E�  �k
�      ����_-������{+L�G�}є�W\%�t��Q���H��Wa��R�'���="��]�1?��(>���y��6`���њ�s�#����̝۷�~�n�-"�忾�d  hw      xA�##{l��K7��v�G<�TR��Sr�[���Y���"�{�P��]���?�U~��e��?���x�6$,i֬(v����WZS��\�n��wD넯.��E�)S���� @WPp     ��������?�.h��<唡2ޜ9��H�}�r{��iӆnZڒ��y��o�hM��B���-�sO�������놾����*�Y���qB���;J��SO�����V�W��E-�����G1qR�'���T  �M�      �J���E��N�?���ͼ3��w��~>�(:��͠�ܕ�ۧ����*��ٳ�x����>�C�V�OD�ݣ��7"RZ�C��ӣ��#�{�C�G�=;Z�v�M�)Ey�	�����N�~)E�C���iK~\YFy�yQ�{�H?�Yg� P���  �Nϯ��+R����    ��l�5��OGc��#ƎzcQD���(O�v��]��N��Ə���'FVw��)��h��q�5&M�族�h��~���k�u�s�֐l�5��*��)b�U��}�9�F�S��h�jH68�W�:�g��*���1�駣<�(/���(��v�hqxd���Co�7/�3�<�Hw�Uo@�.�;��K�! �]��k
�    @%ƍ�h6#�x�E7��Ǝ��GD��Z)E�5+��^婧�����������l��#,��I'Gy�	u'���lF��҈��"�����@�Rp��)����     :#[s�Hs�����5v�P�֫w P?w �Z^w        ���?����կ�}  �.Ө;            D(�          �%�          �

�           tw           ���;           ]A�          ����          @WPp          �+(�          ��          �

�           tw           ���;           ]A�          ����          @WPp          �+(�          ��          �

�           tw           ���;           ]A�          ����          @WPp          �+�u     �3'"�ϤȞiDz*E67""�4��l\iLD4�ġ    IDAT�����՘     z��;     ,�3)��"K�dwF��9,���~��'�eHZk��<_�DJ��#eo�"�[D�nSn     �Y
�     0�Y�8K�q}���ܜ�~�s+:4��'"�g/�'""��/����ٻۘ������߹�s]����8�9N0-2�e4�Ӯ(@ԭe+E�`t��:�Vt�Tc7E�Z��A��Ҕ@"5��MQ�
���5M��BӐ�!�ulb�I�:7��@�4ʍ�|����|���O�y��R���F��E���~     ̻�=  Φ�`��5�-�;   ����Ԉ_��'�:�`Ƃc�]6�O�uQ��qU�   `nܵ6�ܟ= �'�    ���G�ǣčk���=�%?<��"��`�7#ʏEĻ#b[�2     8�z�     �z"����J�k����mn���ϴ6}im���~7��F�PD�y�&     8W�     ,�'k��WW._�~�['�7�:�������{��kć#���M     p�	�    Xh5�f�쯯��\y衣�{NU9p���h��NK������=     p6	�    XH%�@-q��h�-�z0{��ڱ�y�p�.�?����     �� p    `}|u6}����x�m4��?�^5n��     g��    �Er<jy��h�����c�cΖr�𱵃����w    �|�     ,��kԫ��1{ȹ���yS�f�Q���     g��    �E�����_���r��:���d��5�粷     ���    0�J�O����9�X��,�G�X{��o��_��     �c5{      ��_\�~�Dt�C��{�׈wN6�G��?��     /��    �O%nXm�W������������-{     �w     �P�������+Z��~*jܔ�     N��    �y�;�����۟[�����?V�~6{     �
�;     ���������������y�dm2�."���     'K�    �����t��r���!�<����?G��     ���    0j�������!�f�h�P�G"�fo    �"p    �}%nX?x���3�ն��ֈ��;     ���    hݗ�\����cۿ����w     ���    в�����{��C�]������#�fo    ��"p    �]5n�on~1{Ƣ�F�E�'�w     �s�    ЪG�������_����     �l�     4��l���gX��|4����     �l�     �����Of�XT���#��     �Lw     �S�ʝwN�g,�r睓��d�     �g�    Д�P��Od�Xt����Q#f�     ���    Д^�Gʁǳw,����'zQn��     O'p    �%��R>�=bY���ƈ���     O�    ЌR�7����;�E9p�H����     ��;     ͘�zs��e��p�    h��    �V<��җ:M�[���[#©�     4A�    @+~��s�8{Ĳ��5����     w     Qk���˪�    �6�    hA�V������f��GD��     w     Z��2}#{Ĳ*�=wg�      �;     �j���ް�J�     ��    ���dOXv5��     @�    @�:���	K��{�'     ��    �l��m�����"�]�     ���    �l�<�=bٕ�G���;     Xnw     R����o�Q�     R	�    HU�ތ�C�     Xnw     R�R����T�    �\w     R��U7��     d�    �JT�     �M�    @�*poEu/     H&p     W���	|K���	     ,7�;     �j}I���ە�     ��&p     UU7���^     �J�    @�NT݌��     ��    �����Q��     ��    ��e��K�     ��     dۗ=�����     ,7�;     Ɋ��5�D�+�w     ���     d�U/�{i��ew|8F���     ,7�;     �+S��'�G�     ��    ����2{��     @�    @�R���]W�M�     @�    @���5b%{ǲ��%�5�;     @�    @.�ll\�=bYM�ë#�y�;     @�    @J)�foXV��    �&�    hB����˪�µ    �	w     Z�O���G,��ᾨ��;      B�    @CJ-��ްlJĻ�7     �S�     4�D}W�(�;�E�(����     �"p    �%{�{��!{Ĳ���F�Wd�     ���    hJW��doX���7     ��	�    hJ�����eWg�Xt�={�+"�N�     x:�;     �)�9Y�,+]�`�     x&�;     ͩ%޶���ײw,��={^[#ޒ�     �I�    @�zQ�G�G,����Q�g     �3	�    hR��}[{ޖ�c�l�(Q�?{     <�;     �*�~�^|�����^tѮ^����     ���    ��]6�����b�_�P�f�     ��"p    �i%�OO��g�w��ˮ�?��     ���    �֭F�[�`pQ��yU/���(�/E�J�     x>w     �W#��K��F��-�F�ƽ��5b��     ^��    ��Pj�y:�?{Ǽ�n�D���     p2�     ̍�?l��0{Ǽ��QK|8{     �,�;     �Wj�<�n���M��7�(��     0G|�    ��Y�Q~m���?{H���]]k�FD�go    �S!p    `����֞=��Қ�pxe��3�+{     �*�;     �jw���M6.�&{H+&��yC��BD\��     ^�;     ��Z��m�?�=$��`��W;"���     /��    �y�^j���`���!Yƃ=?Y��zDl��     �C�    �"X�(�}2�zݻ���1�J��]���zCD�d�    ��%p    `a�o��'_��󷲷�m������]��-     p��    X4{��_�������s��������D��#��{     �L�    ����(�ir��ݓ��{�ǜ)��ˮ�:tW�����     �4�;     ��U5����O�K.ٝ=�Ū/��x8����Q��=     p��f    ��9�wo|�ߚ=�9_�Z��S�Ξ�)Q���j�����ӈ���<�=�d�K.�=^]}�d2���ؑ�     �6�;   ���W���]�3���C
DD�z�x�jď���_�"�������G=��^�w��{�$�{JĶ�=     p��    X6kQ��"~x<~1j��?9qK��7�U���>���G��K�����    XB�    `Y�"�uQ��&k�o?��ů�lm�޹������m�z�\7���J�K���    @��     �3J\�ո�[[���;j���"~wu}����ř���w����ꮔ7��N"��E�F=;     �?�;     �U��=���Ԉ59����p��7j����]-ktO���D��VV����f�^��Y�;K�v��Ԉ}Qʾ����x�;�D�    ���    ��5vG�7�Q�F��FD�E��V�^zQkD/JDԨQ���v     8)��           !p          �w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	��    8sݶ-Ff�h�t:͞       ��;   �y�ߏ�G�f�hN��E�      0��          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4a5{  �����j��5�ϞA��~8�����=        x�; �t�\[�+~�G�g�쫟�L��        ���            Np   X(;f�عsg���w�D� 8�f���_|q���>~<^����3    ���   ��'���_~y���x { �SO����G?�=�d����kn�9{    ��^�            ��          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          Є��   0��O����f�����3�3;~<��'�����      �  �I��J/�����++�S��}��7ޘ��M;vd/���6��O&񊚽     �=��   0��5�N�o�Ǳ�*8u��͢7ފ?�]�     �f	�  ��Q��6ފ}3q" 'g="�O&񿧓����      ���   N�����l�'��g��i�w]�lk+n�f��(     �&p  �aZk���bc<�a'Y��E�U�i��d�S�     N��   N�}����8��N�d��	�t]�bk�Ϧ1�     0g�   p�ND��i�O�e�)� ���i����v     �c5{    ,�?���p�����VV�� p]Pk&���*l `�}�g�k/ّ=�D��7�s�/g�   ��   Π#Q��t�9����~/%{ g�k�.�N�.o�  `I���s׮�$z�ǲ'   ��=    ���m��7s�/���WM&��8�     �w   8KF�Wf��?�x���������㸽���     ����:   �E�Z�:�}�����<k0�Vj�+���_�,��c      �_�  ���v1����4J� ^�Kk��'�M�     p�8� X:+ǎ�;�g� �ۻ.���=X2'"���4����H5��;���r:���Y�5{
     �B� ˧�8t�p�
�m��q���3�%��unM���c*rh�t:�?��      KA�   	��G�����z� ^�K�͞      �4�      �L��я},{ɮ8�-�    ��;     ��)�Y�z�oe� ���wD�~�    8%��           !p          �w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           ���=        ���ɽ��c{���ײ'   L�       ������h�e� ������.|Y�  `A��           @��          �F�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&����w7=v�w���}��x2v\�Nl�q��*8}�(bK� � �-kĂv���G���] �HTm�� TK	I�3��9s����*iK�p�\���?�7��"���|��          A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A���6    IDAT          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ¼�  ��V�����?�z�=�����3        �� p &�?>���?m=�ƾ��/E��[�         ~B�z            D�          �y�      lV�|��w�z�}�o���z    </�     dSJ�@	�    0>^p  �3�E�+�Ǳ<؏\.���/t4�ū{{��Λ!      �$p  �3pi��������i�9 <��}ߺ?�=x�������ͽ�X�     ���   ��\��������A|�k� �wRk���q��q\������n=}1~�X��     ���   6��2vޏ;<�7��� ����:�88�88�W��慽���^ͺ��      FM�   p��㥃��{�ժ� ��7W'���9�������������]_�      xw   xL]D|��(N�⟏��U�0eǵ�W��"����lw�z*޽x!�Y,ZO     �;   <����x�� �������u�9 н�:���G�����ĥ���ޅ�X��z     ��	�  �!�j���?�?�Y.�[� <�>"�u��X.����Wvw��ⅈ��5     ��-
   <�?Z�q2?�ܥ�S~lu�||��?�zF3���/D���3 �/��m=��,�����ϛ���qS
     �g�  �C�+%�Ji=��Xv]�vvZ�h�ٮ���Hf��3�?W�Z�Ο$      C�7           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           �0o=    x<��899i=Hd�Z��l�zƙ��U�	  0J����Fw~������7���   )�;   ���|�~���3��.��o=R��{�b=������ `�~�7#.\��z}�_�  [ӵ            w           B�          � �          �y�  gmo���~�g�����n�	        �����[��w��K�g         �]�           �w     �t��u�׷��z������    ��	�     ��[��w��OZ�     xd]�           !p          ` �           ��          �A�          0w           A�          � �          �;           � p          `�           ¼�    ����>._��zF3��� �+�<�٬��3�X�[O      ��   0R��:�^��zF3wؼ�}6����g������      ����            ��          0w           A�          � �          �;           � p          `�           ��          �A��[�e�	        t�z  l����j)Zo        ؔZC@jw r�ա       H�x���� �VJ}��       ���� ��[ �m��<��z     @���ƺ���AC7��� &��; �	�ȭ��p     ؘ����� ����; �u� �6��9�       ix���� ��uu       @� ;�; ��u�^�        �2�� �	�H���u       @����7 �6	�Hmg��       i�R�[o �m��[���        �)}���  �$p �w��       i�#�Zo �m��Z�XG�I�        ���l�? R�0n.       9��: R��^�ps       �`]�|s�z lӼ�  ضR�(j�  �7[�������fJ��<شW���X��i=���O�   ���z; �� `�N�_�Z�x��       �'���{?��z lS�z  ���      �[ �m�0w       @� =�; ��Z�       ��G� HO�@z]q�       2�� �	�H��       @�� L���)�       ��E=n� �M�@~����        ��J�ZO �m��_�       �Wkh  HO�@~���       ���� �; �U/�       x��	��_�;       ����� �W��       d��  ?�; �u�:�       	x���� �W��       0~�b��ȯ��       �_�@ 0w ҫ���       @^p`� �Wz��      ��+w ���_��       ���J�@ �������       dP���� �W}�       H�� L����j�n/       �W����ȯvw       @��HO�         cPJm= �M�@~]-�'        <���  ?�; S�p       d��  =�; ����       ����� L��       �@��  =�; S�p       d��  =�; ��2       �@��������w       @U�@z�? �+w       @�����v ���<       ����� L��       0~�W��O�@~��y       d p =� S�p       d��  =�; S�p       $�i  HO��8�       )h  HO�@~��;        �Z� �'�`�       �4 �'p ���       H@����;         �	�ȯV�;       `�j����v �W�E�	        O��n�z l����J�ϵ�        ��4 �'p �R�       ��+Q|���� ��W�;        ��? ���_�w       `����������       �Jh  HO�@z%z�;       `�J��= �	����       @�� �'p �"p       Ư���� �W��       0z}�E� �mw ��y.        � ���^���z       ��+�[/ �m��^��T�        O��m�  �M��8�       h  HO���;        ��W�HO���      �ѫ�k  HO��T��      ��+�b����;        ������	p{       HaQ#�G �6	���*p       r�|Y@jw R�ѭ�E�        1�	�HM�@nn-       ���T� �Mw rsk       H�������Ԏ#�Zo        ؔRw R��Z�X\l�       `SJ�k! HM�@j]�P       䱮U@jw r��C       �F�B ������έe        ���  9�; ���       �B �����jy��       �M��HM�@j��:        �R� �&p ����       $��  9�; ��Z�       �D� �&p ��P       �QKh! HM�@j%|�       ȣT�; �	�H��C       ��ӭ �6	���R�        �\� �Mw �s�       2�B ������       �L.�;wε �"p �1���w        lԻ�>�z l�����]{6"J�        ����|���� ���:�9        ��M i	�H��p�       �)kM y	�H���V       ��K��  -�; i�e�0       �S|���� �U��      �|4 d&p �һ�       �S�&��� �ջ�       ���  /�; i�p[       ȧD\j� �E�@Z%��        6�F}�� ��; i��9        #��������       @F� ������       @F��;wε � p �z��ND\l�       `J|�� ��; )�       ���z��  %�; )�k��z       ��t}��  %�; )�:sK       H���F �������q       @Z%:m )	�H�tw        �Z� �$p ��3\       @bE@Rw R*�\i�       `[J'p '�; )��˭7        lK���? R��R-�Z�        [�B� �w R*5^l�       `���  � p ��U��      ��v�[϶ �&p ��o]��y�        �tr||�� �4�; �'o       @z]�i$ HG�@:])/��        �m��; ��H���       ��J�H ����tJ��       ��j��r@:w ҩ�8�       �y���� �SJ8�       �U� 		�H����       �$h$ HG�@:5��       0�jDi= 6I�@*5bV"���       p�ŵkj= 6I�@*�/�t5"f�w        �����{ R��ʢ�o��        pVf�j% HE�@*�֗[o        8+�V�d� ��Ew��       ��R������Tj��       LG�z�� �$�; ��w       `J� �"p �R��       LG�����d��n       �Q"^��n�o� 6E�@�ƍKq��       �3T���7Z� �M��ƪ�}r       ��Y��	 ���F�pX       &��z�� ��; i��	�      �ɩ��  �; ���       0=E3@"w �(]8�       S��  �; i�Z�       �	*� ����H���        �^�Y��9�z l����/<϶�       ��ly����# `� �p:��n�       ��y)�	 R��B��!       ��^;@w R�n!       ��k' HA�@
�!       �0������C       0]��v�� �P�       �I�p�{w�z <)�; �W�_�PD\j�       ����^n= �����[���v       `�f��P 0zw F�:�       D-�����0z��       @D)
 FO���U�3       ��54 �����s8       ��� �I	���c�        �+����# �I���7�G�s�w        ��d�w FM���-���[o        ����q�0j��;�7        F-w FM���u�j�	        C�E�0jw ƭ��       ~�
�9�; c�w       �+�w�.Z� ��%p`���/��Z�        ��ɽ{�[� ��%p`�NOO}R       ��4 ����Ѫ��i�       `h��
�-�; �U뫭'        M�!p`�� �Wq�       �g�T 0Zw F�8�       ���Ոy� �8� �R�r�jD\n�       `�v�ׯ��z <�; �t�X��z       �P��|�� xw Ʃ��[O        ���� �q���       ���x  �$p`�:�0       ����x  #UZ �GUo��]�������       0T������j� ���U��C�       ��:��?�z <*�; 㳮���        0|�����0F�j=        `�jT� �#p`|J�]       ��i, �; �R#f���;        F�#���/� �B�������G#��;        F�;],>�z <
�; �Rf>�       �j���Q�06�j=        `D� ����Q)Q�*       xh���Q�06�l=        `<�k���E� �� ���՛�D��w        ����޽O� K��h�Y�k�7        �N)� FC��h��?�z       �蔢� `4� �Gu�       ����\ 0��  x�����у��i�       `d�"�r��;�� �/�w F����n��       GYwݯ� C��8��SY        �i��gZo ��!p`j�_���M����S�U=3		Yg��2B��-A�M�[T""�\Xr����Gp?p	�x����9G�	��Qnsk0�$�]=�$��LWU����$$=���Z�?��yU]S]5��~��d       �0���d       ��Q�f�)�� ��}�RD���        �b'��9?; ; o0X���       �iW�Ge7 �=1p`���
       �x�b���3p`�_��        0�J�` 0���h5�Q.��        �_]O=��� �J��h�N�qbv       �h�v�|Dv |%� L�Rʥ�        �b\�%� ��0�j�R       �IJ�/�n ������U#5���       ��QU{��� pw��X�N�qjv       �Y�zQv �w &W)�f'        ̚q-�d7 ��1p`b_�        6])��� �;� L�ѨQ/��        �95.����� �+� pW���i�0CF�o5�q]�r]-�O4">Sk��;�K�L���h�P�'����qm�\�xwD�_������.�      �f���GE���C �K�0����(5��ٝ5�W��|_�ԓ>Z��v�?��z;G���Z�eQ㢈X܌�      �����0p`��  �+�N�j�gdw���%J����?����r�5��x���/��xvD\QOڎ�      �8�x{u�� �R� L�Q���-qzvL���(����=o߮Q�ݩ���X�Ќ����he�       p���ڭSʍ7��/d���Y��R���;`��Q��j�~��t�jv�]9��tv���(/����=       |�2.��. � �P#;  �Tǥ�0�>Y�����<���_5��������7����Z�}5ʫ#���&       �@c|Iv |)w &N)՗'�r��5���~���W��o�5;��*�ݲ�_~Uk}t^D�)"jr       Q�\��  _�d ���a�{KD�����|����Y<t���K6ðӹ�F��xpv      �������'>�� �<'�0QF��Ea��w[�x^��|ɬ��#"Z��_��+��?k�=       s���j]� _����2����0�5�f�핕7���]��JĨ��6�>:"���      �W�(�g7 �2p`���KD�_o�r�w8��씭�����5X� "ޖ�      0�F�d)� �y��3wZ�p��H��hkQ1    IDAT�W�� ;$à�{yD}]D4�[       ��8��;���;  �	2l��~71�n+u��y�GD���o�Q�����-       �Q�g7 ��09j�e��T����VW?�ݒm��{i�'G���-       󢖱� �d @DD�h;݃qzvl����������C&ɠӹ ��YxO  ��D��KĿ�Zo�w֨�n���(u�h�c|J�Ɖ�����~q^D�ʎ   `�i5�iey�Hv �0�ޣb\?��۩F=X�͋w8���I����?���[  `��Q#>؈���h\;*��n,��A5�]ZڻP�y5,�~}�qI��   �/��oX8���� 0p`";��Q^�����(qi{e��C&�p�wy-����n �-T#�J�?��x_ke��J�h�1�v��Z./Qͭz<    �E}C�߿*� ���N�����&��)�~�=�!�`�ӹ�D����n �Mv�F}Km4~k���fEԳ�^ֿ9J���� �   �tk�W� � ����i���iq̋�k���9;c��uz�*Q<�  6A-Q�u�u��Q>{z��t��WE�s�    ��x�y��n�!����L �jyR�3?�hܾq���OD�{�;  �8�k�G�G����h��~h���핕h�W^��܈���8��   ��i4G�g7 ��; �J�O�n��Q�mE}iv�4*�ְ�܈8��  ��m�f����S����g��;������U�a뜈��X�n   `��(O�n �� �|��a�ۏ�3�[`����#�|mv�4v:��Q�,\�	 �t��D}i�ߟ����.�h�r�xdv    [�p+���?���2 �hO��0ng��Ÿ��}n���  p��?�ڵ�0n��h��^�Z]�ڨ�]qkv    [fנ6���|3p Um���� [�^��g��+fEk��+k�jv  ܍�j�\�ZY��r��k�1��D�۫+�6*����    �Fi�gf7 0��HS#JDyzvl�Z���k�f�̊r���?��  _��ﴆ�G,./4;e+�ZYYn�W.�Q^��    6Y������� �/w �{������;`��vky�����������  ��#Q�핕o/���g�c�C�-��_���Dħ�{    �T'�>u�c�# �_� ���[Z1���Ɏ�E%�F#^��  q[��'�WVޔ�a���j_�[    �<����� ��2p M�����bo<���~vĬj//�MD�'� ��U����VW���B����<l6.���f�    �Y��k�Bv ����k�ރ#�����Ǎ��YW�姳  �S%n���׵WV�!;e�p�@��м4"�2�   �Mq��׻8;��d�@�q�������X^�>;cֵ. "�"� ��R"��k��g�/Vn����`����    �_���� �|2p E�����Ju�xmvüG}Mv  s��Q��߿9;d�O~����"�_�[    8>%�3jD�� `������}��xhvl��w���SvżX���U���  `..%���߿.;d��C�nE}\D�n   ��Ոް�{dv ����m��l^�� [��;��D�J)o��  `歗�xfke寳C���~�@�xjDܙ�   ����xfv ����mW����,�F��ˎ�;���N  `��(?�Z=�g�Ӥ����e�    ��M� �w ���^���R"�Un��PvǼi��^Q���  `f]��/�dv�4j��o�o��    �X����zɮ `����>{몒�[�F}Gvü��x� �
�Z��甈��i���'"�9�   �c4�Wd' 0_��f����J������U#�}�  ̞F��\n�i5�c��C��WF�(�   ��+� l+w ��ѳκD\��[���n�!;b^-�ZG�;  ����ZXY���Y�^Y�Ǩ��    �s��#�# �� l��x��Q�;`��f̳r�G�Ƈ�;  ��G��Ȏ�%��ڏ����    �A�Nq`���mju�*f\���N�w�ԫ�  �%�v<xcv�,)����ߟ�   ���Z�]#�� �w �Šӹ "��[��ov¼G|4� ���KK��1���ߋ���    `cJ�=�N�� �w �I����b�U�ǲ#��x�5  `ԟ-�\3̮�U%�'�    ظ��� 惁; [�F4Kĳ�;`�(����y�>��#b�� �T��u�)��1�Z��{#���    lTyV��vfW 0���r���jD7���u�D�k�D�M�  L����}�d���Lv    UO��� �>w �\-�y���5;�Ϫ%>��  �Ժ��h�Vv�<X���8">��   �Ɣ���n `�����9�O�V#�=���*�~*� ���;ey�Hv�<(5��fv    ��#���� f��; [j��veD��ֈzGv�W>�]  ��*�;�	�U�["b��   ��4Jynv �����U���	�j)��n�j  �q%������󤬬�{�xwv    Sk<�F�� f��; [�h�{^D<*��CUO�Fq�>  W"ޔ�0��N�   �F_5�t���2p`˔Z�svl�2v���p�  �bX��g7̣�Νwfw    �15/�n `v��%��������mJig'�Y���  �:����dG̣r��k5�_fw    �Q��u߾�fW 0����[o}FD���ۥ�z��>k\�� ��z_v�<kD\��    ����WfG 0���%ʋ�`[UO���  R��u��p�   �T��]�	 �&w 6�ѳκD\��۩4���>��I�	  L���>�1�Z���D�m�    l�C��#�# �=� l��^�3"Jvl�q-F��T'� �%��:tKv�<+�qMv    �`/�N `���������y���JԽ�|Vm���  L�q]v��     �E}v=�T�����T�[o}VD���	����8/; ��Q�'C-^   ��t�pǎoώ `����J��g7@���V����D���  L��	�B   �iV^��� l&�T �4�N炈�(���:��t�#�ݨ9r�>  bX=F��   `z}ը�y|v ����M��v�[+���z~v  �e\�jv;�s�~v    �n�e� �w 6Eݳ猈����4�ƣ��  ��hܑ�@D�����dw    plJ�7�v��� `6��)F��#bGvd*1�,�aޕ��n  `��<|��}r|&;    �cV���� f��; ǭF,��K
D��j��+�b^�vϫ��  �J�O}����ç�    8%^Xw�>!;��g��qt:�gew�h�".Ύ�W�pz;  v�D�gG���   0��;l6_���3pตh|vL�q4���0�J�� ����|�qv     ǩ���� ���; �e��>6�^�����J_ַ_=眓k�'gw  0uvU�G:A�I�    ����gfg 0�����2�xEvL��u��fw̛���D���  �N#�8cWv�W�]    ��+?�� �t3p���u:��gw���5���0wJ�� plv�2��^   �YP�k�KK_����2p���(?%�&���3N̎�G������  `:��FF����ߎ���    6Ii~v ����cr�Ygu"����P'[�oώ��F��b  �Qs<ޝ�@đ�n;3�   ��S�>u��9?���d��1i�Ư'��WP��ϝ@����i���  �W-��"Z�n    `S5J�ʎ `:��a��=-J�(�&�Y��n���Y7�����  `z�hVO�Z��   `�<�����ˎ `���a���;`������ΘU��SO*%^�� �tk�a���:    ̞V����� Lw 6���w�R�%�0%�,��̎�U���/"�� �t����F���    �(�ý^7;��b�����×E���05J}M=��f6���{�)Q]� �f8�g�\5��(dw    �%j��� ���; �Zݽ��Z���0MJ����џ��5���E���  fBs��ѯώ�g�^�#���    �H��ݻ�� ���; �ڨ�zYD���ӧ�d��<<�bV�u:O/O��  `v4j�,�a��qx�   fۮA��w �5w �z�9'�p�(8Fͨ�W���C�]=眓K�_��  `Ɣxlv�<+��   �u%��Գ�^�� `:�p���7"N�U⑃�C?��1�FG�~3"���  `�<�v:�X��F4k�K�;    �r����WfG 0��Gu��SJԫ�;`ڕ�?p���O��j�鼤��"� ������y4Z�=!"��   �v�/>�{���+ �|� ܣ�h�C�ͰJ#��,-9�|��z��D��fw  0�J<7;a�2��   ̏v����� &_� `��3��=\h}<"N�n���V�Ǖ~�pv�4��w�9l.�UD�?� ��VǍrގ���C�E=���ۋ#bWv    �f8n��8 �'��^���.D����2����g�l�i� ��JǷeG̓���¸   `޴��# �l� ܭ����Q�+�fQ�xʰ����:w������ �^�� �|(Q��B�mT��    �P�t:dW 0���[����DD;�f����͎�D5�9���7G��[  �+�K�ggG̃a�sqD���    R4"�k�# �\� ܥA��Ȉ����u%�:�_�>���z�N�-�-�-  ̟R�+}>�z��n     ��F{zOΎ `2�C wm\6"Jv̇��Q��?��.f�d�g�q���?
�  �灃��ӳ#f٠�yx����    r���k�Bv ����/s���O����'��3�����qƉ�-Y���[�E��[  �o���.��2%?�_    "8�t����1p��Ԉ�F����yT�>q�j������[�۰�y̰5���xXv  D��N���h��<�F}Zv    ��D���{�	� Lw �Ȱ������q-L��Ҹf��{Qv�v�e�Ի�F�:"��� �����v:�gW̒��F���    &G���?���dqX �Cݳ�a�y]D���DD�[룗�C����
uϞ3�ƛK�˳[  �.������wfg̊�R����Ogw    0q��כ�w���� &����F�ø&��ͅk�:��e�l��,�^4l4�ٸ ��V�;��E���Ȟ=�j���    `"�h6�?���p�; 1�t.�(.~�I���/���_�r<��â�/Eģ�[  �^�xk���n��V5ba��?"��   ��*�<������ �15�D��~/�${\#�Gֺݟ�����1udi���R�W��߅q;  ���ãk��1���O�q;    �����zᅭ� �9��t�ϋo�� �;#�o�Jy���옯����4���"�wF�bv  ���^]1tߠўޓǍ���z    �R��[++���  ��;���{��2��sD��n6l-j�)���n//�Mv��Ոƨ۽��xqD\��&  �G#�c����g�L�#���f�k"b��B   @�;F%4釽����ܠ�������q��Fy[]o�yǡ�o�X�tΏh<���ܨqNF  l�O�K\�ce�c�!��v��k|("��   �t)Q����?3��<� sl���u�4>~�,G����k����F�/���x�z�'���qI���F��Eă��q  `�\�/.��r(;dR�ݻO6�e�    0�j�g,��o��  �A#���������������`K�E��8��(וf|l�ټ��t���5�]ZڻP�y5⼈���k"��ܺt  �Xi=ri�ԧ>�2i����o/%�!�   ��U"�k*����- l?w�95�v����� K�tD�DD�-j����L��L�h�K�Xj91��%N�{"bWv1  L��l-4�Zn����IQ�=wqt������n   `�7�����+ �~� s�h��U�q�hD��n  ��U��Q�/����.�V�8��Ak���O�n   `f�K��[++���jd ��jD�Q�o�q;   ����(:��< �$S=����V����    l�F��7�}6. s��`��z/��dw   ��8��/���c�C2�݇[�����g�    0����eW ��Jv  �����4�����[   `���5�~�GJ�zv�vt��5~%"ve�    0�F�(�i//�Mv ���`NԈư�{D���   �Y5�?\h<���)[��~�}���Q��n   `n�K��zx��ƣ�! l�Fv  �c��~�q;   l�����Y[�=���#å��4l/~ĸ   �mv�`0zuv �c�����[�t�/Q>;�[   `�\]��%�����r�w���8^_K\��   ��Z��WV>���2p�qu�������:".�n  �94�Q_�ޱ�g�7ܞ�Q���9�_Z����81�   ��w}k�vA��'��`��̸�N�%�+�;   `��Q��j�~��t�jv�=��w�0l������5���    _�����gG �u�fذ�yB���hd�    qg���Q�����Ȏ�R��9}T�w�WE�i�=    pWj�o]��ߚ���0p�Q��9}�%b)�   �2����ͭ�ѷf�R��{�����OlFyn�xZD��Z    �^�}}}���[v ���`Ո2�t�Y"���   ܣ;���Z��=l_]>q���~��w�)���R��Q�"�ԭ~L    �d��\R"F�! l.w�4��^Qߐ�   �zmD���������KK/�\3<��\;�}���k���؈���hn^3    l�Z�WW~,���e�0c�ޣb\?n'   �b�V#�+%�/���|����Qo��-�,�q�o4�%��Z��R�~���#���	    �M�Ƹ<e���C �<� 3��z�����ؗ�        �����х;��� 6G#; ��Q#���-a�       ��8��\������`s�̈�R��%ʓ�;        `�=l�^_���(� �Q�����.       0������+ 8>� S�h�{^�Ƈ#��        Ht$j��۫�.;�c�_�)VO=��F-��        ����;w��� ���;������ηF�e�        �$(K5�Q;�]�- w�)5�t^_J|Cv        L�F��v�(�! l��;�t:/�(/��        �ITK\1�v4���su��v���5���        �`��x�����g� p��L��^��e\?��n       �)0(Q����7;�{��`J�v{�]#z�-        0=ʧ��K�++��]�=kd p�j�{�B���       �FՓJ�?9��tvv	 ���`��^o��;"���        �F5��,�w�^��� �2w�	V/��5�ߋ��d�        ��{�p\�Y;�]�! �=w�	U#����7Ո�f�        ��x�0�;�};�C �k� �F�a��+�[�[        `�<~0���{�bv _��`�|v�������        �E%�G����^xa+��/f�0a�������        �YV�>}�?�������f�0Aֺݟ)Q �        �A-qŰ���jO	01�!L��N�ե�gw      5���    IDAT  ��y���3r�%; ��a����        0��o������]0�\m�l��~�q;        d+�1�t~!�`��$,������         ""�����+ �Y� �W��ދ��_��        0i~��_yEv�<r�;@�A���(�Wø        &���uz�ʎ �G�� �l��>?j�V��        &Z)�c������ �'� �h����R�-��n        �Y�������fw �w�m���^Qj�5"�[        �{�D��V�����y`��֖z�,��^�       �4����~��e� �:w�-���<�D���he�         ǬF���WV~%;`��l��R��Z��#b1�        8n5j|w{u�ײC f��;�v:O�Q�;�[        �M3��o���Nv�,2p��N��5�;#bgv        ���k-�[\]����Yc��Ɇ���5ʻ"���        `ˬר߶��-;`��l�a�����q��        `�k�oZ��ߑ0+�6ɠ۽(j���zRv        �m�W����(;`�l�A������qJv        ����\XY����ig�p���C���"���         ͑R⩭��?��f�� �i���=$j�7��       `��5�9�v/��fNp8FG;�����({�[        ��q���7�. ;`�����y���K�Rv        0q�,u����ꇲC ���;����m��jD'�        �X�Ǹ����0M�6�������xD�KN        &�mQOh�����ia�p/�t�Z��"���[        ��qkD}|������i�� �����B����       �:%��{m����! �����3�ܽP�=q��        `*�Q��[۳�A�! ��d L��{���f���%        p�ը�.����0���p7�=g�ܸ        �$�Q�st��s�C &��;�]����w�h�;j|uv        0;jD��\�������n�D%; `��}��;�Q��        ̬��������7e� L'�|�z�9'׆f�        l�����;�:��0I�>���}�������#�[        ���U�����쳗�C &E� ����5,�O��%�-        ����ְuY�č�C ��s�v:��Q�8".�n        ��G[%[VV�=; S#;  S��v��3��       �\�xo��N��d�̭�{0��#"��        ��{�޽�d� d1p�Rݿ�=����Y"�1�        �<|8Z��z�����`�̝zᅭѭ��~�xjv        �]��a{����3N��n��\�����7רO�n        �
=l��Uw�>!;`;�s�F4���oGĳ�[         �ͅ��^ogv�v1p�B�h��7F��d�         l���x{ݷoGv�v0pf^�(å�/G��f�         lT����`����s�[ ���;0�jDv��%�3�        �X�(��~k���Vv�V2pf�g��_����n        8^5�3F��F,d� lw`f:����/��         �,�ƳF��[�܁Ye�̤�n�gJ���         �l5⛆��oV;P`ycf��R�'K���         �B�3rf�75��ٻ�7K�����9u���@�]]�}z�iDi��vB6��B��QDVA�eT��`��$�lt��F�y���ˌ^s]>@�:�,��5��:w��̓ ��KU���z���9����-��r����⍥;         6���`�H�C ֊06��~u���         +��t���� k����~e�xg�        �"R�{zaᕥ3 NV�t ����u_n�        L���W�;Jg �,w`����OG��*�        0^�\u�t��H� NT��^�./�         |[J�+����.�p"܁�ԯ�K#�G¸        �{���Y\xK���e����~F�qyD�K�         ��u����Jw w`�,��%)�1U�        `�����^�=�C ���;02����?��         �*G�N�z�+p,܁����{Ѡ������-         #&G���^\�`��{b��fn�s|6��        N� r\:����! w��jMU]�#]�J�         ��՜��f���t�]1p�V37�؜Z�Gĩ�[         ��j���^��C ;0���zt�tCD�V�        `̬�ϜYX�T�����:M]?2��|D�^�        `L�����׻�t�w3p�J��9}>"߫t        ���R\<��pm���`��~U=,"�g�n        �˭Az�����K� D�C�_��7G���n        �0GR��t�h� X�v9n
�v        �N�9�i�u_:�w���Uu�q(E�V�        `�ݖ�����_�&��;P��n�~i���"�J�         ߌV�pz~��J� ���(�h���=ȇrD]�        �;�5r���/�u�`��n��v�#}!"v�n        �N��ϛ����t0YZ���r�����u(��        ������,L܁s���S9E�}K�         pL���O�9|��J� ��w`C�[g�r��v        �Q�5�����J� ���Xwyvvk35} "~�t         �m��ƣ�;v�Ɵ�;���m[����#�J�         pbrD��^=�4;{��-�x3p�M޵댦վ!r<�t         'mG�=upi۶]�C��e����{���~�ƈxx�         ���v�}�m۷W�C��d����{�������J�         ���tV�Νs�C��J �%�Ξڴ;�G�ǖn        `]��N�9'}틇K� ���X3��Nir�6R�S�        ���禅�+��V� `<�:��t�q;        �Dyp����U:��I�{���S�LD<�t         �� ߔw�8�t0�܁�����Y�L�qQ�         �yX��z]>���K� ���8ay���[n�t�xJ�         �{D3=sC޲��!��2pNH�h7�����c�[         �j:���'��8n9��TݏE�3J�         0t�t�������!��1p������O"�O�n        `h���Uy׮M�C��b���j���"ҳJ�         0�R�����yϞ��-��0p�I�H�\�����-         ���I+G�\����nF��;p�rDj��=��ť[         -9�SW�"GL�n���;p�n�w?"^R�        �єs<m��/7r;p��U������         ������?��W���ܥ�~s��K�;         �3rp�����J9^_�        ������~(G��!��1p�GSU��R��t         �*�����+]o� w����s�w��         `�x����+Kg ������\��H��         L��^\xu�`8�J á_u_f�        ��K����3����;�����C�         @!)ův~�tP�1+L�~U� "]��         ��o�,.��tP��;L�~]?/r�a�        0$R��uz�o+��a�j����r\��-         ��R��tz�w�� 6��;L�庾$�""�J�         �����ӽ��J� ��&��\��)�OFD�t         ܍)^2�����!��1p�	���{Ѡ������-         pr�������J� ��&D3���9���M�[         �8��.�Y��x�`���h����0n        `4���ϙ���(�/ws���csj]��n        ����#?k���d�`���k���9�qZ�         X� �%�z��K� ����TS׏�9>��n        �5�o�x����5�C��g�c�_U�H7Eę�[         `,�Z�����J� k���L��9n���J�         �:ZJ)��YX8X:X;�������C"�Ma�        ��ۜs\�t��֎�0&����A>g�n        �t[ʃ�:��Q:8y�0�V��Sġi[�         (���JN���U����È;��ޯ=ȇrDU�         
�f���Ӌ_���!��3p�v����q{]�         ������^�oK� '�U: 81KU��5�7�        ����nX�����!��1p�t����S:�J�         ��ْڃ���m{@�������9R�ݩ�"⾥[         `�}%��f��tp�\p���n��ʱ?��        ��̶Rk����m�`��Èȳ�[����#�K�         �(���������}J� �&� �Y޶mK�n�,�         #�K����o>|���C���;��k�Mk�z�v         8a;ڭ���m�^�;��{��������n        ����:8�w�+�5wR�����,-�?\�         ���7����e׶�!��K���ggOm���"��J�         ���N��R����!��Ð�UuJ�ӵ���-         0����J���o���U: ����nn"}θ         ��C�A�)��qf��;�aH�{����3qn�         �kVV��g�}z��v�0�޽��[n����GJ�         ��yD3=s��;w(,���Y���O����n        �	��fz溼e�i�C`��CA9��,�X����-         0��t�������!0�ܡ��n���"⿕n         ""��� �ʻvm*���
���8"�T�         �;R�����yϞ��-0��a���T��#ǳK�          �+Ez�ʑ�����uJ���1p��#R3W�/"��t         p�r�X9|�9b�tLw� �_n��)~�t         p�r��W��r#w�8�A�U�m��         ���Oo��d�[�~h����)�kJw          ' �s���6����~S��K�;         ��riSu?�#R�g���7S�_.�         ���¦�>h�����ISU��"~�t         ��ҋ��~g�
W��u����r��-�         ���^\xu�7.����կ0n        �1��U�U�wJg��1p�5ԯ�/��*�         ���5M]�J�'�t ��~U�0"]~W         0QR�7t�\�Ɓ!.��~U=?"}8�W         �H)��;�����Qg�'�_�ϋ��         0�R��vz����Qf�'a����r\S�[         ��rD~�t����!0���-�u��R�D�         ߑ#�K�>P:F��;����SSʟ��N�         `�����Ӌ��Qc�ǩ��>)�|UD̔n         ��j��ҙ�����Qb�ǡ��s��FĦ�-         ��[͑�3��]Q:F��;����ϑ>��         ��[͑�5��}�t�w8MU=&G�!"N-�         ��f��M��եC`���=h������V�         Y�V��M-,\S:���;܍���s|>"N/�         ��~���:5?]�V�p�U���tSD�Y�         K)�S:J��02p�;ѯ�F��#��-         ��9�Z�ɝ��C�C`شJ��Y�v9n
�v         `}����fn��J���q���rU�@�t("fK�          �.�{������*]��w���Uu��t ��        ������?���J���0p��8��ޯ�@��+�         L�{G�؟��W:�A* �-���l��"bg�         `b}-��Ν�ʗ�w�(�����TU;ڑ��J�          �y����Ç��t��* ������q;         0��V�������RܙHG��z*��ȱ�t         �w�m����۷߷t�`���ɳ�[��ƈ��         �N��V�fg�S�6Z* )o۶�i�F���[          ���V���|��K��F1pgb�:��t "T�         ���J+�s���B������]g4Ѻ!��        �Ѳgj��;�J��F0pg��ݻ��4�����t         �	�_Ӭ�[vm+�-�����:�^ͦ��#⿖n         8I�؉|n���^:֋�;c+�Ξڴ��E�Ǖn         X#�Iq^ZX���!��K��Nir�6R�S�         `���N+����Q:�Z�t ����nn"}θ         Sk��|�Y�*k����������DĹ�[          ��#�M���g�}z�XK�t ���w�t��[�,E<�t         ������������!�\pg,�}�:+���i�v         `�<��L_���ͥC`-�3�rD�Y<���c�[          
8����]�6���e��H��>?Y�         �����UyϞ��!p2�Y9����G�g�n         (-Ezbi�J#wF��;#)G����9�]�         `X��,-]�#�J���0pg������?S�         `�����W�3�R� 89"5U���xI�         �!��No�)b�t+�)����0n         8�h����f�����X����ȯ)�         0B.m��eF�
_TF�r]�)Ez]�         �ѓ_�T�rD*]������\տ�r�r�         �ѕ^����JW�=�C�����H�S�         `,�x���«Jg�]q���������         �P�W.Wݷ�΀�b��P��կ�9~�t         ��I����_-�w&����_u!"�^�~         ���⍝��7���f@�P�W�#�e�	         ��R��wz�o-������ѯ��G�GD�t         ��H�_����^�"���~n���0n         �h9"��t����!`�Nq�u�����*�         0�r�x����J�0��)jy�����'¸         ��9������J�0��)f��~"E�TDtJ�          ����f�?^:��d�N�\�I9�"b�t          w��#=w�7y�&��;���s��FĦ�-          ܩ���3��'J�0Y��PMU��#}.��         �]3�|ɦ^���!Lw6LSU�ɑ����J�          pL����t�����Tգr�χq;         ���Z�S��וa�����u��ȱ?"N/�         �	YJ)��YX8P:��f���    IDAT�κ�W��"��qf�          Nʑ�JO���*��2pg��������8�t          kⶔ[?�Y��a<��.����A>�W�         ����=Zq����_�.a���斫�"�`���t          ��1h]0}����t����5u���?�8�"�J�          ��n�<8zq�oJ�0>Z�G����s4n         �gDjݰ<����C.��&���v�S���t          �y�>w���O�F��;'m��v��u("ߧt          E|%��f��t��U:��v�����         L��Vj�?�}�}K�0��9ay��٩7F�ݥ[          (+Gt[���Ggwؖr�R� FS���ڴ;#�J�          0T��:X}��Ç�X:��c��q�۶miZ��io�          �ҿ���9���/�a��J0Z�g6����          ܍=S�|��۫�!�w�Y޵�fepcD<�t          C�~�����e׶�!��T:�ѐw�w��|c����-          ���D>7�z_/��s��{��:�^�����         p�D�)����a������UuJq}Dz\�          F��uZ�4?���!/ܹK����5��          ���6�|cޱ���!/w�T�v77�>O(�         ��xx��zm>���K�0���y���� :"�-�         ��yd3=s}޲��!�T:����^�����-�         �8K�Ym.J_��m�K.��my߾��-���q;          �/?�iO]�w��T���a�NDD�v�x��9�n         `b\�����{�̔a8�s����>?Y�         �ɒ"=���t��;�/G��������-          L��㢕���s�T��2p�`9"5u������-          L���╹�
#��f�>�rDj�����gJ�          @DDNqIS��#ڥ[(��}�>n��AD�\�          �O��T�����D�O�~�}kD���          p.m��eF��>a���-)�kKw          ���/h��9"�.a��O����S�ו�          �c�^����JW�q�'�r������;          ��xy�~g�6�s����_̑�^�          NT����kJw��\ps��~�q;          �.E�Ŧ�~�t���1֟�<R~w�          X+)�;o*���0pS���"���         �1�"��ӛk�֞���W�"�e�*�          �!E��N��;�;X[�c�_חF���q;          �-G�_����[:��c�>F���)���.�           G���^Xx�ֆ���X��KR�+"b�t          l�9������J�p�����\���'ø         ��4�9=ofq��C89�#n��~"E�TDtJ�          @A�9�sgz������f�����U1S�          ��j���^��C81�#���s��FĦ�-          0D���3��gK�p��GPSU��HWG���-          0���ȗl��>W:��c�>b��zL�t}D�V�          �X���⩅�kK�p��GHSU�ʑn���K�          �XJ)��YX8P:�cc�>"�u��ȱ?��         �xI��������!�3�Я��E��#���-          0�nK��#��/�y������C"ǁ�8�t          ����ъ�����t	w�U:�����>8r���          p��b�?�߶��K�p�\pRG���)�P���t          ��[#Ο^\���!|/�!t���?�8�"�J�          ��zn�sg����tw�*��v��s4n         �usv䛗���[:�;r�}�,���l�֡��U8          &�Ws�3���ϥC���C�HUmo���0n         �����Z7ݾ���C����8R�ݩH#�}J�          �$�ukup���ݥ[0p/.o�:;��ƈ��          ����^=��mۮ�!�.��dyvvk����(�          Ŀ����7/.�k�I�{!y۶-������          04v�S��۶o�J�L*��g6���づ[          �;�_gup ��9W:d�o��k������xx�          �NݿiV�[gK�L�T:`��ݻ��,-���t          p����⼴��o�C&���ɳ��6������[          �c�w�V:/���t�$0p� ��NiR�.r<�t          p���3�>?}�K��w���.W�)M�k��         `d=�YY�6�}��CƝ��:����&����-          �Iyd3=s}޲��!���}��{�����8�t          �&�tf�˳���W�� ��;�r˭�IO.�          ���ئ=ue޵kS�qd���}��[����[          �uqA�߿��}�����n4G���-          ��I���o�����)�2N��H�h7U�'�[          ���r\���ty޷�S�e\����j���"ҳJ�           '�x�w��1U�e�������}��9�[          ���S\�T���v�Qg�~rDj�����ť[          ����T�G���I��;A��ۻ?W�          
�k��eF�'�����[#�ϗ�           �I~ASU��t�(2p?�u�����;          �a�~���w��E��iy������;          �a�^֟��Y�b������)�Jw           # �+�U�������5u�����{�������{��g8�z�oZ�%QR��֫�:����(�] H
��&m��i�)РF�I�4E�^P�]4��8�^�+���^t[�V�V���;���~��y�ɱV�.�g漜�|������ ��{�'�G��          �W~����!W)�u��A�P�/#�           ے$����q�sd���]���E$�?�u          �����&�~��9�L��g(勿��^��          �$ҿ�0>�?�:GV)n��|�7#�ߏ�\��           �F������k��d����(
�i���          �4�������Z��OX+����/#���Y          �}+�4�ۍ��W� Y���1k�¯%i�QD��:          ��U"��h���Z�
������$����          ���H��כ&F���A�@�="��_���?���Zg          ��4ҿ�4>�ǵRk��^��4��i(�          �SN#��������Aj�@������H�MD4�:          p��*��Z�����:H�؂{yp��4�}5"�j�          �R.�_���Z��Yp/��?�F�8T�,           ���$�+cc/�:�^;p�r��4��GD{��           �˷K�/�:�^:P�R��L���#ҎZg          ��夒����їjd���{)�<"�fDt�:          @u�����GGP�${�@�K��c�Ʒ"�H��           l�|Tr_j�y��Av۾/����$���u          �m������:�n����|��$��I$��          p�f#�_l��AvK��v�j��@ɋ��          �>q8"����чkd��˂�j�x�����D�:          ��Mr/���u�ݐ�:�N[���E�RD�u          �]2�F�Ŧ�����������P]���          ��֟������'jd'훂�r�P���ň�x��           �4����xq���t��E�=���O�q��Y           ��Ѻ��W�kd'�������\��BD��u          ��Kr�/�k�^���t`��\_����L��           �������Z��m�==v�����Z�q��Y           2�3���i__��lWR� ۑ�8�Y^]�fD�Wj�           c�nH�&cc7jd����':�+k�Pn          �T����fZ,v�:�V�W������Z��H⳵�          �a�ʕ�����õ��M�=��[˹��>[�,           ��'�������:H��Z�F�Ϸ�#�����          p�y��\��dzz��A�&�;���N5���_�r;          �v�\���i[���M����7��W�U�Ɨk�          �>��r]���ǎ5�:�ϒق{��Í�s�o�+��          �|�TZ��,��3YpO#�ʳs�F���          �_$�>W*��$=u���Y>M�
�iD]9_����J��           �7I$�����G�O6�:�'e��~�ܞ��#ҿQ�,           �U�__����4���Y>.3�4"W.����o�:          �~�����?�R�=�4")�y���:          ��r����<D���I�'��          p �z9_��,��k�V����D�Z�           [���|�_�I-SԴ�^��7"����           @DD�[�|���2A�
�k���D��k�~           >)��R��Oj������]��]�w          �3���J���T�W�y������$��f��          @�~g-_�o����^��\(�N�FM��           lM��?l��{���zQi���"��W�          ��%i������ݓw��KJ��oG���^�          ���D�_5������]V�+"���x           �"�H�q|����Kv�t^��3"������{           �uiD�w����n�`�
�B��#��3��          ��4��;�c�b7�+��B�+I�2"�v��           �L%���Ɖ�?���x�}�P��$�?����~6           ����ɯ7M���N>tG�k��_M��#�a'�          @�l�������?ީ�X�}}���J.���hکg          �i�4ү4����x؎�˃C��&��;�<           ��J���<>�g���{.����/����Pn          8�J�$~�~l����!�Tp/>�&��FD۽<          ���Z������ѯn��.�����K#�ZD��3           �W��$~�al���ܼ��{�P�\���#�};�          �o-'��5L�����\p/��OD$ߌ��[�          �a)I+_n���w[�iK�R�p.��VDto)           �|��GG_�����B����#ۊ          �A3i�K�#�UsqU��b񑤒�=�          ��f6"�����7�v�]����Iķ�Hv&           �tZ����ɫ?�Y�~�W���"yA�          �{Л�6^X8�.��;�����*�ӈ��g          � �J#�b����O���ྒ��U���          �A��H�_�?z��~��
����P]��v9           LQ��m������?K>���B�X�Ʒ#��^�          �@���V~�eb�ʝ?���=���O���          ���Kr�/���A.""���+��+"N�,           ��������$�-�սi��u2           ���_HJ��X��           p������)            W�            ��          @F(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�       ԅ��    IDAT   �	
�           d��;           ���          @&(�          �	
�           d��;           �P_�  ��ب�����X���ήXik�Ֆ�Xk��}��-J�MQnj�4��4I�����r�mlDDD��jD�PZ�敕h^^�敕h���}v.��E�͛Ѱ�V˿2 pIs�X>t(nvu�RWW,vt�ZKK�����~�+Mr��P���0J���DDC�u�rԭoD����1��qJ��J4--G��B���š��h]\��� �߬55�bWW,vu�BgG����jKK����ZkK����zCCDQjn���J]]��qm-�4�$M�a��|I��J���D㝹���h]Z�5�27���7�c  �j��%:;c��3::o����YZ���4�(��l���z}�_�]*�hX+EDz{M�֘es첸���o�]nތ�� �i��r{���e��cs�rg�h��5*�X#*76F��ֈ�ף�������4/�D���ͱK��RD����l]R��_ ����������}1��������ˇ��<K��J�������==�SS�}�Z�..�y  6��b��7f��b��7f������X��Jno��[_����蘙�#���=u-��]����H*�=� d�Rgg��퍙�s+�==���kMM{$M�ui):fg���tt_����hS අ����5n����#Gb��3J{<vI�4Z�cf6_��y����6D "��F �==��,��]n>�Q����,u��qh~>:gf����>��ttܸ9kD�I
� p٨��냃1U,��ѡ�����ZǺ�������ѱ���Q_.�: ����B!��ŵB1�t�y�}���ף�ڵ�������= اJMM15T�k�BLō���/�oá����������)�� p ����T�׊�[c���=/�oY�F��\�E��X\���_��   7��o�Y���Z�sG�d~��nc#O]�5�2:##Ѻ�P�X@(�@���\\��c����냃�G/��r�J����+W�x�R��8� �S��b���;q<��Jkk�#��ٹ��ŋQ�t9���k	 ؆rCCL;�'O���p���D�$��u�J����GE���虚r�6 �����8~,F�����1w�H�>�4��E����˅螞�u$ `,vu�ȉ1z�D\*�J[[�#툶���:�K��x�r��	jB� 2f��-FN���S'c���Xki�u�]�P*m.��p!�nެu$ ২������=y*FN�����ZG�uI�F��D]�C.F�Ą d���#q�ԩ�R��y]-��Q�t)�.^�Ѵ�V�H @�f�zo�]N���P�w9�	mQ�p1�.]���K�P*�: P�J]]��ة�q�ĉ���u�]��i����K��������	w Ȁ�������31~�h�;<y��������������а����w�������Q�T�\.G�T�r���뵵�X���4����8��{q���~���r1v�x\>s&�<�`���Q�uuu������Q__����c�;c�\.�9n�ccc#�ۓ��||�����y�Ni����'�{/z�'v�� �����O����L_ߎ>;I�hjj������[��=����'�V�4���'�mll��x�Θeuu5�����؈¥Kq����?�Few Ȝ�ޞ�|�L\<}zǋaI�Dss����θ���>�n��$Iu�����.���c��Ϸ���l�����(~x!N��~}�a���� �7�\.Ə�K�OǕ�����}~]]]477����;㗈�ֈ>�g)�J�����kD�q���q����l̆H����F6����Ň�<�ǎ����������hii����hnn����N�T*�����������p��I�F��H�z��8��,���V(����G=xϧ�$I������)��4Mcmm�'�*������+++������8����3o�33;� ��Jkk\x�Ѹp��10p��kjj����hoo���֟��)�����O�[Y\\��Y��z/^�ϼ�N}�a�*�J l��C��s��Ň��lｗڛ����إ��y��.w>������˛�,KKK���/����o��K�"1v�����o��~(Vwh���Wkkk477Gkk뮯�J�X^^�Kc��(�������ߏϼ�Vt]��C��;�`������?>rv�E������舮������,�e���j,..�͛7cvv6��涽0�P.���(���76��I�;�ZZ��#g����c��w[ϸ3Qyg�r�Ծ���۱�����������������=,M#�j<������Qw�� ��K�$Ə����+>�O�<Z����ͱJggg���GCC���7i����J,,,���|����͛7��͢W��b|歷��7ߌ���N |�4���'�'��S����QSSStuu��Ç7K�Y�,//o�]���b~~~�ű��7��7ߌ�|+�n��� ��Ykj��><���O�K�$���~b��5�����M��Y��F##��?����;|�T
� �*�\\>}:~��_�k��ﯯ��ÇǑ#G6����5�4���Ř�������~���
����q��Wぷ߉:�0 �q}` �}��|������/I�D{{{���n�v��ݴ��sss1;;������ye%>��[��+�Z������x"�?�D,tum�������������ꊶ��]H��*���F7n܈��٭��4
}��j]����`ǭ����O>�x<��۷|SSS�����Ç���Ù���ԛ������-ޓJ%�.]��_y5
�.�RR 8�nĻO6.�>��X���舞��8|�ptvvf�x�*�J?�gYZZ��3�����[o��W_��ٹ]H	��; �RSS|p�\��٧b��sK����Eoo��?r���#��4�����~�zLOO����oYZ�ӯ��_{-Z�ᓴ p`%I\=y2���31><��[���g�k7�������ͱ���̖
d�J%���~<���G���.���k��+�}����cQnj���$I���3zzz���7:::v1e��o.�^�~}���~=���w޵�  ����x�����G�R9,I�8|���<K�6J�������q�Fܸq#�]�kkk[��{j*����{�E��y po�$FN��w�y:Ǝ�ҭq�ȑ�N�~^#�q�F\�~=nܸ[$�J����}?���v1%�_
� �V���g���O<�-,����EơC�v1a6������DLMM��-�vZ����v<��w����.&�����ŅG��?�L���T}_CCC������@9r�<Q�^���ǵk�bjj*�_����{�������>ڽ� ��������|\y表T���$I���+���?��0'�_������dLNN���j���,-řW_��_}5�X4 "�����?Wx �*�K���������t��l�499SSS[*��.,���g^=���]L	 �O��Ņ�g��=s��U�������188x`׈�_�[^#���^�n�pa���� ;h��%�y�x�OE�ʉ����(
188�ow�؎���������Ѫds����r�..�rB ���I��>�?�l����$I���?��|����	˟�\.ǵk�bll,fgg��o���x�b���]L �����x����ӧ�.����E�X����Yj�i���c||<���c���ٛWV��}/μ�Z4(��]����k?�����U�]��ۣX,�������t��4���٘�������wGm]\�G��r�~�N���H�$.�9o|�٘?r��{�$�����5�\���w155ccc133S�}}����K�_._��t�(��(55ŻO6�}��vlO�$�9�B!����~�4M�ƍ122��ӑ�w�ԯ���7ވG_�n�,-�AJ ȸ$��=��٪w�hmm�b��B�b�],..���X���E��"X�ҥx��/E���.������������ųGZ�bi]]]������Ptuu�A�������&sssU�Ӳ�����8���b �)�z{o}(�*�������`EGG�$�������d���T}�o��B��w߉�|3r[�M �$���L�����پ����y�	����r������x�'��	��� � ���s���_�b���������(�144�U\�OZ[[�����R�t������w^�����*w� ��f:�����sq�P������8v�XtW��;�R����T\�|9�~C�����}�h�r� ��RSS�����ݧ��J]�]�oii����(
Q__�	����Ÿz�j���Uu�����x��ߊ����A: Ⱦ���x��<�xT��P^[[[G>���*�:���7oƕ+Wbbb���:o܈g��f]���  �����瞋�b���{zz�رcq����i����T\�r����� ���7�}����Qp�m���=������MMMQ,cxx8� ��V�Tbrr2.]�KU���1;O��b��=H ٰ|�P��/�����.;��r���ǏǡC��(��6;;�/_����^[_.�ï���h��C| ��IΞ�W���+U�?:::bxx8���J�R���ŕ+W��]�o|<���7�oll�@�Tr�����/~1V������+�����CJ�R\�z5�^�Z��y��>������b^ ���5�s�����$Ibpp���ʇ�r�J�~��x򥗢����Pp�-Zno��>�\|t���^���'O����K�4����p�BU��._����עcff�@mTr�x�s�ě��|���������cǎEcc�%<X��ŋ155u�I̶�����>���G� �6���/�rU�tww�ɓ'�.�K666bll,.]�tע{����ߌ�^x!�VW�(! ����c��/�R�����ڞ��8u�Ttvv�A��gcc#�^��/_�k�=W�ęW_�'_zɆ �\.�y��x���G�.�>uuuq��QkD�hyy9.^�XUѽuq1��ַ��;��Q:�>w �V�ćg�����R�����K�����ɓQ(����yp\�}'�ﹽ�@7���  �$@-$E�vK�i˒��e�H ���o�R3U�^ޛ�yy%˲=���Nfۙ�%oZ(�)�ľ;�h��z��
�Ⱦ�"ٷ�流U�s.ȯJ���9��;�,l��ӹ�BwM ��'N������(�#""����l�q��r7}N���|TTT�`0D)]rs����������c߱7`��|DDD�$���܁�x�[v�Z�(--EVVV��%�P(���IlY螲����}��.E)�:�>z���j�8�Z�����KyQ066��Bw��*���&�{�P����|v6�{�q�n󌨼�F�1J钛�����0&&&�,t/¾cǐ���tD���DDD۰d��wO<����M����(//Gaa!�U �2�����ߏ�-:�e�������T���>�gރ��{ڤX����[^^F__���6}���b�o~����-6;�����XE9��Q�n��4--UUU�o�C*�z�`�/_���0�[4(��ž7ބiu5J鈈��g��|�3�7}�b����QJF����122�˗/o�v)�ԁ;�k�x<QJGDD����wl댈���Y]]E?�N���|>4���>:�3"Jb,p'""ڌ��҂��߇�V��c���(++�N��b@R122���a���I�O|��ǏC
��������q����>��-Rm6jjj����d��Ӊ��^x�8TͿ|�����NDDq�o0��GF_c����zTVV�6���z��ߏ���M;��^���_��"��Qb��w�?�ᚚM�3����D^^^���f�����ۻ��yF��Cq��Qbp��]9#���͆��j���G)mfnn===Xݢi@��8���O����dD���DDDxRSq��'1^V��s����0�7��Aѷ�����>Lmѥ�19����ߐ>?�dDDD7O�$�߷��ߴ#GJJ
�������t��,cdd������gX[��_CiOO��<gA�~�i�dX#>æ�myy���X\�� ���������dDDD��DI	�}�)x6i��hPRR���h7i�D�XXX@OO���7}���y��_A��G)ѭ%K��}7��s`�3"�Ʉ��J���D1m�,���� ���It^/���Py�b���)+/�{O>��Փ�555�"���	���m ���B����������Y�X���Oc��0�3B�����1������g�.c/aߛoB��E)ѧ#K.�y��{驪�iiihhh�3q`rr===�����p�O�ܑ�(&#""�y!I����p��ț�$����;v��QGOO��`�g�q�����QLFDDt����Q���������k���8v���(%#R܉��>!���ÇDWs������_�H0��� ._�����e��8��_�kŬ�5�8����IOOǎ;x�d����Aww7��t>��������(&#""�>Oj*�z�YLF>d�h4���Baa!�&Ed[�^/���133�
a��Ǳ��	`��""�X�j��7�{�M��t:TUU��� ���f������.W�=)���v��ŉ��j����gDl(�\.�����I{�����}r*�Ɉ��w""��yRS���=��M6(SRRP__���dt+-//���+++��p����QLFDD�9Y�p��A\��. B!�$I���Dqq1�����Goo/&&&">���p���Ү�(&#""��ta!�z�YxRS#>c��QWW����(&�[��t����Mn�)�������M^�#""R�xy���g��ɺ$++uuu0lRDF�mjj
��ݛ�DSq�����͏��(Fɒ�3��gD())�Q�
������h���4� ���KT�?�dD�`�;�w ������:�t�(&��A�ebhh(b7w�׋�?��{z�����(�zJ
�y�/+��Ljj*ّ#A8�NtttD>|�e���C4��D(�pDDD
zv�GAH�Q��!kb��|������L��<��ᜍb2""�m����$)>��h�6�������/ba��FV���ǰ��E1��xF�|�����с�����T\�t��@ �Ɉ�K��ҏ����HM=�w�瞍x��N�CCC***��pHK�E���Պ��9���g�Z-�kk �ccюHDDt�B��x�E�rs#>STT���&��(&���l6#77+++��Q
���B�����DD���F��O>����G,KMMŞ={��������h����^����ޔ44 cnVň�(6t:���3�ji����b�����#���v�j���˃F������3�&�a����DD3�{F�s�N�%�Ʉ��<��nx<�g泳1YZ�~�|���܉�(i�B���G��9�&��jEKK�Vk��Q4�L&���ceeE�K��*)�J�E���.eex�����N�]�v�����b	h��U����V�V�TU�hp�M:y�^����0R]���B�ڵ���	�b� ++��|a�!�õ��y�Ȟ�P!!�ﭥ���/}	��%�)))�Ν;��룖��C���8���+ޚ�j1�cL+��OO�������&JK��6?#jjjBqq1�M(~}���\�f�����A��e#��3�QR
j4x��г{w�g


����N�dm�fˮ��٘,)Fq?�
�DDD�C�Νx��g��IOOGKK,K��Q4m�fdd��r)�<�5�0�Ѐ��q�./������ъՊc/� W^��$I���Cyy9_�Kpz�����x��P    IDAT<X]]@L��Ó����A6 ""U,:�ŋ/`1BWv�F���F���p�����"6?���hU�����H[�����(IX,8���!�p���hDC=2g�a�-4�`X�NDDIg�d_z�������<�M2HOO���B(
�w[,��DQ� �^�
	��(i�3�݋�>񖙼�<455��XIIIAnn.�UX�t:��@���K��ѭ2���c/���7ޥ������d�x$IBNNΦ\�9���Aq_$��""��e��o���O�f3���a�٢��Բ�U�刷����c9ӆ��~��GDDѳ�3�]�v�(����byykkka�!��uuH]ZB�өBB�ۃ�DD�T<��8�⋘��Q�7�hii��n�r2�f�999p�\�WS��L��AQ� �
_���n�8�Gp�;"L��֢����M&!�V���<x�^����͇$	�55H[�&�>SE�x����MIQ���lhii��d�r2��Z����Ul �����B���B�p3ѭ6ZQ�_��
�����g���('#�	!������t���BV(b_�ʂ+7%=�|A���n?!p⑇q��;#L�����(Ii4������cii)l^�$�TW�����
	�n=�Q�p[,��K/bɞ�8�q���l�r2�%:����X^^V���o0`��×��v������,Ix���г{��V��Ν;����dK���ʂN��ܜB�v!0R]�wY��$"�[k������7�7n��h4QNF��d2!;;;b�U�e�(��Va����V���o?��Z��|AA�vIrf�����a��6f��Q�������Q~~~��Q,B��p�h4��r)=���r �##Q�Gt�������ªՊ_��"Vl��v�{���N�ʵڹ���z�X^^����Q�ܑQ���ݨ�$���O�g���`�U�t��
�٬�aL���A��#{|\��DD�pF++��C�G@�S�///Gmm-D��)��t:���aqq���a�4�VT���:�O��DD��w����>�P�����r���p�B �����`~~>��ɪł��R���@�PODDt3dI»O<���;�yFD�KOO��b���T��f��A����*�#�uX�NDD	o9#?��?�ے�8_PP���Fv�kltG�������V��Z�]�ye5��(��$	�}�Y�S�OMM�޽{y��IMMEFFfgg���l!0QVM0���1uQ����o?��b��(..V!�2�F������­p޺ٌъ
�u�@�N�DDt�56���OA���9I���Ԅ��B�Q,�j�������2�����=ii�,+Eig���NDD�HH��ֳ�b(���l�)2�L��̄��DPam2SX���E��X�NDD	͝��c/�w�rq{II	��Ѧl6�z=�����Z-.�ա`h�U�э����O?��Z����4�ݻ�!��(^����n�cffFqs��:;�ѧ7QV��|�s�ۛ������B2��$!''���XQ��k2a��e]]�JDD���j���ӊ��Z��v���P!Ń�~#���IM�tI1ʺ��a�;�$Y���S �������gD��hDVV�N'
�*3��2�;:�B:���w""JXkf3~��X�pMSii)��������b�^����
�j���AQ� ��
鈈(n	��}�;�-���������`@VVV�"���R�VW`��V!ų��B��_@@���h4,�mٸ%���cii)l~�l�TI1ʻ�Y(FDD7e��oEx1O��bϞ=�E83"� �@vv6���_�s��c6?e]ݐ��Q���h��������v*No����(�x��둝���}��Z���(.�����ҺɄc/��E�]q���
QNE��b��d2��t��t:�TW�����u�Q<����ݼGq�f����Z�b2"%z�YYY�����c���#cvV��DDw���x�K�ïp���j�{�ndff������@0���b؜'-΂�uu�P���>���2����T�K��thii��bQ!ţ��"�B�b�b>'�]���BB""�w<�0�[��xFD7J��!;;.�~�?l~��&�*�Sl�D��DD�p�Z-~����U�������QNE� ---b���`�XY*:y�6m�¾�q~�>�9�͆ݻwC��m�h3:�YYY�����.F���=6�4�ΩDDD��d�ፗ^��h��(ng�S�4�v;��b'�U�vʺ�!T�FDD�k.;o>�E^���thnnFzz�
�(�mU�d��m����_�tDD�.�}��߯8�3"���Z��N�aE�B`���',ss�$�X�NDD�E���S�Н���eeeQE�$--F�Q���k2�Y���NH��ADD����GDxَ�jŞ={�qI��F����LX��,I��Fa?R<�Q�[OI�/��B��v�b�v�)v�^����asKv;=
��THFDD�ȓ��c/��u�9ln��<�ժB2J�n����ass�ـ,#wtT�dDD��kk��c�gD����<#�O�E�J���TW#o�2�
/��"�QB���ѽg��\qq1������Qzz:�z=\.W�ܪł�LJ{zUHFDD�n6/�>�y�6'���x�$�:�������F(�f.��b���]���|*%$"�X�j��/=�P�:B455��p��������Q,s������I�Q<�8��XVx�N��`Ϟ=���P!%!�������BÀ��"�-."S�1�'񌈢A����p(6B
IF��P�����J	����DD�0zv��G�߯8WPP����('�Df�X ����|�܂�Y y##*$#"�X����c/���6g6������U�D���`@FF���!_w���h�tQ*.u@�� �����x��Oc��\aJ����
��D��YYYXYY�����(+�}z�}"""�Jq�o>�y�������6���~}1���@��Җ��	HDD1�gDM:�v�]�R@��Di	*::��� �(ְ�����LA�z�YȒ6�p8����p��Ͱ�lX__Ǌ��M�EE��faU��NDD�ǯ���_���z�{��QaS��f�F���bff&lΓ���tJzy�]qa���ܻWq���
�
�cD7C�Á��9x���'1VY���^���	HDD1�������Qqnǎ��ɉr"Jt/�����wݭx�$a���]��_��!"�����N�CKKψ�����X,���
�[7����@YWXIE���DD��RSq�/)�隚��={�@�p�ѭ�p8���~-���@q_R��$"�$"�}�)L���MI��={� ---��()��fh�Z�^���Άѳ��
Ɉ�(�L����O 
�
QUU�B*J�$!++333���ZL�����%v#"�k��T���+�]���Q��Ct+h48LMM!x��$��a���/��<""��-Έ���yFD�MJJ
�f�b#���LH����Q�m܉�(��$	�����p���F^�D��f;B&KJPu�W;%�Kw܁�;�B���v�]�T�L�V+�~?��ɞ(-E���H]^V!łU�o��%�O�v;oţ�N��"33S��l�Ʉ�Lʺ{TJGDD�f�a�/��E��ڰ���\��֪����N���f���dY�fn-5k�T�������bψHm��� ��������"8�&a��#�,p'"�����cXa�R�Ѡ��f�Y�T�l$I�������A�͆��%���b���S���*++QXX�B*JFv�]��Y�0^Q���|~���ZZ-����X���3��hii�$I*$�d��둖����鰹E�Z����*$#"�X�3�Ƌ/��q��'Y,�ڵ�/�QT�F�L&�n�s�90������!"���3"�6�n�����N���r�uwð��N8�Mpg�����HU:[�����x�EUJJ
v�ܩ�y~��ݻw�����Դ������,B
EaYYY(--U!%��n0)))as��T�)ū݉�(��z�~��䄍k�Z�ڵ�F�T���v;����N�f�r�����b�����l��q�^���&��GQ���q�G�����DD�<xFD�����j7�O�n�w�Hm�[IDDqi�l��{Tq���yyyQNDdff���Bq�Ç�<73������~F����dB}}=;�Q��t��Ŋ��e���(%���2t5+��������*��ˑ��6�$���3�*�""�X0\[�����q!`4UHEɮ��v�=l<����<��V�B*""�<#�X��h�k�.h�'��|�߿O�TD�c�;�!��SOaM�ˀ�jEMM�
���(++CVVV�xP�ŻO?���%��]M���膪��THE������Vq����yDDIb�lƻO>�x{GYY�b�1Q�Dz�b%#>��
���Hm��{�qŹ��*�c�h����,N�{P�TDD�6�Q�2�LhhhP�;�?f
���hs,p'"����Ҍ��q�N��;w�MWR]}}��f�\NN�wo�QT-�l��窫���#����|���Z-�fw1"��'�{��"�LF-Z�6�_oS.�T������"K�y�)�n���())�~(�O���hllT\�t�q&JKUHEDDj�ź��,��o��&R܉�(�,�l8}���suuu���b�N�CCC��f�;��LA�
���(d!��O��ׇ�egg���#jkk���6�����{�Q!EK�Ν���j���E[ZZ*����{�&S��Z:���tQQظ^���}�(�222PVޜKǟ|~�%�Q����BZZZ���ՊS��<�,p'"��!N<�(
%��򐓓�B("e6��
]9663���(1u77+^�g0�c�)۬3�;kk"���I5��(�����Ģa�!%%%���_7��![���ªՊ��P�۱c�
�cDj)//��jw������F?Eψ(^H���;wB�ф��4��oI��w""�=��Q)))����~ �-TTT�b���/ef���w�����n'wz:>��`ظ��t*�"��b����<l<$I���!$qۈ�(�|��#�*�~������<E��:z��c��]R��(���L�jQQ���TE���E�P��yo�%"Jp<#�xc6�QUU>�q�Q6m�X��J""���T�z@��X}}=�\XQB���^�3��}��ఫ����n��{T����B�ΓD�������a��\t�ݫB"""�]F��0�� @�׳q �,�����Ź�}T�葈�C_C&nI5�L���T!��L&�b����!��w""J<#�xTTT��6�d���囔����DD>x�a��(.��bEjj*���;��4���c�B�;ş��VT���F�RLB`ǎ�/�=x�
��Q���t8��g�jkk�E�bZ^^���&�V+����V"�D����S=�8W[[˦G�
o�]t8p��;UHDDD�ψ(����AR����]w�i#���DD�f
1�Щ�`0(_�Cc��ˑ��6>]X���:ѭ�jq�A�fx�J� ==���a��'�_�DDDt�]�w7�iia��999*$"�1uuu�(t<�hi��_%����zJJ�x����b���b��c3"��3"�wf�Y�i�$�GQ!������b�,N<�b�kv�x�Ygԓ�߇ �ŵ�w܁U�5l<''YYY*$"�qHQ(���ta�
����VY�XpI�S�V�Ŏ;THDt�RRRP��/���d��DD�v���6���Q���(��f�����t:|t�
����v�%���2�)4ǘ,)�(�����Ŵ����S�$f�ۑ���B�������x�v�����@  �ߏ`0x��F���K��A���`0 55f��/|
V�����f�m���]wa���*%#"���IM��}w��k4���`n��kkk���W�0�@ �$A��@��B��^]ǘ�f��f��1b�F�Amm-Ξ={�������}B��	GDD7���#��-����������:�n7�n7�^/B����_�,_�_�����a4��Q�:|ҵ���199����k�G++1^V���!��ѭt�R�\������- ��յ�����C @(���i풒�����ĵ�6���arrkkk׌4ԣ��idMN�����n��z�,_�g�X�|�����Cq��V��N����b4�RdB�����ɓas>� 
!�*$�d�w""�Y>���!�e`��� ���1??���e����������� ==6�6����PYY���i�k�/�u'�ϝ���Z""�}��z}�xyy9�nR(���\.������w�4�f3��Ү�c�F�-H��v;\.�5��\��܉���UJFDD��ta!�jk���f3���TH�<��籰����U��no�Oq��=##6���������裏��>|�A<�7)R!�*/-]�b� 77W�D���vcaa���W�.�����X�����j�r��$I�����s箝>�0��� �L��(����Ȳ������,E��M~>
!`2�������dff�l6ߢԉ�j�"77SSS׌/�l�hiA�����܉�(fu�݋��԰���b.>7����Ӊ��y,--���_������"1::
!��"���,X�Vnd*���(++C__�5�����c�TJFDD�ƂÎ�������(���n���`~~���7],�$byy��˘�� ���d��#��1��՘��[C��� �/]��:�������>�jjj����F�A�����ra~~>�� �2��ְ��v�E3�V�Պ��Ldgg#%%�����f�!;;333׌/:��G�ŋ*%#"��%qe�k���p:�W�.��Y��>�v���pe�Q@���â��eee�f�a~~��qg~>F��P�ӫR2""�Y<#�t|>���177������[�gȲ|�����i ��`��f��ϢU�퐀��*8�ΰ���F͹s�{�*%�d��Oi�G�ADDt=���w�}���:�MMM�h4*%�M^�������n˦�V111���	����h4r�:V����a_�泳Q��C���ѧ����b��ohh@��Kz����cjj
������Z8v;^��,���2���1::
���N���dz�>�KKK׌��<8x}6Q�//��}���333QQQ�B��������!ttt`rr+++a7��N�P�sss���,B��fs���c||<l�8����3g �	��(.�؁�={��sssY$�Y�������!\�t	��Ӫ�]\.FFF���g6�!IR�r�"�Պ�������gς�n�'�m_(���,��ى���[r�̍�X]]��������� ���l拔���j!�r��yA��@ ���*%�d�w""�I����5���հ�l*$�M������BOO\.|>�ڑ  �@ KKK���4RSS�� W��2W�� �ш�޾?IDD�d.;>�PXGԌ�TUU��*�,..������p:�Q9/�P(t�����ujjjR�n�^��<�����g Eqә��>%!��g?OZ�u��v�^��l���122���cii)�����z�p�\���*L&S�6��t�X\\�f�g4¼��uWiQ�%	�}�xM�k�%I��ݻ�a3�ߏ˗/�ҥK���rTlf}}�������lN�5�^����:����_7���r!��.�DD?xF�=�������VWWՎ��ˁ�333���GZZZ�7�`�X011��}.75g�Bŗ(��M���bΚɄν-a�F�*$�-�,cffCCCXYY������, �ǿ�dY^B�HB�AKo;    IDAT�Ȓe���F����E,..b`` ������O�B���l����mf���c��އ康a��(����`��% vC݆��y�u�A~ �B�iY�� V,!ܲ,� 0˲�*�HB�>^�Xo�q�������� JJJPXX���:�%%%�fܓ���={�p�JɈ�h�F+*0��6����.b
6��65o��0�% ˸�ײ
�+�0˲l��+�+y J ���i0������������RX�7�̉{���;l=�*/\��q""�m;v`�n/((��hT!Ql�z�W�.�� '��]Vpe��*�p�˲l`��+k� E n�@0���&''������R����L�T^^���ɰ�'��s �==1�R%mψ6������aLMM���w2�1 㸲��Q��eYH����z%C�e��@΍�!>����E~~>JKK�~���hPVV����k�}:�{�~G�`���T����Nǝw¯�š��<�:g*������ �n����4��dY>%IRO 蛛�9z���}���.
�U�,W	!��`[w�z<tvvbpp���(,,L�B���
�={��1Y�pn�~��ӟ������Õ����ʰ���L�4����9�u�܆E �eY~_��^I�z4���Ço�����fV0��$�J��B���m�g}>���0<<���"���$|�{qq1FFF�.�}jϜa�"�w��=acB�^���chh�����g[�% o�������/���o�ꫯ$I�BT!�eY�/��W�l��t��t"33IU��B����5���t�55�����э�%	��96��hPZZ�B�����088�����e&(��9!�;�,_�e�����~��_��M��~��Ƶ��*Y��$I��B�� ���YY�1==���i8TVV"�ۆ�F����k��v�֢��S�dDDt�xF���F?�N����P��w%I�
�B}Z�����Þ�M^}��t�FS-IRU(�pPтm���A���bllyyy���Lڛ�+/��ݾ��܌�>�!Fne��'|y��qG �����x�[(������I[�v����u#�N} ~	���$�}�ȑ�ە���_/ÕB�<�mld@ZZ������z'O�+�B!|���|s�����6z���bpǎ��;��E�D�m}}�������p����F��f;w�С�҂���F��� x��v�SRRPSS�����+f���/l|��7Ps݋zDD;&KJp�������Q__�B��499���^�|����4��e�-�V���Ç]�#�ѣG��c/�� <.��k;?'�@AA*++���nG�����q������׿	���Q]���o�{.l������*$�=�,cbb}}}۾mF1
���,�o���wo��}�~���N�B��%IzR����̇��"TTT$|����x���^N�OO���Rэ�Q�`0���!�Ha{��'�`�m��w������nG��|�;i^��Y��B<�l;?��hPQQ���⤭SG��Kx�o����O����܉�(�tܱ>�P�x}}=���UH��@ ���!\�|y�_N�~(���v���來��?'��2�����d<|�$�˅3
�?� {��
���h+n���ކ�u����v�ٳG�T�I�e���b```�Q{eY��V����ÇG�~��������{\��/x@��B�q8����ɴ����N0�����
�,ss�ܷ�͢1"���/~c�ujB���HIIQ)U��&k ~"I�����u��Ѩ_a�o}�2�$�x��mlu:����fmppa����(��U!ݨ���`����1�V�@�p�o�Y^^FWW������*��
���r�޾�[|o��^{m�$I/	!^�e�`��F#�������x�������H��c��OȻ|9�������(���DOO�ֶ�O�eyF�?��kmm=�x������_�'IҗeY�<�-�1&s�FY����ϵ��M�����_�&x[zS]��DD3B����b�����`�����ȥ�%\�pa;_| ���h���Ç{�m[���o�W������z����p8QJ;N�8��뺵�^|�կC�������"9�Ѓ�t�a�{��EFF�
�b���Ο?�����q�h�9r�(Dۖ�^{-S����,�_�i�v�F���jF)]tE*{�?B�Bww""RעÁ��\��������F�R�Y�1<<����-�|����j�ڿ?|���n��a�B�{ �l�|FFa4��N=���g���ɿ��R�v9
��?����"��֪�(vȲ�����vBB�������׾�F��=zT���z��Ǖ�H�r8hhhH�fH���8~�xؿ�<�V)mψ~/���s����B��333?S�y���~��F��sH� l��,**Buu5$i��	gtt���a����稺pA�D�lX�NDD1c��o=�L�xUUJK�lP�P._������6-=B��������W^�V���k�e
!�T�l�lII	�����e���)\�x1l��_�'O�����"���+_��`�f<==w�u�J�b���4:;;����e��eY���_~9�~���o�
���,�`�
����ر#����|8~�8��u������J���(���������.�����(6�|>\�t	.�k�G �?v��{��m��Z���o5���B<�Mn����hhh��n�b�������h�@O��? {<f�̈��o�{�kk�B`���	{[�v�����ŋXXX���. �t:+�bJ��o�B�%�G7{�h4���1�/^�����ke�������-׫DD������2Ο?��f��H��9r�����i=zT���~�_ʲ�{�g�����ԔT7$?~~�����,����x�/�f,p'"����?�2���|��hp�����ذ����ҥK�����1��	!������h7��W_M�j������/�b����)�;�m�eǏ����5�i��8��!����(ft�4�Ge666"77W�D�%
���ccc�>'��1�F�gG��R�����P?;;�.��� �"=g2��s�΄+ ���R������-2gfTHDDDJ�F#���)׽le����ҢR*�����ҥKa߻�3�?����:t(n�W~����_�e��H�!PZZ�����m(������{/�QDyg'���S)mŝ������.����hj
a/Y�\.\�x1���:S �����P��ݴo~�{eY~@�ũ(--Mص���2>� �"��3g��7UHDDD��3�+FGG��ۋP(�DqI�寴����h7����3�,�5��H�h�Z�ر999QL����~��?�����˗���Jrݙ@DD1k�n+n�����)n_]]ŉ'�*n� IҾ���O�� ��+�,������Ph��x�疖�p��	,..F3�j�(.�~�b�b��$����(�����FcRmbE���p�ԩ���Ǆ϶��?O�� p��!_{{�_�� ��x<8y��v��%%%���J���H=�a������'���1�>}z��v�wB�Pu[[���Sq; ���]<r�Ƚ�,� �}"Y�144�3g�lu�N�JIIAVVV����j�'QW5"�x���V�$��exxgΜ٬�=(���������Sq; ����r:�w
!� (���e���8�|�mr�"==���a���$ə(Q<J�3"Y�q��%twwoVܾ*��I���[q; �����F���W o��p�����NEEEE���I�R*E܉�(&��ޥ8�T���q�ԩ�\�eY�s���|�ȑ�q��_������3~��O�ު�?a@�ф��h��(v8��1�p��%l7��Z[[éS������\)��nwmkk�F1�-���|e���틒$=`D�P(��/btt4��n����U����������b2��PX�$���tuu�u�� �r�F��_~y.��n!�����= 5 �6�ssss�裏��)��ƽ������V���z��VdIB��ư���tX�V����g�B�sB�����?=|�p�M�Xw���Pkk�7�5 ~�9�ӹU�\SZ���֪�������gD�@ gϞ����f��<Զ����Ç����Ç=mmm��hv8���atttD�wJ$�A�E��5�� �f,p'""Յ4ԇ6eff"%	Csss8}��f�t}�,������G�M�V[������J��A�;w���QN}Z����a�#UU�4FD#z^�B //O�4���v�ԩSp�ݑqI��D[[���}-�C��ȑ#��h4;�?V��e���	���P�%�ш˵5*�!"��9
��~�ZPP�B����bppp�G��%ޛ|R[[�B[[۟!��x-���2N�<	���t���fCjjj�x�.�DD���2�-���d\�Ȳ�����(�G����fkk�h��Z[[�mmm��Iq�haa'O�ܬ9T�r80a�M;UHCDD[I�3"�ߏ3g���rEz$ ��v:�O���+	S�q�����yP���@�e���Ν;����|R~~~�P4�����T7\S�5�)l<62���q�̙����`04�����f�h9|���n?(������,���s��݄�T4�j��РB""�$���Ẻ��,Ń�d�����!����ȑ#Ǣ-*>�t�ȑC�,�9"\U9<<����('�="��
�������G�0!���S"�e.\��˗#=�𿵵�}���}5zɢ����_eYn�X ��xp��)��&�?�Ra���g�1����F�I�"�O
�B8{�,&&&"=��P[[ۗ>�xo�hoo���N �J����֢���B(��Nb�nW!E��gD^�'O����{� 0,�����~��ѣ�E����ѣ����� � �X�?;;�U�OB��l0��a�J7J�J,p'""�)�ѧ��;Z'�˅�/F��($��Ӷ������x%�٢�СC����?�e�y ^�gzzz6��MV�U�A��5�DD]#����ta���2^$n�gϞ�������<��ښ���J�ײ,�`N陱������Hr�� +Iz}<Q�j��	�Q#;;z�^�D���������b<������(Ǌ���������eY�'�y�׋ӧO'\�X~~������l@DK�F#�**��sss��hTH�Y�q���ͺ�Ȳ������h�RCkkk���n�S����5|��G���ĭ����l|DDc���(�̙3�����������z*�������F �%���4����s��E��IJgDY�rsUHCɂ�Dq&���o Rr�`��4l\qS'�,..���>Y������j�s��������XV�������l�SE�җ���l,�[�����V�v�[f��6l,%%���*�Q���:N�>��]��������ѣGQ�������, 0�4?<<�Y'ٸ��a/���G���`@0�
i(�W�ï�_�l�����"�/�r�$I���(D&�?��?Zokk{	���4��zq�̙�^X�;�f\��AH�q�/��� �Y(���� ���N�"��uwwcffFqNqV���ooo�r,�|�k_s;���dY�;����5�>}�@�l7�L&�l���: ��H)�$	^���)a$�Q(¹s簲���G��կFl�h^y�����{ ��4?77�Y�˄���0ψ�6�nQ�b�n�rf&33����UK:�:|�O|P�^h�~h�~��W`�����u~ֹ9�..A$�'%���Պ��|�����s�"m¹eY�\{{����Z[[���׿�_�Ѽ	���׌�ٳ*%��rss�����g����S��DU�$a�fÒ=�6ە���	Oj*�:=�:�5�5"�������C���.,ss���>7�OBެK	�k4*�������/�E���q������yt�u'�ﯪ�� h4��b!� IpߴY+)j�i�v�ĊE@fƞ8s�Λ��s�e�L��-Q��O^��S&/NB-�-��%J�$R"EI\�$@����"9`�-� U]���s�ϯɓ�6�������MNNR/'�����+tvv~�{���d�e �+X�9M��l����ב�hi��}o�c�R����/�+���H��	��iӭ�T
����Ih�����C��/�,�}}�I6���s�l��+�Fk�3g���ɓf/��L&������<A���3�<sJ� �I`�����`ժU�L�-++3L�pa�T�8aST��t!0\P����/��"F0�����!�i�<��žP,-G���}��Β���訍�E�]�&���|��Ǳc�p��Y���*���w��!+c�;w�L��;�v�:+��?�_�����r�J(�^+++C_ߵ����[V���6EŘ��χ�h�j?�`$����S��5횽O<-�'6��8����t��r	y�P�I��������2���O�.���===�qӐ�+������G?�[Ӵ��u���wwwC�4��:\�7��@t���^{�E6���1M�B讪BWm-��*1����O]nz��\�������qwu���YT�<���n�1aY�d������kC4�/�����7�Fq�ݝ���XVV��w�{�瞻=�J�@��ג�$8��k�"�����|(((0<,�li�wf���0�jk�U[��_LݸN��)W��`4�3i������/�S�0���-̦����Zn��c����&RB�on߾�﬎+�l۶��O~�;���^��~��a��~r:�S�����JK1� Ϥ�͘Ut!0XT��˵��uu����TZ�2-��?s%w�8y�Nq�;�]B�p6-�����u�5�ŋ�駟�������}?��L��v����?{�g�B�g�_������nGhWTT��c,q����YV�^g��`&��������Y��p����?�;0���gQz�,��G��,,�L��8�`�a�����`l��Յ�I/'��;::bVƔM.�۹k׮�?J}`` �F[[���̓��b!��N��p�;�
qM���J���EW����^3�q6W�!�HAӆ�y	^��ҳ�P~�$�Μ���,��q���>3�e��o��o��'��ر#�s��ǋ��� ����ٳg���yePVVfhp���Ų2�?oSTLfb����]��D ��[p�m	.�[[�	���a4<���K�����d ���7�k�"���.�)��u��\�x�ziJ��:;;_�:�l��϶뺾@^�k���X�f����gΜ!7�۽����e�JJp���[[1
Y��X�Q|�<}��Ç��c,����8W_w�Z �-��bSD�9r�N�:E���zggg�.k#�^�w�.K&�o0�v�����u���65�I&''��_�Ұ����h�-��bn�[^��mm��u��n�H�Pr�:��O>�7��f��MMx�ˏ�W�^-��g�MLL���F<�^������v��� �C���F�S��СC8���ꛘ�7���@I�l����@������6�[9�E��Ѝ������|��
��/Û��oX_�~������;＃$ݼ�����]n?�7ݳ�>�C]׿G��x�bTVVZҼؿ?z{��l(84�ǟ~���1[$<�ilı%m誫3���'o,��#G���!��>��f3�������?4{�/�o��ۗ�����?�����#��;�5!V�^�p8lGh�*�c�޽H��W��}k~���b2S�}n�N��`Lv)E���f�w痰o�&�]���"�eq�=UU�t�J�ilD��A��>x�,�ɩ�&�lj2�777�7�){Nq��)�9s�zI�u�������꘲�/�нe˖w |i���b1$	��<���8}:}N$A�����ݴ�P��Z��6m[o���J$�n�cyy8�%t��    IDATЀ�׬ƥ�Rx	���C��,�	�^/�m�=��_UU���B���ǥK�L'�
!vvtt�g�C�j{��}����R��
!�9)�H$0::��+L=.]�����k֓>/0-|3�qc���x����~|�~=z+ʿ�f%!0���3���x�j�35���[�Om؀���k�|>����;3���>�8ݰyV��;;;;MG���/��Ɩ-[
 �M������șí]�J����k֒���S��;4dST�m&�~|�b�m��~;������-�ssq���׬Aoy9�T�:7�1���6��j�z4]2������ӗB�����01͞={^���j ,K����hT��D]�ñ�99Xp��c|ށY�BM5�v+~�e���b8�Ӵ�LHz<�/)��%Kpt�RL������dl^�}>���>��MNNb��������\�x�w�q�������=��?�R�/	!��_���CEET� 'SU���K�Qb� ���MQ1�q�;c�(��8�ڊ׾�>[ގ! ̌�B8W_�OW��D0�hSSv��\�u�1P|�&l ���988����������V��/��©͛7B|���uhhyyy�6E7?TUE__��ȭ+*��1v������m�����zLf�gJW����8��O2�H�Eހe�:�Ѐ㭭�uY㙙�����oV����guLN�gϞ�-[���� ����(����L&WP��Bh��x�	��e�H8���ފ7z��j�pb�LtE�@4����p��	��)D.]�܅�+]��t��`jyy9���-2:z��ٕ���T궧�z��19��U�^	�� Z�_���Gyy��7_�~?Μ9c�_c�8��,���qh�Z���#8��h��x3Ѕ�Pa!N���x[ ���"�j�,�TU�ۼ	���Y���}��'�g����~kGG��c�v���|�E]�� ������@yy9�K���Oޚ��G�]�����C��[�WR���3�_�@��COu>Y���ː�ׇ���a19�Ѐ�]�G4��wTU}��~�����4{���w�}��(�# �9řH$066���2���?�Ἐߏ��>�I,��Ty�0�a	���\��׮��/5MC0D0D ��녪�W�O�T*�D"q�����166���1�n�JlO<��bɾ���l��B�o��o0\�^]]���f����d���3{�;::�fuLN�k׮?`h��47n���)���ԩS8r��5kJ*�o��ὁ�x�(#aذ����J����#\�WTU����な�H�RH&�W�/�]�U��ǑH$���3wpK���E~���onڄ�V,�f������o�' ����{���'_***ڸu�V>);�]�v�6����.��ڵk���gCT7g||��կ�w��g����17,*�q���05i6BC�(ʌ�����ռell���.����ڇ�C��ѝ͋K�e�ٷ�mX_�|9�ѨY����ON��u]����_���I��/�"7���1����R,]�Ԇ�2������HO�����X^>ܰG�.�������k��E��i�x<P��_��LMM]������P�%84��＋�����M��]uux���׬Y�p8lCD�����G}D��pgGG���(�w�.J�Rt]�L����/�#����oe������+�"b�'��p`���������z5o	���Wk-��BQ�R)�������FGG1>>���	�s���:j���7�DaڍM�͇77o�g�ۯY�u���ѣ8I��u�����O\���g�m�u} õx�/Fe�!�q���)�ݻ��=���E]�c�eǱ;�$rf�B�}�=�C!&"� �����O�%�I��������� �i�x�*]�+�x-� ��cl�����H�{��	���㪪n�:'�x����a�z<Ǒ#G�vy�,�i5)E�������/06I��_��֯��W!����|%??��'�MNN^�U̾'�1�͛�骕X���(=s�b`l6��kEEE6Db���ϛ5��7�Ϯ��㧻v�����뺎Çc�ڵYr�����i511q��ٺznpg�zq����x�����]Q��a"� //�'����cpp}}}���7ܸD*,�>�OV�Ć�_B�y��2�l}�aMQD"�O�C�u|��f�����g��O����?�������*���nTTT8>�F�����b��B<��eTJQph�|x�-�k��_�Y���PTT�������Y000�K�.ru�X~>��{�X�/���ӧo*�fC�Y4MC~~��X'�L��>3{y'7��n۶m�v��� �D�-y]]]���t�����"C���S>>b7Pž�6�Bu�u���w�����b�.t]�����}������	��M�p�q!����^��?l���3�9�Y�266F�$@O�RO<��S��>��۷x�g����׎=���b��6z�^���bxx���s�u���2N���y;��1���㍇���n�T��@�Ann.jkk��ڊ��:D�Q�B!x2pݓ�((,,Dee%jjj
��N �I�����z�Y��=��x�ioǅ��k�TUEss���nll�^��R�M�,ɑ��ݛڴiӫB�o!m�udd�H~���o;���CWW����M���1��b28[_���Wq��i�ɧBc�hmmEUU���Z&��=rssQ\\���TTT@�4�b1�����D0��K�`� ��s]�f��݈�hn�`X���C(K���o�x �!���ѱφ�i��Ϳ ���w,���s�&���8����Y�����pV�>�f��ᕯ~���rDQ��������T������d���i���EII	,X���2h�����Y7`�ssqd�RL�B(>{���2��/݁���@"��tS�ҝ8q===�K�z<�o�ٳ��v\��^z��-[�ܟ�������wo:�׋��ͺB���
�?��م���խ8��:��xB]��TWW#�\��~���Y����:�������u�X �cK�`(R��s�M�9f6?޹�n����b�����5�;���>ú��?���ݶw�^���:��������;�_Bee��s�ǃ�g��ԅ@��_2��a�FĽ^|p����\��Ɯ�TUU����-BII	���]硾�!�������������pBLLL 5�0F!�[^�cK� 0>���ޛ���t�"|�=��>����tvv���x���_|����_���eR����Pr�ed�+�����C�;�@��LYq�;cpt�R�򵯢��x�?��xP]]���444 g��}6�� 77��娬������������.[��?�N�U�,���zF��QQQaSD���a@��?xꩧ������_ڼy�i!ė�_v��k���1É�)�����l�⚆7�܏_�u�f9
�P__���6TTT 
Yr�H�4D"TWW�����`ll��!�WR��˖"<��E~�q'��qv�SQ�hii���zNq��Qrz��������?��c���S<��> O ��Kupp��wu�µӨ^/�>����o�`l&1�{~�o��Yn����CCCZ[[Q^^�`0h�s���E$AMM���Fg�<m�5r�yi���*�ix��{�?�����͒N311��R�	� �ھ};?��/�����߿@���x<UUQPP`Sd7��񠧧Si��ީ�����Iz<x��{���{1��g�~?������RPP���j_����,6P\�#���BA/7��̚��ޗ�dX_�`����ddd�1�� ��~���'����U���B�; \3Akjj
^�ב���|8w�aЄtU�nSTL&+*��o|gg" �@YY�����Ԅ��"�f��d��@ %%%���A0D,Cl�	�	��-BOe*N��6�ÐX�li�����Ο?o<���TU���|�]�@�����J5�QUUtuu]��RUT�<�P�p$�n7�3v�^/~u��8p�-3N��4���X�d	���-y 0��x�5�~?���̧w��8W_���'Ỏ��)E����k��TUUI�	���M^�$�8t����޻w/?�ы/�xx������e:55��#տ�T*e�H��A���<����@q/}��8_[;����Css3���2r5�����A4�:ugddĴ�=�i8�҂�?��S��D8˘�W��@ɵX��0���m��Z###8|�0�R�����⋳�wϮ��/to޼�H�f�z*�B"�@�,�����#s��(Jk|gl.z����7���U3O���W'����ٚ���~_=�=::j��$�^|~y�k�3<P�ݰ��*]�԰�h�"[k���СC�a]������m����wE��k�0]��©�g�^/Z�{Ϧ���#����p����9,
���	�/FAA�%Î��|>D�QTUUAQ����6�'=�ln�x0��S���4=��9誫ŉ��zss�����6������|݆�m�޽��-[�� �<�����M�###I�]]W48`SDL
B��ڵ���È��X�(
***�l�2TVV"�6X�� ���JD"LNN�M� ����6D���78ha�Lf�^��b�����$���O��R�'�|��|g����ۼy�y!�c�;�ƙ�|>N�>mx����Giڭ4�݌�����KJ�'���K�L����hllĭ�ފ�����B���6l��%K���c�g{�����N7-�0B&���R$�σ��BQ>�'*躮w�Ν3�a�L���	�p���ɓ�×c���B�����t��/�?}��,*2�3�P+V���u�PRR�U�^�������PWW7ㄳëV�_~�71R �Af���*ÚL�fs��q�9S����SO�d��L&�=����]]]w��s��CN���\�� !ph��/~�g�����ŪU��f�D�Q�]NN���p뭷����4�҅��7��o~㹹�al6=U�\E�4�ɞndd��D�c�d�?[�,������ד�$N�<iCD�C��#��s���筋�O|}���������6l@YYYV�Y4MCCCn��6����Xg�l�r��o��"#d2�r��?�������a����h4���xd�}����Y�z"�0�@��>i_Iɬ7�1ff2�+_݊_�u'R&��BTUU��[o��ŋ�n�p$�Z��>?
��o|�o����0�u{����9s�p� !���'�|ۆ������?�������:���^��="�a����8�Ѐ������+�)%%%ظq#jkk�z���+�6l؀��Z�bk����{mXoq�LF=�À��R]C���cv=����x��xd��OB�I���Ԕ�
$'���!�H�4Ʈ�.޾��y��H��!W�_�E34�gMӰp�B�_��3�_����O��6.^���؍���(q��[�GGG��1]�������!Icǎ� ~����#Ȩ�>մ��lR��7؂w���<�ǃ��f�[��,o��z�hjjºu�f��议�Ϟ�6���Q�9�E��0???�)3�����z*�ھc��{�٬��8����ՅI��i�|��؍��������6*����zlذ!�og�x<hhh�ƍg�	�������6.��+��E�:�����(OnݺU�i=6�u�����Ϝ9c~s�P�	]Qp��̆h�Ӎ��~��p��������b���hii������0֬Y���V������-��c�"��=:,����bL�=�d2I��
�/�L����HGQ�� N8qh&���'������9:��?��r�4�EC�+�l�2GM�x<hllĆ̓2!��w�����?F�&PM/�m8q�Z��u��:)��G .���<y��6�T�7��Y�T{~�W�2�3EEE�n�F�`+W��ҥKM��~?^��7p�����L̦�T��ɉ'��S!��w�����ߤ�����n������9�7���橨lN~�/�ؒ%������jG�.���W7_͆��Bx�~�]o��nr��̹��< ���SO�b��ٱcG,�J����T*��I�>����6����͛q`��?SPP�6�����a�l�����gy�^���|>������"��ݸ�ǃK��2�.���f�����'�|��xd���9�������H$p��;BʈP(Dֽ{�y��Q_I��o����^���lTQQ�[n�3::�h^���1��M�,{]4yft��e&]]]��v ��o�y۶m�L����ׇ����[�D}&b~����36W����Z�{x����h4�)�3	�X�z5jkkM���kVc�C���ͦ��4 ����K�0<<lX�u�/:;;�mI:۶m������I�;g��X�u������L�5�l݊�/&_B`ѢEX�bE�]39���X�~��oG\���[q����Ș,zˍ������)6�011��nc�"�x����B�����W�Z*�r�����^�I�]�XN^���qf�B�uEQ��҂e˖9�;����֭Cnn.���c��Lc�ő1��D#>�]�=�����Xd�����B�C���Ν3��v�s�SP��J�*^}�Q|���|]���z�Z�
�@���2����֭3�Iz<��c��H�2�#c��/)!oj�i_(���������Xd����0RN�>�dҹ���KD��13jj�·~� �z0Ě5kPSS�!�i����V,Y���p��*���o� vC�=�@ `z(�if�Q�WU��ju<�J&�b��I��H�p��-��$�b�:}�~޽�N�!�|�r�i�Nr=�=��.�k�>
��,�M�|��3��W<9��d�����c�c�Y"�x�a��'���>IU�PQ�Ѱl��x����\}�zNNV�^�X�<���cv(/�(����8��fqdL��%�5�7]�;}�47�Y���c����]]]�ڄ��|��e}��6DÜ&���o|�t�n ��5kP%ɔ�@ ��kע�d�^���/��Ns�;��ѨaM!Ume���I\�p�z�5>��9BDΗH$p��Y"��s1P\��e�Y���ʗq���\����b�
4448�9l����Z�
uuu���(�����l�r�cN�_l�]TU5= �tcccf�9�����S��նm�� ����x<���."�*w�:�^j����_3�\^^^>�|�)++�񿧿�/|�70���������L5���nLNNR/��˃Y�ر��/��188hGH��*B�A���]X�pg*c���ex�;��TUŊ+f�x�T�h�֭3�<r�i޺�^��bN�WBo QI�MNN���xc����m�6�ދ��v��1����ccc�!����R�صtE�k�<��tX^^�#���͕CyK�.�7����؂��������.K�&���5���}��׬�GfB]�u�����ǎ�n����%�MRU�|�L&�D"�]�y��h'S���hii!s�����GA7_?�f�_j�U�~���:����&�	!7���SXX�� ����?ކh2��U�|>�JԜ�����zB(�ڵkQX(�
!.\�e˖A��	���״�13T�%
Iq8�2����27H$?`�fwr�B헎��!��Y�5�KJ��[��x�����&�s㕉�Q� 8 E"�ׯ}q�ȬG,�i���wr8��:�]��'����\%��P�D�Q����,�,\�77o"r5M�ʕ+�+bN����f��M��V,���n�8*�dDc������u�.��������HOU����I���� ?�����6��"zs1�`ժU�\�G)--�ʕ+�!
�)E��_~�t:,c�&��V���fz{{15e�Y�?�:7�F���� �Ӧ�Q�.^���B`�C���V���bin�3SUU�e˖���	��|u+��<�    IDAT��& Ʈ��ge@1y����e�֭[����Y�����c���}68_a3y��/���F���|�^����H���X�j��}1d�t��72F nʓ5w�u�,w��������nǎ1 �f���!������3�D-�8�$#���v!/^,���+TUE{{;*++��/����[���d��l~L�� �Y��b�9��O����9��?�utt� �O�����H�R6D�y��ɡ#�n7�36��x�G�"&U\�ZZ�I��׋իW#�����|־�⨘S�>�d��۷o���X�`۶m��/���4p"򁀧��i��z������bŊd�lfj�Ox<��֯`����Ș�P�
 W�b�$�����cu,n�u��$��I_0�4+QM	��Kܜ�n�;wߍ�--�k��߲���O�iS>���a��=��P��d����������u]7\��2�����X��I���4M��h��>G���5kph�Z򵢢"��oل�a�Z�����T�>�(�i�]!�z�����3=�.�G� bN�]�~?��8PRjC4�	b~?^���'jt��bٲe���2����|M~�e��Q1'2�#��p������(8W�?�O�B<Goo��d�:
�E���Θ��ߏW}	����a�ʕ�L����b����o�{/�J����n��0 �����0��
௭��MR�����c��'u�/���Á��ע�(�,YB_)-���<�X��l������c��6+*W1k��I<�ŋ뺮������	BrUUy���ڄ�������3v�N�����U�keeeX�x1q���"�����|m<��?�E��>qM�h~�a]��J:�	�	 ���P\�w~�w�u]1}����|���멪�{w~�|��� ���8�wEnn.V�\I6�O�|x��G�pA�?�9�bDM�e��xNN�?X�[l߾����34�e�`�x��@�YA����
�X�d	�]v��������k��Z����GĜ����4M��L�>���8hu,n���K �+&y�����G�2�wH��_>�c�f�����+���m�^W�ܩ��ǃW{�����醉C�2��0 	!��Z��$�� �������8T!s,/��]���D(�_=� t�	,cɒ%�j�"//˗/'�.����w�eCT�IF򍹊������!*��W6��۶m��{��N�c�� �{3Z �mglnF

��7�����Օ�K$�ҥK���5�8p}����h8 ���R[I���cX�u�����n�q!9L���P~q��1B�����rr����5���\�Ci��B���D������sjO���N�����|�'��H,3t]7�.fC�����5K��Z�3���k---�kn��������k��s7nd3o��%o1�mB�>�<ڶm[�ߥ�_�t	�d҆�2+''�<>�7��q_%���ph�j�&EA{{;9��-4MÊ+�Ӊ�xk�&�bN�TU�Y��l��|�����Pr�;v� ���u�n����*S��qI�pe�GW���#*3m<�E$A[[�(vx�
�nZdCT�)F��F74���n�|��'�Y����7�kCCCH$v�3gB���7^�4IUū�>B����wm�����hii!_;�a�/X`m@,�Q�� Hy����&&��!��,����^0��>00`C47��=RM�ń�=Hސ����b�
r��[��a�:ˑe��y[�Q1�%�,��H����� ��9w��'�O�������ͣj���g��[oy���3.Dee��e���VӃ�^{�!�]�۱�Q{D���芢���y�J��`*��ࠡ��HT�2���,,3ܻsĘ��h��A����z'������e��b�筋q|I�Q1'��''��@�L&͒�W��ōt]�y���F�Ә}>�yҘ�\�j�W,z<����z�����R���_�|��K:�ݼQb����l.]�dX�u�!�3�rvUUy���j ���8Wa����nå�2ú��E{{;9��m*++�+�uE�އBL� vc��G^�W��f����ju,n�u��) {�ם�$F����s�ņ˗���uUU���.e#�\����|��M�����q�H�:�I�2566�K�cq����I_w� $*w�ɛ��;%<���#H����R����UvB`�ҥ�o�PQ޹�o�a4�/Y� �<�ܶm��cq�����6}������k͆t06W����tB����#��,--u�)������hr�ջwމ���؈�U�23��d��kV��F��� ���ԍ��4M��t2�<1�����Í��ZZZ�)�dBCCy81���ݻ�!"���+��$���I�Ca�[�=�䓟 8����&��ι
��`4�Ckא�-^��ƦY�h򈛚�C!|p���Ĳ5�H�g ���C���wz��ō��\�I��LG~F���+�D0��M~g-Z��}���֢��Ȱ�z����$�hT�"Þ�$wy�?���ձ��!w�a�.�Q���ǃ�y?����c�8�����x�b"�N��a�ҥ&��,E��0��{DT�"��~lݺ5	���u'�̈́>�Ǉ�Yfp�;c�]�����A��`��'�A�xe�Q���i�S�L���۷�:7zꩧ� L_�偀ڈ���w�=�ՉUUU(#&���K�,!'�޺�,�>(�զ|>rB��McW�MG�z�{������/8���ʷͰ+��{9H�����)���(X�t)�����-/�!*�md�hMG�RM�l~$�Iä|]�y}���x|]6~}=����UUU6D���hkk#wN76�S��ɘ����ƹ�u���%�LbhhȎpn�Y-r�'�2 ��h�:ú�(X�l������T�"޺3Y�b���0E��p8oll�X̰�J�8W���0����ɤ�d������K��e1��}�����(~��������?moǥrn�cךk�2�����B獆p.�@�Tˉ�����w����T� -ZdCD����T�w߽��̽̾[e�.l�{y���ZG�uC3::�T�pAMV�r�I�U���Z�eyyy��"3��t!��{����7)qme�X,Fn�&�I�x�Hgg�'���A'�ZTU%>OC6DòIwu5����g�%����5}o޾�$x/���j-24��'o9���:����h����]V�z���i�b ��}�!I��644��±/�,P���G��d�
"b�j2D?#�Pw1y�Oz<�_Z�[�R)�>����U�Q��	ɇ�1�p�;c����˵���<yΔ�ih$�tE��w�mCD,�ňϘ,�G�ƌ7L��kBq-!Ļ�k��~2u�h�\GW�s�������M����Wh���m��e+*W��a�pc?EQy����#�9��b~?7�\����w�iXB����ܬg_���D��t�[^��یMx�]&��0�{���~5M��"B]ax����	�w	,���� r���&i��󡨨�������0>^�Ɔ�X6sK�b����4�}�cq�m۶�H_wb�"��k-�/�zgp��ΰ��o��Qss3Y���m�m>̝̞e�#2�=<�m�6�bw����O@�sb����[R����Ę5���1|�$x�}�a����D��PQQA�x����"bيjȕa"j"����$���cq3!���vRc�L���oºΉ�f�����d�6�VKK�Ƀ��!ɇ�eT��lCI&f�M��p�x<~��J��1T����C.wd�R�S�***x��u0;p`�z><�r�W7�o۶�ձ��!'t�ƫف<�^g���G4i����Z�-"�-|�f�4 ��qy���m۶9��^��.T�e�s��p�zr�	�.
�� �|>|�j����D$BHq���k�u���,ty����u�����`����r��(�,Z�H�"�|hjj"�>�e�ѰlEm��3K8���Z���G��םZ����2Ɠ:�E|�~�a���`ѢE6�<~��������\[�Ć�X6��[=�ԛ�d�X̰�y��v��p&}�)y�YNϓ��+�(8�n�a��8f������*��PQN55��
B�����xYC�&1����G�u!���m��yrrr���`X����Y{��l4��!E��܅�����܅��L�]�{���AQ'(++#�2���:�9�^�� ���8W���*ә�q��n7�3כ�������@ ���2"r���\���ֻ, ��;QS�$��)�i�I�cq���� Υ���@@n��iWW9�؈��a����,�1Zmm-���Ѻ�H�ݙ��zo&ccc�uݰNM�`��P�5�V��L�spӘkom�h8lX_�`��߫�T__ONF=�q ������K�2LK��Y��'�I����V�t�kj�SYiX���@0�!"g���&��[����Ml��n��܅�#�{>99�D"aG,7�|Ĺ���Σ�1���A]]�a}���g˗��6�Ğ��,3�zϹ���lp7����3,����ާ+W F����8�g%�a  �]cq$,[MI�Y�4&�z'�m��:C3�7]�Q�$�.PEAMM��8������6���q�'�1 q��U�FL���d4���X�N�uC311aG(sf֜0E|��;P��=9����z����0�����\��f&����V�*G�x��4�|ϩ��Y[�\ŵ�_oXB�7�1s��`�����P��Z��e��ɤv�]�|1{ϝ�ODNp���v}.�����SJKK�sRQQA�:�vBb�3����8��$��*K�R�������$|<���<�uf�wt��ZNN���m���rssQ\\lX?�p!O�c ������n�0p��8 �/}���9�)DA%)��4�>CEE�h2U����]MM��s��͆hX�I���V�;X&&y��֭[������<����#� �����l�.VT`0j�y���J�F��V[[K~���,&��I^"c�b�,ϵ�uuu����q��>')�.��x(�s��� vc*++���ҥ6DòMR����8�NUU2wqJ}e:�90)��*�1G��5 >�7wfã�C!t�td��~�ι���J*�"oZv:w�/�g��E��.VT`��аn�y�fG=D�'x**]x���i��7bu �����R��\�X�q�O�q����c��j1
��&)����LL~'9�������I�t��s��K���̦{�ٙa8��ȷ:�P��U z�����d�k�Ν	 ���N����x�Օ���A'�=p���x<򶼞�
���6DĲ	5H �3w���9w�^,#�sYr��3��RU�hi1�G�Q�������;N��1wI[d�[��k�ƹ��TU�&WIG�]8wa7��w�ըMW!���l�F�p!�9���d���dx �
�B~��p������>&!p�u�a9������*���)E��>��v�a<r���4Psc*tRC�8���6lnR�Jp�F��r3����0��5����S�dSH�y�o`*����Z���]�SP���Byyy� v�\勚���'ȗ�$	r�&�.�۱cG��VB'�.��`����نL��P���x<����O/jD��!"�-��Y���~��*3; 餽 3�$�����鑱90;�Z\\�Wf�$j��Ŋ
G"6Dò	���P������O͘6��TT靯��(1��ݜ`0���<���V�&7sj:���L�&��!�pt�����K�1�t��������~��̾We�.{:���ͦ\�y'E���$&�g���Ri)��Q�:�*7���#B��ok�(]άW�Z���"�.�q� �+8waWP�������Ȇh�A�KhN56��n�g�����:�SŰ8�Β�� ����oa�nPwe%&��A.d޼��2�)F!p�'��^�Hhd=�*���!�B�����0`�9���;��XHSU���6D#����2�@s]5�*2/gB5��<����'m��SQ�C#Ln��4MC�h$csCի�/X�XN��0��&y����̞��b)j-�A�����a�o���=*,$0���'$[�J��uEQ8w����9Iq��uR����z�zii��u����a'��_W��Yd����3�v��I'1l>��
��d����|q��0c7��o�fFNN�Ds؅��e��tnC$�E=��n|"f�Na)�$;��*�����c��F��wm7��k�=g�č߫f���0�T�<��<���Z�ϊǁ���P������5�؁�]tEA7�.��&�g@�������F�Z�ئ&8Wq���faa!�^����,�;O��1�0��a_h:�ƷT*Ź�=��]���y���by9�fX硍�A�����d�3s�Q�����o�Ν���b�D����d��#�܅�<��b�u�h�.((�M�),,4�uWU��i.G5�:qjB:�d3duH�R��kN,\�3��x��]j�~?����|�df�|>���2�����Ur��p�=���cȦ�x܆H�]F
��M(��dF0D1��sw1�^�a�u:EQ�Oɤ1�g�N�uG�(WP��'����$4++뜫d���A~~�a���[r��$�]lcxߝ�4F�.\gq��EUU�7����2��oQv-j�H����^�F��Cal~��J�N����="6_����RB��K�ƤXvc��pB��[a, 3�����pi�1̉��t��DI&!$��0s�j�M�HĆh�D����jm��eY��3�<&{8��o���5kBX���܅��\�쐳��gyUU���~�
r�q��WOe%9���,�C��jj��T�rK*y8���p�b�ݻwk |��N�]��g8wq��M(�H��6fH8&���.�<��~��%8W�X"� ��d�i�8wa��J=��H�*o�fN^^�0p��چhX��6�$~ ��0���N}N�a@~����~�~?�l�)���x(�a��v-Yo��	�1���y�����.�5��%77q�6�1�`��h&<l�-T�f\���HMg����WB���LǇ�Xwu�aM�4�B�ӑ)�SPKJl��e�4�_�@��'�[O�����<�]�$���H��y�#�@������o�s+Y��̞��~7��QE�w����7�3W,2�4MCn.�vg�ٔ���ѰlA]�+����|%���݉��t�0�NT���*(( '�D9_q+j�H�\e&&E���;w:���<�/~�5�n:0kf`r,4��ƃ2�|?��`���39�=�x��Z�Cwww���)9�t���� �oV`7&�M�č���rk-&{9w�X"� �s'�&s�r���|$�����2����s�ŵ�="j.3�K�?v�Q�-EQ�\��:�]ؼ�w�JCD1���3�zO����ը	�2<�|��!����0[,L_��ɱ#���B�;�
O�,M����A�W\��n��R���w�STTTgu,̹y�YsOs!0Th����%��~?�Tʵ�p�T�7P�hC(��i��;%G��������s��R�f�ab�s�zȱ/���mT�s��R)�=�j��.A��<H�]��!����ȋ�i��E��!f7�{V�����5�mư'���:�ƒ�t�]Xp�;s�A�D���n�p5\X8���q�>���ht�š��O�� �;�d(���hs!SfqM�QT���s���S�A������L̾W��,����)�������� �����v�~5DԹ���d��0��I̤V�Mb�3�'�Ǒ��T��q����`��Y����=9�f5l��.��s�b1�=��|��>�Mb�2@�~���Hqsu6!kWB`�o%t%��-C�"� s��^*�r�>�L�ܹ��n7�3W�&�����m��Ԭa����4��%(�pcXv]"����}jjʰ杊�	�ʐɁ0�=g���7^��K�*SSSROqWU���p#    IDATl��1�я~�P���f9�6i�L19Qu�s�����χ�3�ә|p~b=�{��$��h\[q���|$�f0�U2�lp'��3w���P�fs��G�]�'M�B}N�)�全�G���%�� �ǵw�y���,YC�w����c26W���\'��`��q��#ۘ��|�սB�Æ�I	�^<7�e��c��av�ib1�k`dĆH�UF��J!�~��ȍ�W����Cp��ݪ뺔��Q��F�Z^������)ϩTN/R)���l���a� lX�4^��9�I��a����$j+�3�ә�<���V��r�4�Q�J������L����9��u�U�JI��5�˰/��$w��|�,�5x�)��tT��}!W)06�s�yf{�Ü��R`�Xs�e���=B�>�Ũ�ܩ��tf�=���L�w�:S9>r"�Is*�	����]��^���Ȳ	k�t��:7K�R+��rrr�(�Ow��?Hm����z���*�9T���3w�� 97^���]���l�$�I���z�g�?6FN�cr��{6��2?4M3�M�pό�P�&&&l�d~�p[�(�2Զ����:�V\.N<���
��cC4r�r���!%A�����"c����Q��b�V��V�?��
`Y��s�d2I�>0�]29M�S��2?��5NԺ��̞e�i1�jz�g��4ؼx��䥯;eh&T~�ŠI��a��js���N���9?��5��	nn$N�NLLHq�S^�!�;t]�nT�!������oG(GNp'>OLS��+�*�z_t�xu%��8ِ+C�r&�����ҧ�~��a����A��a�{V�1�������i��O�wjj��Mb999�a�T*u����O?ݨ�ze��I,��])�Mb�'�q�2?��W�s��K&��B!�ΘL&��l~���.`������3µw�}"�P����S���r�} Mq�ձ���(��P��\%y�ߚ�2��6��Ѹ�9?��uJ���
����S�����l׮]MV��F�w��1U,1^��D�4�>	bZ�*�,�8�<��'R)����2/gRXH��+B�۬���nO_pRC}F�nD`r�nj�M��An�z��m�LN2ߎ��䷐�-����kB�XV3m�|�5��x�������u1w�[d�]����B�n}4�(�!wQU���%ۙ�.\kq�0;���iaW(�r$�#���%	p�b)C�{^^�Ϧ��\sa����u��B&����BOp�B�[�^dx (,,� 
�i�,���m �'5����bH'�yʘ���j�,�ҹ����� �~?�7�Y��[�&}���AV"�s�m3�'6�x�u~P�.�+���r���v�e���r���<�&�lG�*"������D5(q�e~���f{sL~T�j����~�Ɵ����k$X�Q�K8����:����A��p3G�Qp�e~P�8<�ݽ�!s��]�\%�Jq?�t]p����P��ga��l����4)�;���	����ƅc��BHz�������7�!�!7�+}���!�KF�M��	�r��8W���Ÿ�ݵ�/gBф����$�IC���Ts5a��+A�Zx�u~p�#�͡x<�d2iC4��d�OB�!�y�s�N�ÎN�x��y��8y�<�S�h��:��0�<յ�:�����ɜ���V��6?��� 6��;5w�>#�$�>	���k-���������Y���AB��ݻw���<��3� ���N�UґC��&c7��7�ut�pj�5s/%��|ܰ>N�9�|�~�O~�9��,�s�N���[�ם4�t&��C�:��4����Ƶ���e�,6�I���[iu,n#�x<}-77�1�Qu]'�|�1�q���a<@�|% '�x�u�cq����{ 6����J}>�n�d��ޛs/��s*������!�.����= ����܅��:��7�������s���.2�� P���W���m�|�i��fB}F�j���7�3��T~_�amD�Ħ���Z�MMM��Y攖��#�(I_�F`i��.;wp���1��<1�Ut]�vQQY�O&��aC8��k׮: �In&yeV%?�g�1����� oǓ�����MB����O�q�=K�R)C�i�c�Ć�f��K��0Ƙ����us!���P�_޽{����e���|>��e'�>�}�g�1�XfQum����A�oY��<���*��^XX(���͒���L�w�c�*�hX�x�(??�쁀��Q*�2<py<iܩM�"a�1w�߱�dRʩ��y�^�S���ݻ�1J܁t]� �ɂ��r��1Ԧ��J!��kC4�1&?O"A6���$ eeeԲW����ɏ~��< �����BQ���D}>���c����"0:fX�5w1y��K$Y�[����y	�������9�Z�urߔs��F�Ec?�L{D&���ݻw7Y�[�����Pન��!�̣�Y���~+c7�H�c�E%1��xL�=��s���v�ޝ���w��q_��g
ڠ���b��bUw;�]g�8v\r7��or��^�nVY���� ���b*V�z#%Q"	��D!  0�e ����?H0��΀E��7���y��y�3��'�3��}��t-,,��kW@}П�x(BDD�#kxP�K�4��,7~��\⁔R!~7<�j�*$''���MQ�U2GF`Wt� "��:[�j�Xff�������V��n�� t]f#�������.��(Z "��O{���l$&&��ܻ��@ � ��Xݻ��� ��ؔ5�"1""#�R�Ye�����դ+5lT��H��@���	ِ�������<
�B�����LH)��ѹăP(�� t`�zp.`nnN�4!"�����G���.n��˥������7kB��	�X����5 k�㱶�Q>��+�JRu��^%�ߍ����ۍ���.=�ӝa���`ժUf���E���NbDD��V�Z���"����������.M�vx<--iii&d��E��7�IyDDFH��G���.n��KRRR�������;�G�v�K�Fx<??��y�Bˇ�DDd�U�ð):X�"699YYY�������b�Z)���եH)uw���1{�.��U1-�lŤ�<�[��fC~~�j�^�-?���_1���MS���he��z���caa��lV^��bB���y��/ ����ɕTg+)��H��5!"���j|4;;͢��"L���B��1:��4�w ���#�oT�,�##p�&dCD�T��V�#���dNJJʟ���	!����xqq�	٬չK6�h�����e�12��[�� ���T�$MӾct.V�
 /<�z�j�Y���Ĺ9�&��Ɖ�h�����p�W�f��n�' ��)��G���y]���VV�K"��W���#�m������|�LJ�|�WZZjF:�By���xDD�R��H)133cB6+/---R���x<�F�cU���v �G�#���T�<g!"2��'� !AWs!�_�۷/ф�,�?�A>�?����[�ac ����Źw���w""2��0s�B�yyyp��ӛ����l��}��%�l���'$$���Č�V;��Cu����-��J���, 3��{�f�s�"��_!"ZY)SSHRt����J���*UX���q�ݟB�
�#))Ɍ����lE5����VN�ovE��8ܻ8 ����X����o X/--���W�R*_d򜅈�H�C�?w�tGd��Q^^�Z*r:����l�+~@rx<��:sxGDˋ�DDd�E����	ˌ�B��Rل#UQcp:��t:�\J��d///��n7#�1:��v�30`B&DD�%ҟ��?��(R��f�g�s�"����Rʏ�����bFJ7mddDsMN"٢]������l��{���t��䨖�X[[���|�����!����x,>�����Ǭ�1H6�V��e���x\d�Kvv6222TK_�z�����j~��'	!�_�`/&LMM)'���DD�rr��Zi�RVV�|&���}�������<���R�o��SSS���oFJ+B�{"��Gڸu���X�NDD�+<wN�B7!���@I��׻Ǆ�,��v�J)�6<�p8bzdv�����������?DD��\��H��UżV��LJy����-R����� ��c�xLuxY�����+P�y;66�P(dB6ƈ�w�MJYWSS�0:+����3 [��EEEHN�5�����(��1>"�8Wt�[����d��SJ�R
����ٿ���PRR���2Z�s��!��τl���kbic��+���v�����
�?������A���BXg�ڻ��,��'������=8�D�_�ҋ�%��ۤ��������$��������a��l�d[(���^�!"�?ŊEVګ\˚5k�q)�C��q�����U� 55Մ�n������u�n�!"�CŊ?oC�&&��!)++YYY���rKnn�7MH��^o1����g[1C��B���;����n],(�WZE^^�ӕG(wz<��7:�����B�Ux��p�d�+��.�}��Ttu'"��U�ػX�h����.� ��v�o1:�ؿ� |><�r�PXXhBF+#*�!��w�>
��ᄔ_텱����"dff����������X����,�_�'''���IU�{�� ]݉�h�uu�b������3!�edd���H�Th�������ڍB����v;֭[gFJI��;/����38�D��C��gB6�ٸq��ӕ�~�a�慖
��///WN'�%��J1������6M�ŭ�	U���:���A�ǳʄ�b��iH
�WVV"11ф����R���,DD�P�s[���tb�ڵ�% �6޸|�e���E�i_���ƔӘxGDˍ�)��I�&d�2�/^����6:�X��z� �@�V]]��:�)%���tq�Kq""Z���)G�Y���J6lPv�B|���~҄�b֏��P(�( ݜ�5k� )Iw/�T��飣pMN��Q��
g+Vk��rEz��n�������RLs�ݿ-��Rx<)))滷���`^����f��L���_���%33%%%��< ?�RZ��� �� >w�\X�z�	-���	h�G ,#"2Gaww\����(�6
!����}ׄ�b���r�mJ


���mBF+G��O��F��~����S	FDD1E�5Rw�X������RՒK��z(��bQMM�MJ� �̦��|��暐�ʙ��B@1r����DD�I��A�����*KY�{�MJ�SvI�~~��� ������b�V�!��{""C��]"�XIeee��a���������*��]-���H��p�ҲR�B!��J�1T��GGG���d�ڵ� >W[[�m��U�������6n��M�Tg�΅�����ʋ�;"!�R��k<��F���n���q�ݎ6��
S��vu+�}���'"�����!ezZ��(�k�F�xݚ���ODW����� �[�ˀ���=D~_�	��/U�������JJJ����Z�c����v�����ט��fff���u�bE'a""Z9��X�l�J����xRʿs����R̩��KB�p�����!//τ�����.�30�EWw""2�j�i�r���8�N�_�^�&�������N)��۷/�f��@b�Zaa!���L�jy�b�}�Y��*Q4��;����HM� �z��H��jkk7
!���֮]��D�&����ajjJ����i�:���.\���Á-[�(����_����"p�ݟ�R��jm�ƍ�Ĵ��]����`Єl�����uaa�r:�"��֭[#u����}��b����7	!�U�VQQ��u1!%
86���P�|#���?��&//%%%�%��1�ۭ��%@J)4M��9|-11�6m2!����Ċ�W!"2U^?���F�w)..F~~�j)1
�b߾}�S��jjjl��� �	_KNN���1����abbB/T�M�q��hݺuHMMU-I)���S��!����~f(z�&999(++3!��i���=C�Q�����LSq�M�����,TVV*ׄ�Z[[��S�	�����O�������Ȅ�V���4�
�[ZMȆ�(�wu);<����RRR�*t�+����F�+���Wb��~ =|-++k���ec��1^O/�ggMȆ�(�I��6�����0�q�@���iii��B!��0�V[[�? �~x\�-[� !!������࠲�F9�V��Le�4��=��[��ʦM�����Z�����я~���Ļ���� |1<�ؔ���z�Hg���>'���v;�m��]9���P(����֙�y衇���1|-!!�7o��)�ע�=�30�TŃ=�����iJ�v�� ���Bvv�j�
���z�w�S4s��k4M{��pjj�%�r��
�D��""ZY�`�g�u�x�x�RAAA�.�B�/�������ߟ�p8^�k͑����[������4ffft��f�!"���]L�4�|>�1��f[��u���y�ۭl?�<�7���Z[��*�\�pAKC�E���bIe�~�b��G�N'n���y�b����3���K4!����z�NJ���֭[���©�r��>6fB6DD�(����R�v~~��������III� �+|m�!^b���v�����3�3J���w""2M�/CCC��Bp�NX�R�gkkku/;���-B�*����t8��["]`�<�%laO�r�<��*��k ����pKtI ����~�������N��l/Н/�c�PS�/B��� ��E�wK+r�\ظ1�Q� ������������� �etvvv�Ƀ�&R�dU�E�xk|.==6l��|��������ּ��A��O����Z���Cyy����ߏ��I]�Bq&IDDƋ�;���b)פ���x<cpJQIJ)|>_-Sf k5�<s�R���h9�����L��B`�n���صkW���١P����輢��㩔R��"|M�m۶��r������Q+��LȆ�� ��#�/^�d�ٰcǎH����y��/�W4����U ���7l؀��c�ZfCCC�XQO�����BJT��������4̈́��WTT���*��3>��}����VT�x<_�c\|�x���Tl۶-f�˄��I�g+DD���,�:�����a��Ց�kdd䩇zHy�/�^��B�wIOO�֭[�Oj�(�Y$FD5��h���K�c�7���?���8D�	555���C �Z_��
T?�yH7!�,p'""S�������.����k����] > �F�~�/S1O�so����Q���b�4���������JIIIعsg��z	R��=�׍�+x��򅅅CB������*����ֲ���´����'��̥��i���M��k֬AIII���������52�h�v�k � G�Zrr�R{���:[����G������p7`ddĄḻ~�z(פ�_HJJ�U]]]��i�NJ)�^�?I)��Z�˅�;wZj¯jR^^?RY$FD��h��`zz�^U[[[�Sg|�AW^^��B�?T����b���F�e���Y����
b�;�*�����A22Fvv6�n����%�|�����v�?
����p^�~}�qXV �����u���n$�Κ�-�t���q�h�u��5������v���} �T륥�X�F�~/�����b��;�q�{{�25����ܶ��7"???��n�����?��gU�:�y��ZOHH�Ν;���dtj+fvvccc��j�$�'R�#���U	!�u�VdggG��=���]WWWhd^f���O�z�?�R��j}��BBB�ѩ����IL)��M�&dCDD�������Ν;����\�R~���=OSg��ۗ�r�� �)�zff��&�(��<C+��DDd��f�A��i���7!�`�ƍ��At    IDAT6�N ������ۗhpj�����y<��[�+ ���TUU������v���+���ڕ��t%��H����{{{M�&:ddd��[n��1K��^������Y�f8���G�P�} �K���BTWW���?/��c<""�	)Q٢l422���22�u�����������y�a߾}%yyyoPN�q:�عs'\.�������^e�J��E��a�u'T��U	!�}�vddDl�~K0<��x02/3x��r��w����c�$'[�����G,#"�:�zG����]�v-�0�ד��?t�ݱr��.����V�zZZv��a�)3�B����F~_\&dD��DDd���N���_ ���[�l���S�-���^]]]����?�A~~~�� �;��_��O�Eu��8?���&�!"�+�4kO���GGG�]��ENNv�����#����p���v��y��v�z<�G�?�lcRVV��^/����+',Uk4!""
�>Ǫ�Vf�ٰs�ND��*���K������z���Bmm�g�1 w�֓���gϞ�F��$MӔ��
zz�9<lBFDD�����t1)e\�]�n�c������Q�!���v�����ޒS^����R6أZOII���ފ��4�3[Y�@ ����x�ٳp��y#Q4��;���d�z�HMU�)��r���������R���xSJY��LVV��ٳ�]�%baaA�>���-'���l��r�3==���Q22Vaa�^s��4���vYJ��Q�x�����R��U닝׬޹��������I82""�p���d������Ğ={��q�LY(z���|����2�{��6!�Q ��3k֬Auu�%���Ϻkr�g�MȆ��­����9]��������y����"~���|����n40������n�?�B� (��RSS����e(�P6m0!""����^d]������)�qX��nǎ;PTT�#6!���|�7���G?�Q����/�|
�*�g��Ұg���(�
Ĵ���+���5!""��x�#Z|(����#.!�O<�O�4�w�������^�= �g


�s�N8�eKQ=DM��EES�	�P<a�;E��ǎî8ȉ�/����w�FBB��a�B��x�޷��߿��ܖ����W{��g���P�T[<�-,,48;s(��H�jdE���Q�tu��ʮ��$55��v\.W��8|OӴ�^���2[~�����z��
�= �U�B`ӦM���̝3FGG1==��W76�
���l<�����oB6�B���k׮]�c�C��q���O>�`čL,�x<��r����.��,>L\b�xLS�!�LO���Մl���z�
y���qAQ�nuBlٲ�Z��4��������1���������V �D���b7�%�*�,)�r�>:��N��#�/�N'v�څ��ܥ>�充�V���Xn�X__���z��f�5�D�ϕ��a�֭�٬_~;99���q]<R��r���0""�	�33(on�Ň��077gBF�����޽{�z�
 w�l�c����G?��y����K�x<ߵ�l�R�/D�\jj*���q$���A���.d��"�X����iZ\��KJJ�m�݆��۵E��oz<�G���b�ۥ1�l��ڤ�_E����D�޽%%�I�1K�ϮiX�	�Q$�ϜA�b4��Qu�������ۗ�R����j�z�_42���v�׸���@Ė�eeeؽ{�e�e���+��o�c<"��Vu�	���x�4>RY�~=�nݺ���$)e���?��x>mdnˡ��n���yM�s [֗��c׮]��:22�߯�o������C����vl߾UUUKM���o^��������������>!��� �#d�v;6m�d�	�עڟ�PՍ�&dC�ƚ���(&mjh@ǖ�W���[�Τ���8ީ��]���8�����?�x<���o|�c�eyc���R4M� �x�����z��[�����J"�Qz�,R��1��ܹs(--����H�mۆ��,���"�.& ~OӴ/z<�J)��7��UwuuuNM�~�� B��E999غu��
�fgg���*�[�<3cBFDD�-Bu�14�����SSSAvv�I��+//{���ɓ'�ݦ.)�R>��zC�������������h�ǳ�'����DJ��6m��#Ęw��9]�
aC�1�!"������	�ڳ����&''���nRf�*,,Dzz:N�8�|�u� ��x<��l��}�k_{I�������d�پ�i�o�x�t:�y�f�����񺻻u1g ���O�]7�]�:�f�dee��ɓ�W<V��!D���y���7��E<� �+�{��\jj*�mۆ��TC���������ᚘ0!#�7��NDDQ#��9��QOO��	�C�u��a�ΝHHHX�Y �@�����n�;�n+����gz<���4����Dq��nǖ-[�y��*n�4My��:>�Ҏ�""�%E�F0;;���2�N������[�r���X2�o!�z<��߿?�^3>��C���뚦���X���ʽ�Պ����R�=��񈈢��c��)Qw��w���d�ٳ���K~NJ�C�T^^�I�������K���v���x~��`�����t�~��/n���R>�+omE���	э�>� ����{�˅�n��z&��
�^�z�^������Qu��v�w���m6�I\|�1���L�~��/n��Ȉ.^u�r�E�����,�~���j�`� �x<��x<w�����������{<� ��k���[o���v����acT�Y aw""�*��;����b�����+n��/�����wމ3g������¢K҅�/<�+B�G�~�����w��WX]]�3~J�� > �Z�&??6l@R�5?j9����W�!8B��(*�?~����B掎�E��둞���{����]]]���@�?��l��x�B<"��7c:MMM�-//�.\,�"�k�����Buu�e4�~?Ο?���� O'""�LϠ��E7!oll,�����_�hnn����R�$�|����n���6��?��?=lT�W��~�~��l����v;֬Y�իW��޴��C���ł��Q�vt�g͚��CCCq�� l66mڄ��B477cf�)jۥ�O�|�A����f��׿�uSځ?���E6��wl6ۗ��[��y�Ӊ5k��M�۳g��Rb�#�'CDD7�wD�.!!�v�B?��ڰ�����?����MJ�����o}�[�qlؿ�&���e)��b�&������q�F����]t���Co�~s�χbE#G���w""�*U�O��;1�j�U���^���_����8�Nlڴ	���hnn^j%p����J)?���4��x�B��p8���W��oe�L<�* w!>�i�B�^ϯKIIAuuu\~ �`0���.]<iv�|�JD��fgQ}�(N��{U|vv���(.��YX�X,�***BKK|>�R �R��_<�RʗB�Л�����a.�|Е��z���~ _��z~]BB֯_�����J-*D*���&dCDD�k�{�s�FH��\Ϟ=��222p�m��������K}<G�-)��nw��I)�)))���̭T�uuu���} >>���)((����㦉@���E�Ρ@qKDD��u��Žˎ;L�(�dee�;�@WW:;;�4�P �;�P�;^����B����ï}�k+6*y����l6�} >�~ �%�6]VTT����������p�ϜA��	э��^QQrss��ގ����7�z!��+��G��sPJ�,�����O��ԬH���GAA�nM���l�AJ��z�)6�����-�-^Dj`���w����!�r`�;E[(���Ł�.����ׯ7)3seffb�޽���EWW��y���+Rʯx<�& o
!>B�-,,���?��%[����ե��u���c'��p�{��z� ��W�^������"  }}}�W�[>� Υ_7�ɶ|�!Zv�Rv�(**���#%%;w���� :::0==}�_���B�/��vx<�n)� ޷�l�6���k_�ڒ��*���	���U6�m���\���*�t^��.���(--Eee%����e1i�@>\�� ���MȈ���W�χ��tl�tU|||>�/n�_I���2��磽����׺��b��B�����{���C��[ NJ)ۜNg���y��<)e5�� �p��iE7��LOOǺu�����*���cp&DD�Q������Y��cbb&e=����Daa!���188xͽ˥��[�5���x<�w�o!Nj�v&77��K_�Ғ��*�:����l �%���[FF֭[������ǴH��w8h|2DDt�xG��t:�q�F�����������%6\l�x7 �����^��R��P�Yq�����\����egg�v8�B��!�= >
�҄��?�]���X�v-RRRn4˘��G__�.�x�Hd�Q�Ys�4��y&�����PQQ7��-^��������������_�	�k[J	����3 ��!)��i!�4�I �W�� �M�J�M~#KHH@yy9���`��o�_a��)��'��r�6QH���ƣGq"�C����ף�� ����p����09y�o�ʅ����4�gDJy�f��0
��qq/3 ���Y ���W.�p\+��v�����D����dg"����Atn�Vvqg���KLL��͛QUU���n���);S)$K)�B�\<��4-��x:�0`��bZJ����+� R���B�b 뤔�7���U�PYY���NNNbhhH/��Fa��Ś�
܁�{��;w��QtJNN�֭[�f�tvv^�#�K\ >)����B�|���s@ǥ��ԥs�i)�����\:c�R�!���9���w���������+l���Qe�_yk�i��(z�(���t�޽���������O(ɑR���Xl���xf�mR�\<g��Ŏ���L!Dڥs�r)�: ����!�@aa!***���zC�֊:;;�gd;�q}ggD˂�DDu����_�*��ى6��Yt��l(--EII	��ݍ�����W^�gE_'''������q_ؾ�ܹs���>�3�bSB��hm9��w�D �ع�����q=�d)B��� �����N*�B�����+��ILLDii)���,߱�J333��s�ٽ��(Vd�����g�l�*>11�.�
��ɨ��Fee%Ν;���>n�����_5~PU��Q�.Bdgg���".��utt(���9`p&DD��o��]{U���a||��7�̒RRR�y�f�Y�]]]���G0��M�� 6.�W�*Z������������n����BJ�8��Q,���233�c�LMM���CCC��P�J.)� ;��ܳ\�>f)v�������Drr�M�;����+�������ل�(�������Қ�&��L��V���Aqq1���L�,z!PTT���"LOO���������7;58��塨�(��c_�����{{��,�LȈ��nFҥ�'������,���QYYiRf�#77��������� Ο?����ӂ�fC^^
�����D[[[#toǄl���f�8p ��6"v���҂;�#�/[U�n�:�]���øp�.\� M��N.�(..��ב�u���N��{;Q������Y�}oii�m����ϯ%))	���X�~=|>p��.�ZN.����(**Bbb���jppccc�xyk+����-E�]���4l۶�@ ��������Ȉ�iA��������ô�����8 �L�/,p'"��$B!l�]���/\�R����v�2)�蔚�z�vdd.\���(fgg�!))	YYY���Cnn./�#hkkSvR���!8]݉�(zm��4�ډ@�%]WW������dRf�%))	������122���i�.d��������a���|>�.��ߏҳ�N�DD����P�Ԅ�-[������ܹs���0)��'�@^^���a����all�f:��t������FAA�=\"�DKK�rmǁ�gCDD�)gpeg�꺸ONN����())1)���X?//���0���{�w�ޥ�������w���ihkk�Ņ��q�{"�X�;���t:/7o����|�2>>n�=���@ff��s�Xo.kx孭&dD��DD����q��[1RPpU|dd���(���Ĝ��ˣ����0::���LNNbfffY� !���|��2++)))��ku��������Q}��	�G���c����p�=WŃ� ��ڰm�6s�a��U���`tt���Y�KY!���������,dee�`�H���{^������#���tUW#��*�����4����Dii)JKK!����$FGG1::���i���-���p %%�V���Gq8x����[9��������DD[v��&���thΜ9���|8�N�2�			(++CYY�����������0==�lS�\.�U{�xnIGG�r����	�b�v"�X�;��������JTVVB�4���attccc���Y��			HMM��O����D�k�R�5B��7�`�v2OG��(j�P���
���/�FR���!77��eא��t�%,pqC���1;;���i��~h�M�!���N�v�v�IIIp�\p�\HII���-�e��^�C�՝�����>@�-�0�j�U���A���"++ˤ�b���DAA�U����033��������=��f����v8��v$&&^�Ǹ\.N�����[9��t
zzLȈ��>���ql}�}4����⋏��n�jRf�iq�uFF�����aff���������<4M��?Y��]<_q8��\RRR.���a�6??���DG ��^{̈́���h���a㑣8}랫�@ gϞEuu�I��&!233���y9/�[�ܻ\yW\,`��l����J^���p��������'DDDˎwD��n���# ,,,\u���p��e����GY<oIHH����#oܹs�0==���>s�~�4,p'"����ׇ��O��i��͡��k�FU�҄�/N���@+���SSS�xqg'V�9cBFDD�욆�_~/��o�֚��q�w�Q�2JJJBRR����N�r�����ե�;��q�o��-�mￏ�[6c2�Ru`` ���Xv	K7�n�#==���f�bymmmʉ>[�?�ԉ	2""�����tnڈ��ԫ⽽�(..�߹������ ---�B���w�A�b"��-���$$$��`ʦ�`�M�TlYFDDQo�o A121�Hb�h377��g���6M��/�bBFDD��J::Q�ޮ����(�4E���e���w�C��������P�577Cr�0ŀ����ic��v�	�JI����7��ť�ܻP̸p�|>�.�5<��&dDDD+�wDd---����C��66nBFD������^���8���B!�<y�������.�����>D��	�r���k�+~��ە<��I__���t���Ql:|؄���h���9�R�����i�+.a��I0DSS�rm�k�}8Ŷ��N���G���@ww��	݀��477+����
l���DD�xGD����]��>�
��X�NDD1aӑ#���'''���iBFDק��G٥�55�m�gBFDD���ư��u�P(�ӧO�AE���Y���)����
슮�DD���������n���5E�����~]���egΘ��8)���� ��,�h��Ԅ��]��t
�ɗ�ȒxGD�jnn.bS��_{NE#G"#�����b�-�ޗ_�Pl�;::099iBVDK�����	o�+���8�$"�ص����66��ONN���Ä���&���ӧ�c'+��Q����DDV�>6��￯�U�i�    IDAT/�}��QE�.���_w����MȈ����=8��]\J�S�N!�.��"M�K��í��nBFDDd�Q,jjjB@Q�^v�,V���#��DD3
��`�#���'O��E,E��CvU���S�P�/DD��pϳ�)��uvvbLq�Id���n��e��4ƈ�,j��w��?������=�̲�����f�ڞ��@:��DD���ͷ�12��OMM��ٳ&dD���,Z[[�k���2R��Έ����p/�(���������I����MȈH��DDSv��&���u񙙙�������ى��q]�55��^yՄ�����}}�z�]|���Q����VH��^xI~��Iъ��B�����P<����Ű�̅�,�O�Ƃb�]qg'�MȈ����p�3�¦(������	Y�I)��Ԥ<�+omCUS�	Y���xGD1����̙3ʵ;�0��܉�(��5{�9�af�ׅDFS�R��g�C�ܜ	Y�Qv8��tq�ߏ��2"���i8q�r�{uc#J�����2}>�|�-���ӧ1��Ν;�|p�������4!+""2C�� ����..���ӧLȊ�j�)SS��Ev@%"�';@v�;�HSʈ�
�p��q僋5'O��w�EX�NDD1'gp��ť�8q�����L4??��'OB*.Z7>���n�"""C�4�=�,�Ψ�ϟGOO�	Y��ӧO+��icc��ƛ&dDDDF�|�������Q�L5>>���6����"FD��|����������Ǖ��DFBgg�~AJ���H�<"��b�4�Ꭸ���wDd���fLNN�⮩)�}�U2"���DD����>�Ο�Ń� �?�����J[|d��v���a�[o��"sx;�9�\kmm�m2Mgg'uq[(�{��&dEDDF[j����;��i���p��1e��S�QɟM"��d�p�s�á��E{{�	Y3338u�r��hJ�����ec���(�xGDf����yE���w?���L,p'"��d�p�3�"q~^�633���&��x��܌��1]���_>�<|'""����(VtF�R��ɓ�QD+�����ٳʵ�"O������55��_zY���ߏ��^�3�x�8"{A��.ml{_V��Q|�����וk]]]08#�w��El��5<��orJQ<���(���ŗj�G�������ڪ\�z��;gpFD��w""�Y�cc���g!]ѥ��@�Rz{{��ק\����}���ل����_"ubB�6??��d(�ߏ�'O*�V��a�{����	[V����`||���(�577cB�wv�x��FDD_664`�ɓʵ��&LMM�ų�'ObzzZO�����'�LȊ���������*�Vp��	�B!2�x4??�'N(�J:;���O��:�����bZY{;�8�\koo���38#�G���_�n9|U�N�E���Y<�ē�)hnn6!+�7���رc(.V3}>���� [ŭݯ����$������Q�iD6��ǞY���'EDDQ�_���~}���ﾪI D˭��CCC���p�3� M1허��O��,>��S�;���q��!���+�����_>���X�NDD1oǻE_\�x�nc�������ب|]]�ۋݯ�aBVDDMrq׋/*����p��Y�3�x��'Vu�s��で�F���5[(���|
i����y9r��b�����"6���!T����`��'�D�̌n����������ŋ�����y��~%�gDDD�,{pw���r����hoo78#�'RJ�<yRY7���'�@��oBfDׇ�DD����/��LE''M���بH�Q��͡��A�5ub�?�$l|�JDD �N����G�k8��J�Q-\*�I���^��&"�����_�:��~;;;���F�ъ�8"�����yǄ���(ڹ&'���O��؟LNNFlJC�Q��i�����6l;��Q,�:݄-�+�:;;���mlB7����Sg ��_���kDт�DDd	��'��@ �M�jaaG�U�\9�A<�ēH��5!3""�V{^��z�kmmm48#�����?W;Dyk��Q4˾pw��%�����?�,B&�Y���qGd��{{������Q�:u�{ZVccc����>�g���"���(����̙308#����6�?^����!�=u����n܉��22}>����ʎsss8z����6э�4�Q�@��~�9�H�����B!���S�Pt�^�=22bBfdE������S�U55a����ł��NE�;���P�����L�� �~?>Q���&"�k�|�6=�\DKK���UMMME|��2=�O����;H""Z�-�}O>���*�ĩS���X�nBWWW�� �Ϝ���64���w""����N������֥.Έ���i8v�&''�뷿�
*xhNDD$���3?�9\SS�5)%�;���q2#+9w�:;;�kK헉�� `���`CC�rm`` ���gDV377���,,,��� >��z��>]�������f�Zoo/���Έ�fffG�E0ԭ%���S��i<�#"�����ӏ���	ݚ�'N��}d}}}8s�r����>�KṆ��w""����&�}�����8>�N�tS�� �;����w��Q]@DD��51��>�(��@4M�ѣG1::jBfd]]]s��q�SO)']鎗_��x���MMM��N7��������+��_�x�4�"L�!""RR�g�Ei���wggg��k����ѣG��A|���2!3""�U��)|��ǐ<=�[�hhh�_�i}}}h���3kx��áx�G�X�NDD�����T�MNNF<�"��Z_&���#""
�>:�O��N�~D�4466r%ݰ������K���R��g�EI�B���>�:u�E�tCfff"�CJ��(={��Ĉ�(��B!���ȏ�H������ܻ������Ç177�[��y�����ź��1|����y�Z0Dcc#����n�RM)�����G�b_C�X�NDD����t��rm�C)�p�@ G��8�r��DDD������'`Wt�^,r�p�	�Q,joo�X��g{\95���(������F���r}`` ǏG�#��:LOO�ȑ#��n}��;y�ଈ��J� >��zdFh��ۋӧO�ȝ�����=��-%���K(om3>1""����|��'�wD�PǏ�]���.�D�Ƙ<;�O��gHQL �v,p'""K����Q�Ԥ\[�k�%���8|�0&&&��e����!x(NDD7���w?�l��0)%N�8���A2�X��҂�Nu�ݔ�i|�Ǒa/CDD���<>��_`հ�Plhh�E�tM8|�0��� `ǁ����gEDDV����ӏ�ic�f5����BC�4::�#G�D,n��װ��q�#""�)���=�|f�;�����9s&b���Y|��Ǒ1:jpVD˃�DDdi"�=�>�������Ø�KER���8r�Hğ���<�ē�)^U]���f�����.RJ�<y}FlS|�R�ԩS�0;ub���O��{��H���gy$b'���a444��(�D�~
`��obǁgEDDV暜���ӈ�����A�3�X044���Fh�s:!%�|�el�0=����fT���'��]�7�� �7)%�����ե\O���gyY�@1��DDdy"��^�6xX�>77�>� CCCgF�l|||�fff��U��po���DDD7ju[>����\XЭI)��Ԅ��&v��� �=���~�z��8>��H383""����Y|��ǐ�۫\]�;4ŧ��^444�/u?���!�#""�K�����S����q�/�;wǏW��B������ф̈��������N��3)%ZZZxGDW�4ǎCo��:��>��G"Ne$�,p'"��p��,RG(M�p���/)��������XP���F���,n'"�eUt�>��_ Aq�	\�������Q	333���1a�d�χ���G�݌��y|�񟡸�S�>;;�?�###gF�FJ�3gΠ��Yy�.B!ܵD3
""�����S�=��S񦦦p��!��ax��B8}�4Z[[�{��ᾧ�u'O��ŋ�s���Cb�x}}}��G  �ߏC�axxX��6>��=�(�#�!��Q\�q� v���rm������|���z����Q�����!"�P�Ӄ�<��"`�|>vG�s>�~�ağ���A| ej��̈�(8|��X�֦\hhh���8��A,R	
�cϿ��Ǐ�ţ��y|���Q��kMG#�[ܿ�?^�n�4���/Q��jpfDD���w��U�gÇO&���A�¤hpDQԪ8?�?����S֢ۧE���`3fd�L��@BƝ�~��ivb��\�������b'��>����ֶx����K�������3�i���g� q��0��]R�E�ȱ}���%��˽�:͌����Çso��f�=_�#�"B�����-v��~�@��vTƦ����	���hj���r�� ~�2�x�?G��������UUUL3�.]�p�؜��x��E'N�y2 ��9##������~>66'N����z�]���[�sݐ7wp0���Ü/w�����=^xｸ�q?w���u���(//����q?_��b��; �����?�!���yOOO|����ٙ�ɘ
.\���Ҝ߳FG�ɝ;���<O�t���#^}���9�����(//��u��cǎEMMMο��G���|���- ��f��œ;w�C_~�����ؿ丙�kK{{����_�/��^���y2 ��=:���?Ž{��<s���8x�`�q2�Jkkk8p �w�E==��[o�ʦ�<O �8{.^��뱢����_������3�i ��ĉ'���2�����J��&	���n9y*^y���1Ǜ����q��!ǮqMMMQVV�r|џ��/��N~W��� �����ŋo�k'؎z���(//�!Q�5����QRR����~>cl,������33�<O�tw��x���r|��퍒��hkk��d�K&�����8v�X�[f���ī��K�; `*e�q��}�������q�twwOx	W��KN�8�9��jh�W^#n��)t��K�����-��FCCÄ/lq��p�B���Dk��X���;�w\��	���uw�˓l`�q��t�����/0,io�W�x3nn� ��1+��'>�$��ޝs;jOOO���:e��hjj���s�����S�]R��� ��+����~'�������h?~<N�8/c]S.߈��ܜ�̚�����{1�o��� �ok**b�{�Ǽ��q?�ÇGEE��.טɖDDl8|$����1�& 0+��m;?������Y.p�lY㜑�x棏�޽�",��%p`ڛ;0�}�a�?r4����(--�]#:;;���8:'ؾ���"^z���<N ��f������cv���###q�ر�������<��mpp0<8�x{z�7ߊ���<O �j�ٳ��oƲ\ۤ"���5JKKゟ��	��������?\���Ɩ={l I�Μ�W�|+�=��̙3g���9�����f�ԩS.�96�|�����g1��� H̝���>�99�]^.��kÏY�xCoo����q[uM�����=� @
ff2�خ]���%�~���3�_�\�:::bÆ1w��)������H���DKKK�3�2����Wqg�Ao����UUqcWW�~��8���inn����شiS,^�8���f�������1����W��c��mb $e~_��λ����Qy��3f�˙���(++�իWGaaa̜i�զ��?*++���;�y}}���O㖓��8 �{���Ko���=�w�5�˷��Y�&V�^3��~C�.^�ћ㶡���'��3��>��� ��s[uM���F�~�g��ψΜ9��ݱiӦX�dI�'��������>#���>��Ә�c�;\K� ����ͧc�k�F����ioo����X�vm���U���=���bxx8�;;c�_v���H��g��߈۷G�[�=������|��ظqc\w�uy������b�FGc���q��<N ?ެ��x�/���>���r\Zpÿ���A���-6m�K�.��I�we��hll����	oZ���v~����8 �4s����O>�������1t���r&��D]]]���Z(p�d2����N�ʹ�4��X��]�bn��� ��_��W���gD[�_.p�ҥ8x�gDW������������gfe2q�7��]�e1òF�	�; �/7vu��o���m��?�q~(����hmm�;�#-Z4��cDeeetvvNxn������� R1kt4���X��{_|!����\{{{tuuźu��[n���Xcccq�ԩhhh�0��ܹ���c�sy� ~�[N���~�����Kq�p͸g�СC�^zzz���"���s������Uձ��-�~��h���q�\^(�r��ذaC��&`�������~w�=:�[" �U�ψc�K/��$ψ
-nL؏](���|<��Ǳ��5������8fe2�e�����ӱ�c`��q�]�p!������o���5kV�'%����hll�S�NE&��yn��`l��X]]��� �?w[MM�W{{������HTTTD[[[lܸ1,X��)�HgggTUUť����f㎃�⁯��Y��� �C����׿�}{��8�m[�͜9����j�*\2<<������2����ɏ�K݈�UlAoo�x��8���q��G�]~���]]]�~��X�bE��d"���QSS�|'Y���?�K�4�b$ H�m����7���_}%�n�m�3###Q]]�q��X�pa��d"?楼���G���_~�-kd��
�����6�}aG4�{&��FCCC���Daaa�z��N�l6---q���������x���b���y� ~^7����G~8�>�52���1���;JJJbժU�v�ژ;wn�'�Ο?uuu���=��}}���ϣ��6O���kF6�*.�U�����g��㞻�R^SSSŲe��<)?4::������8�Ҁ�fc��c����s���7  \!3�������U��qa��q����ǣ��1֭[K�,������H444Dss��]f����c˞=� pM�������q������h�fzzz���4V�Xk׮�y9���/^������e�y����_����<M���$���ů���h.*��矋�E��=7<<UUU��������M���������/Nxn��`lٽ;69��l �r3�����X[Y��?g֬�\6��3g�DKKK�Z�*��������[���O�I,��X{�x����� ���[[���.*�/=�D������G���n�)���bq���+��Ҁ����$X_��[?�<V66�g8 ȣMM�~��8���q��G#����.���cɒ%�nݺX���WF&�����hhh��I6�.���v}7���i: ȏccqwii�����瞋�k�=��f���5���<#�"q�ԩhii��D���<#z����'���; �Huu���1�>�X����Z{pp�[�
c���y�t���鉺�������ꪪx���<? p�Y���}�a4l�%�=7�0�ˡ{GGG�^�:


bV���<��ɓ���2"�;[w}�Μ��t �3�����q[m]�<�|�.�����o;)//��I6����������I^��96���ǽ�|�&�� W�Y��q��}����(��|��~{γ]]]QZZ˗/�����?~���.��W__CCC��=2�������̱�<M ����/��K    IDAT�x����~q����q�]~F����f͚���v`~������MMM16���E==���b��w ����-�w�m����;�����y���/�;��ͱq��X��~�����������I��,�t���*V46Ɓg���͛#r�(322������k֬�[o�5ϓ^����?��'���쑑���ocsi�� \��?�~�a���({��X� �ٮ��(++��˗ǆl�zzz���2���&=���)��Y��ݝ��  ������?��_��o��y�r�moo����X�re�_�>�̙��I����Ψ��������W=�/bAoo&�4���/�os�o�5���ψ2�L444DKKKFAAA�'���ꢩ�)2�,	������%qwq���w �	���ƫ��U��G�n͹!5����Ν�_===�����]����l���d 0����?�4�=�~*ή\�����`�>}Z�~�4N�r]6k��b˞=���|^f�~W�ԟ���m����L�e���?��^�dI�������O�/8>�|�uVTFLr \���X�h�������{��^�.^PP p�Z[['��o����۪k�4 �e��Pl���Xw�xx��h��������+���aқ}o�����m� �C� ?�̱����`�;~"N<�@�x��I,�2��t�P��mq\��T� Sbyss���[Ѹ~]�?�D�.]:�#�+�ݻcik�T� Sb��`<��ĝ���ǣ��;#�##���t)~U\�����@���G?�[l� ʟ�7�9���������u; DĲ��x��w���(ʟ|2z��<�#��O��-_�_�93գ@�� ��34����#[����˹��<�fc�wq�7�Ă�@d�q{uM��E��w��m��҂S=մ���#ؽ;n9yj�G�$����>�4�*+��'��梢�iZ�=2���%�q���T� �Y��O����\��w��ի�z�i���\Rw8sFF�z HNA]]�Z_��7��m�G��7N�H��M���{����ک�����ɼ��x�/c�ٳS=ʴ6wp0�عS� ��̱��p�h�Q^>գL{��+q; ��g��S�h�ǘ�V65�}{���$���Ŷ�;�z�i���.�).��fd�Qt�x�]��G���|���~$�;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�         ��c׎    �[OcGq,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�!K�    IDAT�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�     �v,    0��z;�#     `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap�صc   �A����Q          �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           _�3    IDAT�;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;       �k�    ������8   X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X� �];    �o=��        ���          ���          ���          ���          ���          ���          %%K�    IDAT���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���        �v,    0��z;�#  w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           R�;;    IDATw           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w   �صc   �A����Q      � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          �k�    ������8��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ���    IDAT��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     �];    �o=��     ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�@�ڱ    � �i�(�          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap         G���    IDAT `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap      �صc   �A����Q   �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;          4A�_    IDAT �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;  Į    �Ǝ�        X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�        �];    �o=�� ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���         ��Y    IDAT ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���   @�ڱ    � �i�(�       w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w          �صc   �A����Q� �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �        �P:.    IDAT  � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �     Į    �Ǝ�    ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��         j��    IDAT ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          �� ��v)n#ð�0	8��V��=��J��*130�� �UU��u]?�K%����-	         �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w��q[��~�3Y���ǝc[ך�nwǙmq�����b܁���m��Lch|6�в�����\e�c�f�3�inw�s�i�����m�YͦW�)4��MS�18W��aC���L��/Իִ����T��܅�U�'��������I��⼺�/�W!6Ϸ��N�N��{8�O5�c�Q�1��p&0����������]��� Z���\e.Cc�ɽ�
myU���]�1t]_��А��ߺqe��ʺ�C����\e6�k s���ʹ��C{�o�O9������|�L2���'pgqN�G��Ө&An�к*�� �F=�����n�G�1t]Ol,аj>n=4!*K��|��z��x�ͩ�VW�Q���x ^�j�oL���u�RZv��X���83��b<1w�E��/���/K��|�yK׹G������#a10�)KdA0��+n����:�j9�n�#�6��G��R_j��F�rӕ�T+�W��%,��b�bL����}!W�XM�g|��U;�BI��W<8C˪h���F�����	�Y��u�YLahtl1@��1f�'�ld��U�c7D��ӓ,Q����83o�`)��L�)Ө����9�S]W��z!I��{8��Uc��v���8��|��\�D�s���X�4Cp�w��5j�]w�d�.7�noo�p6m���{y��M}Zqz}�s�3�j�9�v��3�q�+l,L�GN��#��l�7n�2����^w��sS��\�V�v���ٴ�W�n�]h�ٍ��9�}�����mMDcN�����j���ٴ��O��:и�b�1w���c�.�Sk"ZtZ������Z�iZh�POa�2��=>v?�P��8}ߝ��s���U�����=������α��;q������P�#]g�r
�|��E}��o����b^bM4�r����������E�<O5����A՚�zh|�ժ|�К^���B����k���
p�y�wn����m��������W�w_�\�.-;���;)s�h|�5=����C�	�Y$��yT����_}���U޾�-F6���w6x�^�ֽ*6��W�WFb6.i��v۽)�5ƌO��R�_^vEd`\_���������b蚾�믙��u�^{�L<��R��<��n���Ѡj��E�)�]g���}w^��Գ���Gti|�B��"U���ĕ���1�i��c6h��Ƃqd\C�KP�έ��W�1�t��t��~�9n\�f��V���q�Ѣj���l��y�j�rzs���:Ӡ���*���M���"TZ�V��;�j����;*�H/]u�sh_����.'�uw�~����>����	�Y�j3������Owuu�s��l9�f(��O�t��<�l���~��������qd\777�cq�ÍW���Ab��j�*o���&�QU4��X�t߾�ksZ4��6_ח�>�.w�A�q�\e\www�����q_�a	�1��{s��Us�!ZeM4�j>���늗�AK��C�~��yxx(���?#pg�>��q�X��墘�Y���h�?�^{hч?��9vi�:��z���Sw��(4�������Ud�4�����c��?�������]�U��l�fh}��X�B>|��@n���Z��Zu���h���M�S�[Wu=��9�����y���ud�4�>�A�w�|�����y��|ѝ_@1w�н�_>chӏ��ݛ�7_���鬉X�����Cw}}���iӗ/_ʽ� �	�Y�����u�G�b`<C��?��6��~���������/E�dh#���:���D�q�[�U�W>��{w����l�?{���u���� 9D$"�����m9ɒ眩;s^ϭ�/flɖ���
�$[�#�sj��� �"{5����T�T�wX�W����y�k���r���R%��S��~"��Xu{�2��m��3��@>0�X��@ `�m�ly�cf����Ӄc�]6���<��h��U�J�m~>�9�����3�`�<�a8ka^98�pXa�:Ŵ�M�����?:8��ee @w`�pG�2mv�����~��s��t�̦=�S�����0&�D�|Ҹ��rC%e:F�9�y��,V��j�s�D����r�,S����H&��d���٣pDL��`PQCuT�i~��[��h��W���P4����a�Bg:W�z�t�< �sq{<n���Ӟ?*��`�P��3m�� ���:a���v`�    IDAT�����G���k �����n>
ɰ7�e��t�=� ����U�!�`�H��3�K	�6a�qe�,�ͥW�Y[[��h����
���w�˥T*u��3~�߸�4%A��8�T��b�s�.cmm��Җ����Vb^9(����˲����ԡ��t�����|>cR���G���eY�NL�;��u~AE$ ����I�u
{��a�=6���}#Sa����-�o( �Y.�w��`u��[8/��o.���޶�L4�SS�i���ֱ֨O�eiee%�y�ܼ��l!Ϝ��J{����0��bZ�F�T�AA9iX�$	.H�i�)J��N�/�\�a^Y__W0��h�i^����ࢻ�W�߯���"���_86v��������H$B���d(<R�L�}��(�kk���}X��_04v��a��V��pVk�'���b1cR�t����LwD�d�������Yk�	���U�������g��E":99��� ��?0��,�H�!�'��kl��?<��� �����1q����$�Ic o��PP:fgUe� ��?���NNMQ�y�pP6C���F�ƶ�����Jn@>9c8[Y__��>-//�W��,�q����5>�2C�q�*�cY�G��	��o _�,K���k�өx<���LAb}��Yp���=����������1��p�,-�ΐ�kJ^�ޘ�Gm���;9 �#��߰8�T�����c�TL�
L��j��Ӟsa�?�ߟ=W��XF��hT]i�����p�i����fY�31e�Ȅ�q�݊�8�0��W۬���{�.]���@��6v��uL�x-�˪��5�\q"��##i�WWW��3���k
����9S"<vǲ,�P��*	C�6`^�Ӽ��t��Bu(0}�{���u�)���<��0wD��!���ؘJ�n���YM~X\\Tʰ�:C�"�ڬ����-?�nO$�l�GFe'y�ٍ߰�b^�i�W��}���(<�.^�=�YCpoi4������y%
�ᱳLsr�ꪱM9�o*�~��ͥ=_\\4&�bg.��X푤
�9K2��(�>����P���(H���jXs�=����`�Z]]5w�e�Q���o���{�'��z������y����PZ�H��Ǵ?*ɐl`g����3TE]]]���H&��`��W���G?  �2^%iff�G�fggI�A�955�2C����4�"O��t.M8@!h\]U��|�Jý[__���N{��`D��>Q ���Tb��}zz:�9�VVV�����BbJ���bTqBSSSiϊ�I�>x��� G�m~^U�s����Y��������wxXE�s\����Ճ��V�
�DL�i�x\�����a�ofO��LgT�T�.�(H5^�Zs��⢱K���^���Tj��`g������V�3˲�x}KKK�*(_�u��1�z�K���7��alK�����2N�:H@+J&���{iϹy2�5^Q2��n���h��p���Ҟ��q-,��`��I�������4U�����>�Ϙ ��2�O�c1��?#��wxX�3�Q����h}}=�y���i?�a�,=}�v��H$B��0�Y�.p΂v��}cq��.c��{��ꋂ�;2�
C�F�D{���!�˕���ؘ*�,�Ⱦ���D"a,p��eZ�]��;"�I���׶�������L�`�J�������s7#rǕk�Ӟ�H�w����J�Wo\���之�}g�����޸�nc0Ǚ�Ac�6�P�T�ߟ�<ӿ�0������j4<�ٕon+v�ڛL��}�@T��x\��6�y$1&�#���ɴg�TJWo���h��9����8g���gU��9P(*�A�3,�tn��2+�r�,�Ȟ�x\EJ�흩��,KW��@��Q�כ�|aa�*�{�p8Ҟw������IW�_K{fY�FGG�0��izzZ�H$����3V) 
I�ܜZP������H���5^�z�i���W���􄱍����eY3����R�r�`��dR��I���b��A����k��M ��x��kX�{<�!?�%�IMLL�=/N$t���Km �e
F����u������#��x�0" {J�Q���^�0
inn.#:~,���Ȉ酮\�q�r��7U�L�=Sʐ�t����R��=����nc�Q�䤚蘌fK�t�F�>��a6::jL���5wD�~�H:95��+i����Ȥ߅p8l��^���[�>�Bd:�ߺ�*��<x`<��z���2$������x)2>>��Xw477'��Bu���9 IOݹ��P(���쬱z0���$�a.99m�k���us����1%k<jzzZ!ü|��]Zf� �F�:�}z;�X,�e�.$�Ic¯,KWoP����7��n8O���4���������ҞwMN���F@U~���=�B�b>xT"����x�s[*��+A�ʔ�Ǟhw2&��|��Lݮ�Abَ���U���I��� w�����磣�\�� S��k�Uj�"
Q�Ԕ���Ӟollh�P�����j�Ի\:30���Q����o�I{�Ǎ�=�/�H�x�[�L�ٯ����S����eY���x<n�t�,=�a�	�z�K�CCi�#���4
�Ơ{4��7�@���wƄ<.[w655e��RÚ3#��<��o�M{�1!e��Rz�_faD@nz��uc��Lɬ����	Ew���ݧX	
��o�U9{�'233c,��5>����,��-Eɤ����e���m��vE��⋣�gp~przZ=����p���m,//g<��-���,K�~����������b1����~�@>{��/UH?�[ZZ��������ac���7�~���;j2T��z�Z�?���c'����Q3��Q�^��c����Yc�O�+��TH�ٯ���Б(e�^�<�bв,��@Z__7&͔E�z��V�+�o�f}=��ᠻ�6<x��!h���;jZ]���T���+��;�$�IŶ��z����C!=��daD@�(�����m/hzz:�yI"�W���,��Mg�j�7���i�*����f,*�>O�K`�p~�O>5V����0� 
����w�~򩊨|<����C;�D"���3��������au��B*�F��知=�,Kƪ6�nvv֘�W���2m'�G�R)���G��$###�T�fqqQ++�A���0�I����eY�w�10��MNN����=op�t�B���}.�C���7'��x<���A��s��R�@F䎒DB�~������EI�0$FWz�V@�+�|�:�٤��6[�x<���/���p8�r˹�����~?]h���ݻg,�t��k�dG�`Y�^��cc����q���%���0�*�F�"E�A�;�#����~}��nhhHa6��R)ݿ߸�R��* �ٯ�6V���|:<fffƘ\T���?���П���X,����,�#>���2[�^��S�	�ҜX^��{�Ӟo��/T�@ c ݋��KW�Oߺ���i�#���0����x433��²��'t�$I��W>����aaa�tY�2�6;z���,��=����e8;�.ȲPm�z��ύ�{�BW�L��O�f|755%�%144d,ztbyEg履Wɲ��_?2����J7�G���(L�\�����faD@nkXs����Ҟo[�`ɿ�B!�=��/UIQ�@�<��w�3^�3i�������H{^�eO���Ѩ~�+����q��ǣ��	㻗��w6(x����������TF�{b���ݻg���RW�9���矫�P�#jhh(#�=�x<c����I�%hx�fY��_?RI"����tj�yI�����߹�v:X5������w���
pf )s��DB?��/�q�<��ǟ�ܐBQ������vML�o��@ꜙ�Sw�=�+磦���k��x\?����j@�jt:u�z�=�)��-..j�Pt�(��O��WΪ H�}���M8���I���ɤ�ݻ��ai���� p���ߚ��/ۃ r�ͲtrfV��/)a�?�.�(���M6�-K#̾��I�.Vm��~�ޟ�h8| �/u^��%%Z�:����t���AYYn����}��1��`P�}�UF䖲pX5>�f�~*���Uyy�jkk�0�ܐL&u��-�!n�ǣ7�{O�T�2*I$Բ���+Wd=��	J&�jnn���/�J��ݻ��|i��~��λ*��	���`Pe��ΜI{��xTUU����,�,7��qݺu��9����/��>�ہǴ-,h��)���y�J��t:��֦���,�.�VVV422b|��#�xLi,��KS.H��|>�JJJT��|SH��@��GU쁀]蘙���s
WU=�<�L��v���]EE�[�pyy9c���?�D'���xD@�k_X���[���G��R)�\����\.�=������Iq2���M\���c�`0�h4����,�.�,��ݻw�n(U�����X���!�0(�FU�t3�����Z[[�4��Z\\�X��ٯ�����M�G���k��i�=t�,Kkkk:q���ʲ4��	�B�u떱�U�ǣ7��A���N�jj�joK{�r�
6Pl�P�����+N$��;���
�QU~��I-����[__Wqq��0��ڪ��2T/)J����S�� ��ʊ|�M�.?���TWW����,�,��ɤn߾m��bz��wUA5j �ͲtrzFS/)^Z�ȻD"!�˥��vgi����x2v��ы���Q����Q��T�'O��s�ݪ��(�b;���Gջ�Yp��Rj���ĕ�J=�>��b�x<��r�t��}���a=��퀀cbsO4�ɋ�xlO��zO���t��c1���Y����t� vP�,���w[瘍��G=��044���մ�6��/����dx���dP��(^Q���δw~�_�TJMMMYY�8�3Y;�����~�F �%�e���&._R�n�T�a�{�c�,�����ƪ�%�����Um� 
Y�̌�ΞS��?Rav�غt5����W?��J���.-���.����v\�˲�������?���?�~	��ΙM�?�XEyڻ��5555��<�]�J�R�w�<������� l��bjp�i��Ŵ"%�x\^�Wmmm(�����+^�׫߼�
 �h���R_��55i�N�jjjTe8��W;큞��?�?<|ģ���PH�~��ΝK{�F�������޽k\�Թ\����	l�����6n��b��|jmm-�=Q Э[��H$��Uz�w��=��Ȁ���ʊ���Z?q"����n/�NW###Z\\4��z����{��G�?܁mt����n�X__W<WsssA4,..jhh�X�����o�yWvZP{R��uiI�.��vJ&�r8jjj*�J��`P�n�R(J{W�J�~_mY�ۊR)�������iU-˒��(���d2�{��en����z�ڵ#p�����b��N�S%%%q��J�488���e���z�j�����I������J<��kY�VVV
��{"�Н;w��P��ٯ���[��xT��S���,�bzE�H$"�˥��ւ�Z�r�t��%A`��~�_�S!�m�,K�&&5��S���VWWUQQ�C |��*"�8XM��J��Z=u*�]0,�`T�ө�w��.��~��߫2��Ȁ���=�Rooڻp8,��S0{��������Ѩ���;�3t��٩�)���V�P�h��S!Tr�,KCCC��{<�k�|������6l����19����K{��������ښ�A�3335�����o��;Ur9<�j�O��k�9����摭 ���ڼ����Э[��F�_Z�^��c�Q	Ȩ,���iM_��dI�#�,����JKKUgX��x<�m�X��^��#�'P�L����ϝS����v�}��N	4]��z���f�Ry(�����D��.W���+++�:p,���ￗ��3���]����G<*��jY^�U\,GWWڻX,��K���Ě|������������z��?�"�%{,��IM�Z	Cw͵�5���!�;�D�=p�:gg�����-�](*����e�.[A�?��Y��b��h4*�á�����m%͘*�%���{����S)u��i�L������U$щ'���h5ùJ�ܜ~���V�a]`�pvP�J�{|\g�(R�`��zu�ĉ�;hH�Rz���fff���"�����<d��Q������3i��R��G��:�������_��w���"R��f!�̓=˲��ؘw�[ 666��;gf����3�
�>��quMNe���|
�:q�D�U�ú}���*��,.��?��v��U��jZ]����i���f�XQQQ^���~ݺuK���G��Ƈ0�Q�ܜB55r�����q9��թ�w�Y�������I�R)�����>7w�#���HDs�p^�Ǌ	H����u���@�!;59���x4���TSS�J�0ǙeY���μvI&������Qd�9;+}�<��i�������Un�Rs����khhȘ4c�,��������,��%���'&4��ӊ����������jnnλ��H$��w�����79z�we7t� p0pv�$��!Ƚ_QC�H$��������%I(��۷�t:���"���?���8�����Pi4���޴ wi385
���9/�R��FGG5>>.+C����7��W_�Ȁ�Ʒ�FǪ�z����z��x��Ԥ���q����;w�;@Hj��כ��I%* �V���̬fϝ5�������Ae�����p�Ν;
����'�W�ֻPi�9���<չ=�;w���v���������ݻgl�-m����Vc�955%}�<�-i�ɤVVVd��T__���XL�����Ғ�}q2������'&�xd@~�Ժ��٧���}>��n��������ڶ{�f�@���Y�����<�)}}��x<���e������6#<x�Y������59u�#�G�Ĥ֛��~�Dڻd2���e��0�G�DB������5���Rz�Otf`�h��hT]SӚ;w������W�4N�S�o�V(2�o\[��Ｋ��' � w`�Jc1�=x���n�m��.I$����X_�l�E"��J�_���ߩy��v� �,-�nݫ��g�[�c����:pl+�&S�[�e���>��k׏xd��W��mn^sO�S�p����WSS�JC��q�L&5::�����I2�cc��{"c8@��z��5�_1Cbo<���ұ�|�q"���$����o�@`�_N�N,/k��9�A�PH+++Ǿ�r"���А���3�]����ߧ*�6����q��˴��i������;�U��n�n߾-��o|o�F��?�Q]��G<2 ���|:93�����HD��˪��RUUUFx0R�����4::�q�9=Mp;p��R)�?������J�����p8����c]�����֭[�.�Ѩ���u��v`_l����1E�*���0~��v�E�卍}���Z__7�/N&��>P�����_塐zGG��׫��y뎨���X'�X����	���d���/�����v���AI<���ay�۵�hn���x�������c��
�v�p�s�����w���~��4���eaq3�����)��bjll<V��ei~~^� �R��G��۷�xt@����Щ�I͝;k̠�J���jhh8v�kkk�w��nw�Ϝ�{Oo�χ���,Q�ȈVN�V��:�eYr:��z����;v���n��޽+�˕�3}C�����$�8����U�̬�ΝS�P�4�HhyyY�hT����n��"Ӆ�$]��[���'�e8��7'��U�h)C��P(���%����X*�������"���~�]�-.���T�������(V�~�J��p8���p��m�2u���a���쁀�P��ZR�I�  2IDATQ.g�=��/�á���c�L��522���Q%3��V����Q+k�@�$����,i�t��3�`�a��Cq�\�H$411�����J�Q���H�Ai4���a��:�`]��3.�KN�S����.n�����ݻ�5JR���~���TJ�5�H��Qq*����������X,v�._S��fff400�@ ��s�s�z��wU��g �_���:gg���gN�6[�.//���\Ն�\�r�t�����d�r-���������#�*B!���j�t������0����6�:�ᰆ��455����fYz��� "{,�������h�L8��⢒ɤ���r>)/�hppP�Y��޸�W?�TE�3 �L�߯��	-��(������Ʊ�|����L�@��TJ/}������#��Z��U���b_��CD*������Rmmm�wʳ,K�w^o��5�9����Q�6�� ��,V�ȈV��̰	ZXX86�3�HD����vt�o��ǟ��Mҩ�)'Z��6&�%	9mll���^vCrp.�,KKKK�{��ɾkN����~�B �L����6�Z��e8�M&�Z[[���96�Jǎ�I�����;�ui�G��DB���Ԥ����D�Q---)�����X�m�b���C����}�����Y��-��I���&/_����R|�ž�nשS�t���;lH�RZZZ���L�j��f���k�����d�82��J}���[����~���^===jii9�������Ԕ<;t}h�_���_��Sx2ɒ����5�ܳ�~���Z���jkk˹�H$���---e���@P?��u�����Bg����/����Pj�����R�>}Z]]]9���5�,..fL6�~���NMM���/-յ���ԥ��~���F}}}jiiɹ�K8�������2vǓ�j�O�x��P�8T����?�S�'Nd���fSKK�z{{U[[{��ۙeYZYY���̶�I��NV�|�)��C�**�����_|������R������ȹ�J4����=g)�����P]G8: +�]�����kޖ��"uvv���GG8��Y����UMOO˿�}Ϲ{��ʧS	�O�C�jk���?��А�36�M���������jN�S����&�H���1���U��� ���կ�����n�����:u�T���E"���iqq1c�<i���O?����Ǝpt $܁}�57�����lsI"I������RWWW�[�$�I-..jffF���Yf�i��uk��1i3ȣ��W���Y�8�,K.�kW6���7�̗_Q8D�.��o�Vl���/`��I
��o&I���z�>T]f��X=yR_�������ݮ��n�:u*�����fggw5Ǵ����|@"p�ƞ������%%�~���J���joo�z�X ��̌VVVv�W��������m� 88q�]7�~K�/�����f����a�����L&����caI�G�z���74|D�0������K�K�����ӣ��ά'���a�����+I�����jc�F���UU����]�}��~�f����C===���:�љ�R)9MOO+n�Y{4��?�D}�CG4: ��2]���j���m?g����ڪ����'�n%����hc�5Iq2�?�L��uD��c��v}���!�g)%%%���Io/����%���T�C���A�;p %%����4��;��l6555���C---Gv�iY��n�VVV����m�ٖ��Q���'�l��9;�u������m�ϖ�����M��!�� -//kyyy��I�s���ǟ���H�t�ok��g����v�������H;��VWW���,�׻������k]��[�v$p����ؕ+�V2�6�D'N�P{{�ZZZ�,�&�keeE+++;&�I�=��k�t��7$�Y�=Ѭ����N��Y�ݮ��v�������F�ik^Y^^������eѨ���:���8r3���替޶"���Juvv���M���G0���[�׫��e�������svV�}��jw���kku��4�̎�-..~x^���pd�y�D�s����J	]�~CW�_gd�e�i���u�g?۱h�$���=\�eeT�ϧ��%9�wQ��}nN������#��M\���~�K�w�ǩ��}x�r����pws�ܼ��������#�Lbee���74�쳲r4nn���ŉ��ܸ��?ڦ���E�;p��'�u㭷��ݵ�����E���jjj:�6r�XL�G�GN�S�HdW_W����O>���������4��s������ABUU������ب��F��Pq/�������x�r�vl7��$����u��7l�,�>^���W
������+=�H�U��n��n�\.׎Y�[zFG��S����v򤮿��ܭ�����nd�r�d�e)<�c�n��[�G�������]�8D6��/]����|�6�@[k����� ����@��W,K��Cz�/�8dY��Lw�S?����J����=\�t`ꓞ�Vz�w���@�͟9��yS�]&ٕ�����EMMMjhh8�@�`0�ȼ����k��^��S�x�J�Pu�����4u�®>�UT���I�����Eb�^$	y�^y<���)
���*A���g�&�ȲhE����=���]�m�Q�bZjjjtO�L&�+N�S�]��lx��]�H�r���]��~KΎ�]}���D���癃.2�u��uG��{�S��z�ӿ�f�� ��A��4y颾����e�ؖ��
544��������+Z��H$�`0��������M��F��t�]�yS��9+\]���sM^����Xi� ���N��ժ��z�����m"~<ǄB!�A��~����:HL�l��ӣ�z��/h�dY��Lw~�<���{X��l���U]]�#k��$�%�ɇ�H(������U�kp���g��)�\e��������: uKEE������D;����G�C�`P^�wW��~���ҋ��S��{�: �+Z^��?C�W�*�����=��ڥ����h'�D��%(���*��i���^����>����p�<--���_k���=}]qq������l�-;�+�e=<S���|�=�ߖ$z��-=��5��q/��$�v��5����{X��l���yxf[YY��e���T*���x<{>g��x���_�{llO_�h-�>�o~�<'N���JKK�o�]***vU���獍�|�=�'�z��=�嗬]������߼����=}��nWCC�����_���v5�D��G�E>�o���E�����?���`pOcp4,�Mc�<�;?��B�U{�����;����]�m�1�@@���{>˭�x��_�{���+pI��X�/������а��e��U\\��OQQ���R�����Ğ��+�u��u��T��pl��u���4~�Ҟ�<L���T\\������(�H(�L>���TJ��t��u58]��^ V��Z�/���g�U��􉿏�fSII�#k�T*�d2�p>I$�k�ág�]S�ظlT����ݮ�g����/�kD&[���#�=�~5;���`]���Ʈ^�S���攭??^�l�[��viY\��k��55E�B ���<�{�����>i�UKJJ9_ٚK�{v+I�hT�����o�����~�E=x�y�vف���k��9��k�d2��}P�ӥ�ׯ���UO���f��ٳ���kru���[m�-[�-**zd/���KI<������7U���iK�����kZ�������|b��UTT�H<K2��u�d��dRgu��u:� �D��DcW�j��������ۺ�.))�eY�7��F�SW�]W��# ���TQ��/����/��ښ��<�����[�u���	l��`M�_yE�/)��J�G������.߸�ZZ79-RY��_��3�(\��L�CeYj�_Х�7	��dq�Ư\���/h��9��y�fYj��ӥo��)��X	UWi��5v劢��$sTl����]�qS�����=p������h��9%�YD� U��z��]]������l�.E�����4��s
UWg{8�hY\��o�!�8��z5��Z���w��A��t��=]��[U�B��=p�:��W_�B_��=t?leѨ����7ߨjc#���REE��|YC/� OKK���/����]��;u��sG�(܁#�ii���K��x1k��e��zFF�74���0�<�,.���3��tI}}����$�R)���R�а���T�Ϫ� �V��H�}}��tQ�g��2�~Ի\�R�а�ש��WG�&.^���YK�it:�70���a.E�c.Y\��3��tI��Y�IR�����?<�J�?+c p0���>^��/i��3+c�ѨN���o`Pss��ǘUT���Ӛ�xIsO�S�n��8j�^��hX�OV� �p��5q�&/_���1+c(���=>���!���VUO�c-T]���5q�R�Q��I���T����&'U�}3�7<����|IS.d-n���R����s�Y`i��i-��i��[��Y�xYR�����Y���V������C�Y rC��R�g�j��[+=�usP
�mnN3�:=6��`��~��++�ܹsZ���r���#E���WV�13���1�X^9�� 7�����ۣ��^-uw�{�{��dR-�Kj��S�����C�9 �+RQ����i��i�tw+|�k���%u�����WW�gȞ��͝9����rtu)VVvh?�ƻ���Yu�̪k|\%�^@n���j��-��
���ϲ�Rjr��snV]�j]X8�� w�uth��-ww��٩�!V`��>;���i����)�S��͝;����Z��<ԢH塐����1=�ޑ:Xyn+nn��G���r���я�rOML����� �� w D**�8ݭ�S��kl���I���'j�T���V�ǣ��%��Ϊ��3�����H�9!_S�֛������)�T�v���V�ө��Y5:��k
���I˧O���&_S�|��
WV����R����#��j���(p��J�tu��١��&�76��ظ����DBu���P�˥օE�.,$�M��͵���M��͵K��b�ߪ(�R����].58]j��S�����+@A����lk���[��M�V�O0�T�|��xT�v�yš��9*���Р���r�w�״9������ʖJ�ڷ�z�[�.����67�2�Y��/-���VOu����e�	�Y$�,V�ǣ�������C5�\�()��ɓrtwi���}���Q�'�W��ν�'jZYQ�ܜ���^�hy���Z�ؼ#�55n�]�8�'����̥��R��g��1G�;������56*P_��ݮXy�b�eJ��e�$UY$*{<��hL����n-�Z��L�����+VV�xi������U������4�=U�׫r���H��B��&���/-U�^�XY��e�*J$d��d��T��$SͺO�^���&`REE�74(PS��k�xi����*JY��6�D%�����P���E��"���k��J��뗲R���U�H�$�yβ9�DU�]W����R�l@�
WVj���uJ�b�e���J���4��*��d��T
����R@FѲ�͵JM��b/ݜWJ�T�Jm���hT��S��C�^ ��**���^�J�K�(Wܾy/�,)�=yd�R���VE(���QVQ�uu�54(^��~臻�Di�J#����xL���j=U�:�c UT�@}���J���r�e�*�6�J���1Uol�z�;" ��                �	{�A                �! �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��              ��v�X    `���4vG ,�           ,�           ,�           ,��z�{>
=    IEND�B`�PK
     t$v[T��T$  T$  /   images/8ade0660-1c92-4b58-a3e7-adda420d3982.png�PNG

   IHDR   d  6   ��7   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #�IDATx��	|U՝���-�CBB$� [E(T�E֪�uԪm�Ng\:U�^�m�ڙV������� (*����,��@BHH ��{�����}/yyy{xd���9�r߹�����}{����&N�:<�����@Z�W������@�p&�i���4-��e�xd�=���4-��v���3	ߗ*�P ڔ�Я�
槟���#=�ȑ0w��Ćb@N�!C`n�����π6b8���- �W ��/g���sxg��eX�����d�&]6�;����}�2�~�+�K�v�z�r�n���~>�7��φ}����g07m���a�t���8�O���ۣ�B�:_�N�N�l6�Ax�8����>���؂�5G$�������6��5+u%���u�jBn�1�OF<�������:�s�(G�����������c���|�& �:�@DB��6Rc�l,�9��
D��y}���,�iM������gb�r���h���r�w��5�1��-!aY6��5������r�YGZ0��0h�ՊSʊ(3ه��ro�[M� 9*+PDn<��h���iN,��*�?���>��z?����]��n�ױ����no� k*
�t�Dx�-v��AzN��a�~ݴS/`0���$"�����I����#)g�^�p�15�˼{��o�𿗡�r��^�
�}���K�����F����d�j��r���^"���d��)=p���;qJ'C�2���<8ݞ�)�����8�^cߐ�[�J����e*��e\%<NG���}Q����]5��R��q����G�?���8��r�������݇�w��tת�c+ҧ,h�$�J�r�E�)�����3�=LTE��ܥ��_��>��jP�ź`��۰R�r#qi,��O�Tپg�2|�C�&��z,7%�V 䣺�h~����d��YM�pST]Q��zI[f�D��W�\��5� ���8�ꊢ�M_6�g��	�O���օ~�<dKk�7�j����=4���f��$4PVP���]F��}�D6�<�Ο�(w�J��>���8�f3����;�wj�"�+b�E�2���>8�v��\Q�q�=��;M�u�M��3]���zA��P��P)�*ˠ0�ĳG��hc��ѭX�B�3���M�"
�Ѐ��p�	�O��Cqj/�q}�ZВ��$ퟨ	��r�42���U�QT� _Eng$9�|�/-%?�:�����#�1��*���a�܄�<�Fw56�1�g��>�,}�O9�1\0t�^�BO����#�>���*z9�L"��p��yVq3�`?AP����D�{8���"g������	�9��*�␙����H�f��"��&,݌��G^�NsrN�P�Ɔ�����%�2q�&����J�1�vN�.�M��e�Q��F<7� �B�ǒ�:���e�vD.񒻗��p~��k"����2����E�����ĝ=g1�-Esvz&�'ʷDz�[*4�r��b�!�*�mT�؊���w�(z`�=��j����W�PC!��!e;kE'A���㨮
��{�>��
�P ;�m@�
�­3.�΍uC�<چS�n�.hVN��i����{��e�k6��F|�{�\tUl���9'	ܪZ�$d.ڗ  �ȵn��g[��^��5��zmZw?�
���)��c�X��+i��w|�
�0�6cV��j�C
�9��P G�:5����Āa`�$�<���p�˺���&���ߛA�y���Y#�ћ�\�u�W��ć�� ���)�Ǖ�h���}�������De�ڟz
��"�r� 	���a2�8G����7F�ũ�m�C��Kf�oC���N�x��P� z�a=�� ^]�����H��"�7�	�+Qo^���/~c�<�;���G9�����BT��k`��
̚+W���\4;��7����⺠��ְpC�%7��&CO��nEp�j|dL�� ���Ϯ:Dӡ�v����=B}�����- ÇC��zo�s���EV0Ԁ(i�'C���0^x�?�G���
���	�lX��*$�����p~B�p���ܯ�7t���9�\IO_�5�����5a��o�$��g���_��w�����Hu���������q.�C�������ʏɽa�sҹ�Ƕ��0����_��7P/uz��T�e�cF�[5yy�&L��⋩9a�'�����J���^/M9�Њ��gq�������y��qC	�T������D�|X�ʨ��wF��"�n��C6ޱc0����;0-� ���\��J�F�~��|�CЇا�?��9��v�i�z*��
�C����xtw2�Z�#�}J����_a��U���o��m_E�-(+̠b�x�䧈GlJپ�o��'`��u�>�U)��~>���S
��}�����r*�2a+)0�����w��K���+���u��mj���v7�X���#'��>\���ד{<ڃ��_B���M�>\� ��AFD�a�ou�~�s�.�E*���^�n���n���o���wÍd�v�W\m`9|>d�6xh��i]�ǘ�|��H��$[���Jr�$�z�b�0��`�FU�	*n)�P��k8��.�3.�N��J."��DE�**�9�S�r�b������E�9�!ٱ!���οC����wo�8�B�E�?�V�*Q�乨���z!�i��x�.��L��Z��=�N�FTd�?�!̃a.[.���x�m۬�:��4k����/�c�R���q�$��ĭ�S:�H��.r��E�D9����9B;�\�������*x#�L7}o._ai�N9q�T�ӛ0^��\x�e�[<��'U�[o�J�\���p.�z����}ݞ���ˁ{��3|)\x���0nQ�����3tf��+�g$�G8�jQ���ʋ���)��h�GA@����j�����1�J�+��8�P�XC���dq�����o��gx��=�g��=��X�z��0�A} ��LW�ܶ>��I���0�y'~#$�OY�fZ)=�{�^�;�kz?���?��e��+)x�W��rG�����վڂ:���'#�R�F�ܑ=d.�'M��\ı�+a����.�.�@�F�Ӏ�-�$F�c��p���9)�,�AP���rEsN����i�=-v:��Hw�C�R	�}X�������=�B��Y���g���xQ�E碽��m��pa��k����� y֊ǖ�����n��(�)��@bcT_gqg��z^�2���`�mx)���#l\%��@��7�Z�Wac'����'�ieC�Ŧ��HOG^j!܂�1����pC�a{L!Pxl�]�V%tR��o�m-p��'�]���I��F�`�蜬�4���X���q2�W��& �e%��hkA/Ž`�]L��c
a��|;��-��*M�����}��I����7W�寄U�Ś�9������Wp������\�?G�Ԣ�t l�I�[l��?�{�k�=
�%<9���-�ݼJ���;<(��~x	@��de�@?\Ӟ�L��w&�xW��J�'�{ �����
aA�[����3,i�౭x���ԓ��,Jv�"X��zS�<�;��~��g#ѫ�L`Q27&$(���
�_����0KaU��g�9X<����9��l��:хt�٧έ�� �����%�@ �+����+ZQ���0׭������"I��N�N�3R?�*��m�t��71O���0x%��w�E�Qh�Ӿ�
<�g�̇k���-�0��w��w$݄�[G�u����%�L��Ze�8hF��q��u+��ˡ�v��,���ef¬?���eg�1�k�Y���
���R,��"�7�Y�ۛ"�,S�İ��Z�J�^;��V�v�b?��i�X�h�m�Ǎ�Ͽ���y~^�ޱƎ��f̀>s�8���Zo�G���Mo�|�$)6��J�}�Z2Ĺ�O��΃���k�_���^7�E�O��F���/1���:>������֥�m��1jo�k��X뽸��U����3���쯂>v,������:*���ll9H۵�r�*��7���F�FP���Ӯ�)�����n��\�%`�(�?	ۏ��\�&���L*���β�����#���~��3a,]B��50֮=.K�N ���U�gn�w'��f�
�{pN�����R8gk`(�(#�*��	��е$�sU��/�8��~�[���YsK�V��[t�L��g9NKi��9W���:�W�l���k))��	?FKNr��PXUm���A���J)],X�Z����3lZ
���3��/G��7V������� 	�Ny����ϥ\�S���/��.)��v�,���oʹ�>�}�|j�D��c2��P鿎��Q��K}�(#�ňǡy�)h�N���p44 Y�Jt�MHq����/e@�`�E�+#]��z�ɔymj��V璡^Jw!M�d��/��{�>lmj�k9ٝ�4����lw�]���T�QN�\\�UcO��r.NSL��K	��L^�Ά���x�D?�ad�Y�����JX)	�_M�|��?a���y���\��Q�?�v�j��+σ��Bk<"@}�N�'�47��4��|�ƻ�����_�6�¸�o��1(�{p�;/'�yy*'���\�B�p"IO)r�b��*m�������d�w�1��);�������1�������fvՅ}�0��XKR��R%���b��Q$�"a��'����R��:�R
���|"�?%��)P�Ǜ������D��3�7��R %��(�58���(u�3 o�����V����CƢ�f��<aR�ߨ"T��Q��gN�]����dV*� �Ann��&������7�R-��6|/�q��_s���h��s���1L^�L��
�VQ�ӁӦ�C��d	���(�H5]g_�='g���B���B?�/�"��	�A��5^ܜe�'l�a�r��G<���jP����:b�;�<���>�;t(����}��β�����q8����.'f~��m�с��k֠��ݝ�c��Z{>;�DCĎ�����Q�6(��/����9�N�H�V`Z�?
_��Tx�8魭��;қ[�A9-�6#Swl��,P�k�e�p]��]��1��}	n P8����?!Y�y9��/�~�-�I�7ˆˢ�Y��`l��,R7��{_���s�ަ����[Hi��=��	>�+��⎌�#zO�8T
�I�~@o��	�H�s``�"���JH���"(E�	OkUorH�"�2�{�4(ERҶIHPq��G���O��#������������<95�i,,�$zri�9�Ϯ�:��#�������\�u�������1�K�`�hI�7�$�,�Hg�o�w�� qk��x9��gށŇ���Ň�
 �䒸�����i.�����~l��+�ˑz��{�n�=Ԁw�r�-��H�A�C����ᩨ?|��O2������m4�6�=|!(Q�����k|4D�M�Kfq׀��֯�ńH�R��GB)Q�)�(b�t4(a���(��3N�R�ˆ||����HPz 	��C �}Y�V��MlC�%C���t���|0f��QJVܙf�v�hg(�N !0��dn����C�^�mʶe(b/b0{�B��Wd� ̳�t��ǒ���hXq�b �=�����@�x�m̶���ً�"���2|����;�ۚm��񑊝@���g+��-�9۞�Rlg <6�����m��%�=3�����P������@y��z���Q�ٰc�q-\����<���^�x��������y�_۾4�J���)�B�*w�wT%a��ŉW�{<"N��%H&N���wc��6�%:�i�s�@L
�f�7�<k���N��/Q����޻W3^i�������r�N?hkGڢE(^� �DS9�i�4���C߾�/���ݻ�%wFj����&	 �+P�ƛp��	-+�@ða8r��0++�C����(\�&���p��:�_q6BV}���/�����.#����ƍ�՜q&p��޷�[�d���>h�&�¶�\T?�\'Bkmk�ݓ�FUY���=~�(�C�I�"N�g������6v��v����{D�	6:K��.V�;���a�y>ũ��d��I���d؁�?�#�������9�a�H�����,.��>�i�ٚ�9޻�A�{�Y?�G����>Z���Vu�ٲ[)E�]{/���߻������C��/�b����ҳ��n/~���ƞ��k�U}�
���f�9a�����ٳ����<x�п8��ӎ���|��`��^Ɨ�������Z6� K����kŞ�����O�z������A����+��o�w�S�q�$dnڄ�;:�$R4���<����ݻ�������C�<�1s�#���zIa;��OqJ㟓�C��W]gQ�����Ν;PVvq�A�4��:�Mvuq��>�Pj;x����0��o�%�/r������VX���G�N�>������MvA�eڰa:��T�`۲�Q��Cp�����8yo �>Bl�nll�[�~�>hooG}]�J�s;�����֙�tO�7���O@w�p��Q>g�8�����`�okn�?eʔ{��׽s�̹��[n��>tX���9�;�xg큻�}�t4o��O���z�~��a�Q�75��������&���myA�K�À?��䷞r���q�ŗ0衇D�%6�9ZC���u���[^^^;���|l�ƍפ���tS�Nۿ�[�S�w���cp%�E��0}o�!�9��?���C�����/����ԍ�a`6"�����������#+κ:�W>yCe�a��?==��.��E�ͽvݺ����G�v����T�:�+�_��uޮp�F[.W�ܹsϞ1c�2��5��t��o��8L�\)��q���A��Cq������V��'>��C����j��ի��^��lq���/����N)�M��}$.��k�s����3G�1���k��6��1c��dC?�>�\�3�����2�TU��������M?~ŧ�~����|"o�ɚ;O���!6��7|���i����������-,�ֻ���#��t������ys��]JiX�hB�y� tj�W\�6l�[[�l�H���d<[�ܹ���@����{ZM[?\
/w�rTSC {���������_�\PZ:���v�P.��@0��E��3:���K@2(����1pР�6n��/�F��Ȧb㕿#�seHŞT+K'����=�]N�͜Y�a��������!��[��6�pݐGEFU���e��ӱr%J��uD�{58N��|
UT49g��NKO?�C�����(^�,F�йT��=��;�@�}�!����5��Z�}��T�l���J���Q���Ʌ����������ʞyF$�Н�Ia�ePV�y�M4�>��`_U5�����w���,�t�e��|��T�sE��`!�)�����N�@.5MgRC���;p }翝T�
>ۀ������Ta�o���T������;o�~p�ee�얂�߀��y�H��p�gwXE��%p��$��K���l�O���ԫ.Kb[�(*��&�8�(�8�s~�^w���('ѝ�cY�	z=�qb8��|ͤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�RDK�Ǹ��B���Y��_���|��@t���`����h�_���;Df��-�{�6q�f��L'�Ό'�[x,kw��ķ[���̦w>3rx���?~����n��la�PX �ݱ�K�sD<do�!^�[ �`������@۾��vq����jh�Q]�10֯���Ѯ���0`۶�����v����v�܁&�zZ�۶A3��qb?55���A�� (ގ�6+Qt��GKL
�[Y	�}p���x۠�χ��_��׵?���`A'�v���p�o�.+��[Æ��t�߼y�?t���>�A׺��f���o���+��j5l0�@iǎ��׷�������'p�A{D�^�����~�8	p�ƍ0�_���R�7��+�0q�C@�o�%Z�E�j��v���?� -B��-ȠD'�߂8|���@��5=l`��ȡ8'wY�?�ZH)�ރ�{��>���Y��׋~�wF.���y�R�(NᲵ G�(�R�I/."iU�λ"'��芖��U��{8�pE$=?�rk�Ĉq�k>s�[�?�+�tʹ��.�j�%���aC���)�����W�o(B#$N%�Go�HDH�~8w�\�Ë#N|�8q�+�xm!%�� ��?��A�    IEND�B`�PK
     t$v[��4k� k� /   images/fd3ac6b5-800b-45c8-a4ce-2476671127d4.png�PNG

   IHDR  �  �   ��g�   	pHYs  \F  \F�CA  ��IDATx���`S���w�)KT���T�Tq�OQ��P����7�� Ȕ%C콡�����ۦ�i���M{o���W�����m����;�Y�������*Y�    @��Hiu�7&�SWUA~�����;{�:    X3G'7v��{e~����.�۰i�T    `՜���V�c�͞���>l��-�    `S�&د^>�K~~���J��    `K�"د]�~ha�"v��m�7��    ���>�ϛ7ϱX��c�_�G�]      [$�`������]6n>@     �J��>f��Qi��/X���J̖    �%�`�rɜv�%E��/�H99�    `�d��-��_h�Z�:v����d    �u��111�E�V�;p"��S     2�ʂ\������w     ��U��Y6�����,�H%%%     �d�Z1�YaQ��E�~S���"     �C����z(��������	     *�|�W�T����{�|�]{     T&�`�|���iO�X��     @?I����z��L_�t     �'�`�������嫶�'%�"     0L��>&�Sג��u��8v�"    �q��ʂ�o�]��~��C     U�\��Y6�մ�̧-�DJ��     �j�
����w_Aa�G?.��rr�I�|}}��ݝ��ƍX�� ruu%�JHH��  `���E���(v��mNq�)$E;v�o��V��~�����������	 ��֭͝;����H�bcci�̙�  	�����SOQJJ
����'�`?o�<G�}Z̮?����4IQ�N��P���FR�������ѣ}�����HR6h� �=�= H�=��C'N>���)11�@�$��Ҿ�r�F��� )��H�6���~�m����ӧ}�ᇒ�����5k�= �)���1HW��5�f����yq����3���ݻ#}r	����#�܃M��>�@8�dذa����{  ��:}��Y��]E��y�l���l���z�>��c�����۔�-��9<<�
E��0r���������e�u�������QXXX��1r ���H��h���kT~b��BQQ%''@M�Y�����,�[����n�.'���}��7n�������iڴi��=F��=��4c�!4�:p� ����TPP@R���O�o�Q�q���ܻ�K�۷7�k�����^��{�V�kG�E�'O��{H�ߟ~�)-Z�� j�N������N+���L�����<��#4g��W�<y��_�������὾poj=���7)4H�uҋ~ʠ�;���t�y���t߾}��+�Paa!I���\_�ǄZ�����B_}��0P���?��5��N�y����������A���/_:�𝋴�4髓`߼�����Ծ+cv��<��c­o}������^zI2��uYk�wqVЧoQ�.$uS^�����yP�?#��Н+�g��0a��B��=��]�r��^�m۶B�Qnu�|�r�_å�����%��>|��y˿�ڵk'|�ȑ#��!>ץ�ZO<� �|�z�_�d΀ܜ�ɼUQQ���j8p �M�;ҷ�~a�OJ�����p�줠�ߖG�g�v
z�@J�L�#���Ț��^˓&Mһm۶m�-q~��2�{ �Z�f-[��������7�r��)S(((�>��3�����.t�cyyyB�T��U�VB)N�z��'����Pz��W%W �W��>fٻM�J��%+�(R�2HJx��w�����?~�dG�tYK�wtT���ck��������� z~j��"���3T�ζl�"��K=�k �H_�|:.����cǒ���01_�g������5y��θ���;q�I�s��I2d�p\!���{����X ���`���=�U%�6n��u��U�>�8��}�{�n���\B����=�|�;!��v���`�����S�i�t#�����7o.�;�C��݇_<����:����)55���_h5����߄Q��byܡ�@�������%�qf��/(33�|�P���%��s}zup��� ��ȹ�ˀZ�l)�0U�{���bͲ9O���b�������{g'G�̝_`���5��M����C�������73B�ٷnЭ۵�n�Q�F�`����^\��;;h��ɼ>����ł�=�f����ջm�ƍ��[oY�ի����%˝�� �a��;�I���|>���?�P`` B=T[����s޺�z{ಕ[IJ�A�n�s(���b��za~�8:���@O��r'���G7S3).�]��DW��$���Y�e'�Z����N�JR���/�S��d�:s^|'�r�-�����K�}���������edd�M��\q�J�P����6�[�������(2��$?�J�oFf.��ʢ��T�t5E8�����P�{����G X��\H��'z]�;���f�`�j٬��g��p��Kk�f���6a��#}NNtw�Fԩ]�:x����Ux����5���cW��_�)'�fo+V������?Iɫc|�ޞdMZ4r�O�ѫ�%�%����U�Y�(..N�p�n��2׎jƋ/��HE�=�>�r�J�={v�����#u�>�G����G�^n�[�����kK!���>���������]�/�s9�= ���ӓ~����>�|�}��F�ѴiS����Z�c��)�!�����װ��V���n��,���\Kǥ+5�����(��@rsu"sp��ѥ�wwS�{��=pF}�a�����.xv�T�<ڗF�&kԩ�+�H�|�wb,��G��n��򅜱֬�W��^x�����Ϲft׮]���ǅ�]Rƭ�j���NAw����[���y�/����ZR��Mh������kt�r����P� @Mq���
���ڵ��9O��9\b�s�N�X,�/Z4ݥXi���=�=Or�믿�(�{y�Ҡ�Pd� Q�GG{!`�n^�V�;@)��d.��I5�?7ć�<n��^�w7w��Q҇�Ŀȍ��Z�i���O�
���-�M�6	�Մ�wo��^xRoMB���y�>��/����h�>ؖڶl@�>Hi��_�����R�='���*�w�u�nݺ�{��a^�_��Ϋ�[�K�ł���ӷ�/�wذiي�_=�;y���s=(Л^|�7��� ���H�dX?/z~�ق�}=)%�XX�VLj�v�k�U�V��>}�Ї~h��Ay����]���Y�c��7��L/Z��>�|5�  ����ps~�Z0�X<Pd�$b��s�=����
qY7H�u���,�c��~�Vz���ne�. mڴ��8߆�q���{jX�S�������](v��t�tY�$;�?�%/��+qE���x��j���a��p~��i�2�i㒜~��Uk�k�s[F�&�c�¿��A���s  ]\%�u�V���f^O���_&�2�c�d���I�D�+ˁ��>f��{KJ>]�t#e��%t�҅�|��J�o߾�N�}`���ݢ�^�ܓ�;j�a�/����Τ��/G7p5�k��G�ڵk��/�(����`��`�d�װ����O�G�y�; �4.��U����+t4���V8�q�%�F�`�r�`e	���v���kId8S�P��8I�'�%�H�������8A��''�P��G����9�Up��ꀿ���2�,s��œ��C����pכ-Z#���/Ƈ=������J�q+97��JAA��E����Q8�C�BM�8pp��=���yX� @�g�}�Ya> 7���-�ϛ7�Ѿ85������M�պ�P��B�{U���K.\���8�n҂տ&�ۧ��<��|߉l8����h����3���N�t�^��j�>\� Y�׷�^.�GIz�!��;�L�����Ϸ�522s�/_IY�̧�~X�Q�=�����t���A�|�ݍ^)pל~};
sf  L%�dV��7�=��$$$�G�`���ٵ���׬�wW��V�{;5�r�sO���x`ٲߍ�{߰� �N�۷�;��~nլ���zϐ&ѡԬI�=�zݪ¼���f_�|s�_8|�py��^ƶ���thU�~��%�����kŊ����Z�rS��������z�7�lZ�~c?C�[ԧ��&���j�b�>�x��0�!J�_�t������,�d��ۥ�n-+LZ����ɫ��[�qXu��e�����ӣ��ӱm�������܅D��U����M����G7��v9�{M_���%�5\]]������/��|����-��Bu��q㿹D�>��G?nߦ�\Wo������   ���K�U�J~X�|3�J7�Ǻ��J�-��3�ϩ�q{��-Z��='�G��9��>!�>BG�KW���s��UT9��W)*m�c�wq�~�U��5m3�YP�5�6�ˉ3q���_�i�K��j۲��BQn��w0� L��c"�(]�~����(دX1ǗJ��~ݴ���k$��������n����,,��ϖ-[�\
�:ڵ�0zr%ܸu�/d}����-����<ٻIth3cߋ-�
!^O�/�؈~�?!�S�_�|��{//�j�+ְ��n��F�~=�f�?n�W�����_Ǽ9ap�������6�� `��g��1f��ӧ�9��V?u9������4h@�����0��]��Yc���A0>!��I�&�II�O6�p�Pǜf�Ék�t�V���J�~Z_��zP���5_���v��S�;v,���&O�uss��>6??��]�&���yt�Z��b=WRJ�����PIϓY��   j��`�<����i/Y����]�)4�������.ߺX��[��tP��)��D+cߏ�y����}���JU��C�B�_i��|R�7ܷmۖ>���8q"ݗ�n���jҤI�c�m�)7���gx�����+bwm����ܼ?(`��FQ�zg�
ߏ����N)#��Tg��^��w5Y��'�qxA��0+��,��?7�`
�,[PPD���[�V�~��!�s�gd/W������ �	��8�kz��
��!_��G��:_�P9�K�իW+|���
�}���&�j����S�N�5	2ޞ6-=k���y�v�Z��Iƾ'{ i���J}M������V5����A�Ν;����;��0U����%���(UK��ܪ��d�u��~��^����9�TvߩT�����F�Bm���|Ⱦ<���&�+��W�W�}P6@��XS�o����)Ő��O?	#J�����;���&S�O1���!G�;�֋���wޱ�?��JA�j��ϙ��?O��`���@�6m*���_�~��uG�u?���#� O�4�222�|?~<4���� ��V�����,P�ۺ�/��'/��rs5~K�@UxD��\�bKf���*��\�꺘�r�ܕ���-�)���U�XY�&:й�PR�ˢ(���ڗ~��E�w�(ߦ�����+�\���Qz�ɷr۴iS�צ��/*���ڹY%���Kn�9����R�.M��Q��\�8��*��o�֭�_�~@x�����~�v��M�ׯ��k��
��KgΜ)�Zxn�F˖-�n7�k����/�m�6�AAAԩS�
�EEE	����煁 �&���:0)b��^x�����m=H��裏����V��1b�:zT���J���W*��,���EE�`�����I�+�B�G7�k>���J]zO!www����/��=VVs_q�^�x�������>�F���5Ǐn��R��p�g�����Cre�`�\),*R-߾�"8��[��z���	��6<���9.\�@S�L��5�b᭷���i��׷t��?��s�z�۷o�̙3�$�?���4l�0�]	5w�9�/X���n�J -&���߼��=h���l���>�%�'��CI2O�� ��~�/*�����)��ꕚ�3�/i��=��������K����ݻWy7))I�P��>�����VW�\!�*)6|�89:*��!�~�Q���jrs5|�]P��/ ��Q�E����_e�1��������Էo�j?��5kݺU�s�BBB�7ިr?���#�|�`/=&�U�f=XPX����6PN���«Jn���x���mI�`?fLW'��
��Mkm(gz�gyiΝ�z��ɯ�>iwʑϨ=�	[;w������]n��s�/��|���9�{����;y�� ��믿ґ#�U����6TyGS���_�/^L={�,��d�¿�O�8Au�zx��v�4c����;�<��._�l���݀4��;%`�*�}̒(I�*f�.�����[�F�{���P��I��+vy�؂XU}O�D3i�bm}Y��rUi/r!�+U�{�Z~�|�<� -�x;OWg�gH�`��������u��K111u���2��c�ƚ5��ￅ�����(��FF���E�]Tvʵ����/�n�W)73��h��eP���b?����PcۓRn���3b'�+UF��:�G�Tou���W��{V��y|}<�cl{R��?  `��{W{�o�^K�v��;���Fr:�������3fx�qKVn�^��5��vQ�[��e8���"� �=��T�ʷhde�Q�,�-&���k��U�W��|����ް~@���Yy�a  �0�c��z1#;���J�Ŷ;1Ӑ3�{�0��=z�߳gO�V��#8�'���p�޹7l~B�6M��HDV0p�����k��'xq�\�9�@��m�wߥ�������3s&��td����FjlϜO    1�����O�R�����QF���nW��W���-�j��x��"��={�^���~���Q�F�9!�%P;�x�	�0a�h�k׮�ّ�W{V?< ���[������0�џ"�ۇ�   ��R�_�rV0S��{�/\�')�K�\���.�\�3r���xjռ��}Z4�wϋc[�݂�O��ό�;�m�����F�m�|5�@G�ұ�]xis��^􉉉5>�ڵkI�RR3�¥$jbp�V�����cK�_�q�9���G���e�'��s-.��lso  _�`�k�t��xŚ���k�苧���B�[]���)ux/_�Y��ZG<����g�Snݿz�N��c�upk��u��V5y��='��K���H�(m�#���S��$[�6�2.��Ug?��#rpp=5j��{Ћ���'�QT���n�x�6�'��x��Ԝcc���XzĈ�^~��[Z6�oUs�w�W�  ��
�>9���I�=V�l'�w�9���ҹ���G�4�I�qs�)�v���v]ӷߠA��|��gDG����r)ʳ�o�]��Y0��c���V��FQ��T5�[~��gyA^P�W
��e��O�E��B�2�_��w����y<�2�v�+~ު�����{�z;��8*�io/�*[	?u��\Ca  O��Ϛe���������P{%-r�#n��NA��F�sws�k�&rpI�rpttHZVN�����x�JU��d���� <�/��$Ym9����Ȗ��KZ��v�0_­HK[]rKҚ�s�f���P!�{{��\Ξ=[�b"�n��0��}=�����j߾m�(��;*"zhjv���}���빻9��6�����\�u�   &!د\<��J��q��-���~��QTTB+���<H��NU�oooG������Y3��V�; ��E��
a�*M-���?�P�R*ȎJ�
(��[?�
�(�Kt�F�5���ܜ2˷�-�����?� �{6o޼:[�E�

�h����ܨ���\�M2��mP/ @�!��7�9�w?g^���  ��aŊ9��Jպ߶��~�4nӛ�{P/]����äpPJ��b��i����n�=��W�?�Sp�/-��/������j�:_���~E���#�
��
Y|���o)*���d�֭���_��|�V���F�F��13�梜ˀ   ��`_�\��ћ��6}Mpg��w��!�����"�QXT,���o����4�S٨=OeVڕ��+�����}ݯ/�W�zͤ[��+р���Hs�Υ�m�
��R�o���p1�qg�E+w�ޔ;o����V�/ ��
  ,�Kq�n�r�s� 1)��Y���LQ���'�r��6}Py��l��0�΋uq�/�'aG����y_��������h��BɎt�Eʻ�K]�t>疖���)??��4��S��w���R�pQ��p���� �JǺ   `9B�=F���u�V�m#��m��͹F�+,,�=���?�Qq	V ��#�kF����p��|i�UY���cU(���ׄz�}�l�رԿ����x�JKC����)~\�;�ݾ��ޒ�\kv��(��?N	ݳ�{  ,́@t*�9zYhgש}����Y�cdf���c���_�)�쌪P���M�Jp�>���^�׭��j�������]w�Eǎ#�>����?�ȉ�ԹC#��.�|}ܫu�@�V��}^>�_  ���5������QtdE�� O��v��'���ʹL�V�ҕd�wSPY���*�p�YuV+�<��15
�R�j�*�ӧ�г�M�<���݅��`��������/��mP/@}�z���[��n_�v+�����KW��z|� ��!����q����z���Q(��=K���n�g�������;T����r�?y�$M�0A�Óh�����ӬY�l���O�>-�1��/��Mw��	.��aaa  `���iӦ	��{��!K+(��@��T�o�!k�	���4�\�A�>z�S��B�ㆾVj���G���}�����~�СB_�)S�Pa����̙3�222诿���s���۴iS���O	  ���7oެ��/���^}��Z	���A��`�
�թ(%ź��W���6�U�rc���cR�k�.a���5e9}��>��_PP@�B���N.?z饗j%�׆F���4]���l����  ��ܕ+�[cʦ����Ӆ�{�=�Tx���_|A���:�ܹ��o�s��Z]���_&9���~�tCթ�Pp�S�׶�~z�g���'ooo�=z�w�}'�{���5x��7���֭[Wx��=�Y���?�$9����������˞�IѸq�h���  �t�R��w���`�=��şKTtý���p�[��>44�-Z��6�ƍ��SO	����ڏ�{<�:~�8�5J���Ν;y/��ef�=���,z���{^���k9���
�o```�mW�^���~�RSS	  @æ�=��p�#�
�իWi[RR�
����9D7��ژ���|I-t<�+�#F�k�Y�6m�r����,[�L�k�����/��*m�~��p��+E  �f���Y[�����N���+m���?�<��ő,�9�ڷt��\,r|)���8W@���j�xŘ1c��?�q^~���#GJ"�3k�|�e���B���w�x12k�  �@�/c-����W��ѕ�ݺuK���\��+P�k�'��S�-C�+�&SNn���˵�\�<`� Q��}�v�k	�!!!6}�i�^>�}�c  �ƜAX{-r�<��C��P���.ܾ�x�"I�������Ǟ��X�Ur��� �R/�3׼y�h͚5  ��`�C����ˋ~��jܸq�m<Q�'LJ1�kX{���PoK��|�[ZFEEU�&��9  �.{=��===�P߲e�J�8�p(8u�I���{���%�p��s|�����b�  H���.�'v�ԩ�6��}��$����B�n�a���B�?q�Ʌ��{�������wnp����%���3�#��B����  @�����&����"V���-u��Σ���\n�%�#��-.A34r/�E�4wښ4iRi���ĠP(��Ύ  ��~��T\TLP��͕�����#�����>�΂}��]�vz�]�|�Μ9Cr%�p�P/<r��]�-�0:th����Oo�;w���H�B!��� �Np���P�� �T*����߄	�n����+�P]ٿ?M�<Y�Q�w�q`��J��p#Gr���1q�D��>;v�Ο��u�V��nƌ�F����;�\   0��\��/���޽�^{�5*,,����_�����J�m۶B���>+���r�������G��w�o��Fo��Q]Z�v�p�Ξ=�*�:滄\���/RNN  T�^�&MV��g���4eʔ:<���̝;W(�֢E!����۷I�8�O��B?�
�&�N$U�!�K���=M�>��|�I��ccc��w�z�K��M����D���܎���\�  `���%Ρ`���z�oܸ��~�m*.�ք�?��C����W_���s�m͚5��K�
���͛$G��:S�pG���aԱ���+��np�������z��^�Z��u�R�e��B㣏>�t�����9w����9  �{-
�{�=0`���j"������{~��nnnn��j���������w�ҧS���Iړ�4�@���M��:�w�>��cz衇�n_�`�ЦV��m�FB�-�;o<gf�����+ײ:  �<�2�Bʣe�z�һ]�@��&�~������^a�j����7���$r	��u�;���*�4�OD嶵R�eu�Ǐ�[V׼y��93��  @�=�����d{��w�\B���Ç��=w��A˗/���z�H���5�kߝ�P��%-���;��������"�w޸�nɒ%�.�  ˱�`���h�Ν+m�P��'���ŋIn�9"��sW�
���p��Z��ő�5�k ��///ar��E�xB�̙3��3r�+�r7�Ӡ{������{��y ��a���C�js[H]��ʕ+-��v���@v
SQQ���q��)�=�q���������\�~���s[Y�z����Z���U����/M�:U�sI4������M�V�ơ��6l��s;8ؓ����A�R�/��q7�3�{�-22�����-R�� ����t�牲�B=w���7�G��� �ES�z�M�n;���Rڭl��J��$o�%5��,��s����p�w+���GR!����e�5j#�7h�@�����x���z�sKH)�i�B=��兩�Z��NA���QTկ�OA���Z��=7��RӲJ�߫|���ra�]V���Ya[Æ����z�\�sI��E  �ʦ���%����=�JYS�.NԹcc��.���ܪܷ^���v��M(/���B���̬�}gϞz���;�����KRam�^Ò�>((H�h+�k2�RSS���w��	O>�Q5����NM��]Q���Zž��vg�½�=�('��+=�sj�r�ѣG�nW�u��~  �ͦ��><�_�P�#|��}����ټ���PѥsS�8���`��S5����E�f7&&���ZC��%�=���
�3�<(,�T|W����Б�W]�p/՟}�{�i����.���R��`ޯH�#���f��ƴ���{��?���q�._�  �`����b|��h���Q�pqFP9d���9�jV�V�|�n$���.11����C����!��믩q����'N�F�ssk~���V>��s�^��w���oݺ�䠦篿�������BĹ�ŵ�|�ߪEZ�v?��f�},���   �"�0?zHwa�]l8^�Ů��N��f'stj��AV�54�~�G7i�?�p�/�С����˗�I�b�zƵ�<q|ڴi�J�<)��>�{[���`>���wٌ	
�q��������7  ��EcG�NN���+�N:<��n�==q������l&�kp��y�[��}׮]��<'��o߾Mb�U�5jDÇ�y�v���G�ЈA݄s�R�wÈ�])旃��x  ��������,�5�~���:Qnn����?[�`nܰ����k�����a�X4�kpi����K�W�+�R  @L�5ē�?y�ɷ�
�T�7��s�/�ĩTT��h�������\e���:ӷ��� �p���'��|Q�_ ��q9�y�
�Jx�GG�wW����y�\��'�C�����[k�1  @�}��ٖ����O��.\J�1�D5eŊ-zg�����9|rT��)�A>F�cr{���D�V�&���u,�Uz<ګ�0�*鷳/]I���՜�{�d�ۧG�.��]�FG�����b�x.��Ꮄ�}   ��N�������O�~�P Ј�=]������i����nݢ� �3$:"�Z5�O'�X�dZ1��¾mkX?�ڶ�0����:s}��s�ٳ���:o�C4U}��n�O�ϭ�7x�K�i�4�G�����   � �`ϫ�6o޼��w�K����7��x���?,��lu�;s&)�6~zd��ڷ���X� ���xXZ��@o�1��;���y��#ǯ|�����sܲ�G��{����0vq���{@�  �H>��B9��9}�44�ꊟ�5oft�g�U7�k[�|���vh=�P �6z<�g�-��zsB���1��:�yw��9~�zluC���˷�tvrk�&�yC�����t5�&  Ԕ䃽T�ժ�p7���Ĵ�����y~\�y���Ӭqx��K��{� ����LO�
��4_��Ϫ�1��vm"�n�r-%����y�-��¤�lb�f�m��   
{35onp��\�~󕥫��5䵤�f�ot���Qo�l�8T�å���(�&�W��P����*��J���֣���ϣ�7o��n�iX?�GG{���wɆ����  �������D!�>�'ܸ��t��Ub=߲5����>޴IX[}۝�),ć�o���PT)Ы���zh�����4��q4#�R�xTXX%&&�~숈�F^�����ap�����˷m��V���7,��b��F��{��P`�7���   ��@�7CP���2�Դ��b?g���e�wmm	��`_��F�(�J�q2:�XQ�eo�{**�{)�ݻwS�޽�9(?���5����E;��!Chذa��t���|�����A�缕������`  5�`o_O��ss׈���	���C�~ƿ'k�/�k�J'�k�W�p�W�n���4���R��o���'�{�I��==��3��S��z��Io����qII	M�<��;F��������<�2��3+7�G2�m��  � ؛�W�4�HQtD������n�tww��;��Ŵ�o�Nw�^_�Wjz~��'��Ԑ��TT�Ps�d�J������{��B�/,,�	&��ŋ�v��Z���s��֭[kt\777�����̙3iǎdM�\�����-��W1��\�ީ����A�O�����  `Y�fp0җ��AQQ@�%�7���H��m341���J�H��?7o;S�^�����c��������C!�Q���lz��h���B=�=��#���/���kג��w0|���o�^��z��_�:��}rckU   �
�&f(*.1��ßCIr���b?�����a���b�%��z��^y�c�9�F4��%:jϸ���^�+VP@@�h�]�z5͟?��Q���G�ǌ�d���b>���d���l������_  �{3������ҞD����suq6x� /�����|^68_9���fvU�H-.���iܸq4m�4����N�<I�f�"k��k���/�k�~�K��z�w��Ά���U�;  ��fH��mt����p�;Q'�z8)��iiYd�4���u�Z�^Y��ڇ�s|~�}�U
��3gΔw��Ro?W]�&������K5��   L�`o�����"6�(�>�������~~C�m��"j値U(á;�����*M�/�J2����=X���wc}���������mOJ���  ,���E��t��������̈>�����7|��55��K�J�iuɟ)�G�}*�@
��%;'�n�fPP�������G�5r�����x��Cz�nP/��������n�.   �)��t�l��`�"��۷�7[�l�q�l�����t�8{!��"L֬|�^��V�S{ԾfOB��2��'�|!� p�A�V����ik�z�����u�\  ���L�O]�^��6\����<*���5y����[al��'��-��N9�����]���s%$$X]���ǯR��Z��盞�S�a��<�K�>��a��c�9q�   Ā`o&�}~�t�m���>͚������~3�W�٭v�|v��_�jQ��}�o����Y덌?��\]]k�N�8au��'�������}Z6��}�3���~��'�y��zda�5���	7n  ��k`׾�Բy=r0�b�M���'Mx����׭�wٔ���7�������SU}��{N��o2iWi�����F�����&�B��N�	��k���<y6�ZF��v$�rܑ��

u�ּI������{N  �X�k 5-��:O=�knt�F!a���}}���f��~��4>`@���>��5����VeC�������$�u
EY���0��
���.�/ݿ��ԠA2Ղ���S([���5�kz��M>>>d�n$��_�/�=ݯIth�za~q>��ϸ��֪u{���oȐ���\�W�?����pQ}��'����T  �}��{�ESx�����\�w�n��:X=ܲE����܄⢒�)��<���CB�}L\`(3+�����:�*�/�sUp�/}P!l�铐�deeѩS�Lޟ۳j�Ϝ9Ӥ�iժ�U{�m�q�jdp"�����k�&�q�R�x�&�YY���E�)J�O���C�:ȇ����s�+�v���  �	���JJ��z�za�C���R��:C�}=�o�ԟ63�9��K�����j�L�W��!�y�����p�Edh.���J�4y�|d_Q��R����s�Z�EŴJ}.=?�Aruu�r�y
��j����9���rW��Oy��   &{��ے�{����ȞE���B�M��/-�)M�&�
a\�>/�g��%�Za�Ғ��DoG� \j�({���{�v35����KO�A�Ύ}���Z�O(  ��Hn$ߦ��v��!�����"ϑ_PD�~�O����:z;;^rV����ޮt�*��?�J��T*��P_�MQ���z�%����篧�e����2�?  �%H>����+=���OR�r3��Y����י�5#1qK<.���JSO_�9��W�����\�	��ؽ=�Y�Vq�X�h}Y���+�ϵKsl����;h�=,��ۚ�
mr  ,E���ٙ3gH.��
iy�Ԧe�ӳ-y{���x����?��X>tB~Y�no�	���@�*ߩ�1e	^;��i�ڗ�|E��딝�O�WZGP�ښ4o��߱��}�ͮ  �G��^�xe��g�]���]4���V��o�g�?G/ӡ/RAA�~��T�����l5Z�R�q.T�=:�/�k���V��*,@��(��}t�]stq�>���$L�  ��T\R"���[P�5�
���)P����k�D=~���ʣ�i��&��s��*��/ou���z^�������?Vy)�Bq��F�q��z��������d�i��ԟ�\ނ���qt(5��O����K}�:����Ŕ���>�����W�19  ���'��[ޙ#%5Sx;���
��֍[���e;��}��c�L�--�Q���s���7Z����b̘1�裏�֭[ɚY��M��!������Ѳ{  @��u̚5�����҉'�6�V(

������Qy�K�ҙ��	��h���+��+*>���B�9?%%�-ZD���?��_~�Ν;W+�W[�oxx8}���  `��Z�lM�:�6n�H֠Q�F��w�QX���z�R�9Ze9B/��T�=�o�X��w��������i��ɴk�.�mڴ.��w  �16�.]J�[�&7���k���|@4���Yt��E�sw��[�������[�+}�^��N�U��i�����Ҵp�B�={v��>����K���h���$g�z��?�Po]QQ͛7�   4l:��޽��.�����
۸��Krx�{ʔ)TPP@r��O�;Ｃ�67//O�ܹs'ə&t���k�qS���y�f���F�*l����I�&QTT���{B��Q�F	�/��#''�&N�H���#   ���4l�0�;w�p�[W�>}���u�ii�X1�/J^|�E��D��7o
��'O���7��&��^x.�����o���͛W��������+���۷I������>�����}��E  �f���q��!<���c�U�΁?&&F�R_,�G�y0w@ч���q��ƍdm�ø9�S��og*i寙�HNN�ѣG�G}D<�@���۷�U�V�K/�DW�\!)�2"� |������2|�.�A  �]�e
���]�vM 
��"��KyR�)�ꫯ�C�z����4a�I�2߱?��=�A���j�����RҋӒ��B����ҫ��*��;��v�/Ój�|�СC$Eܹ��<�h�B�v.�����|  ��^O��ɤ<�ǣ޺�4���m��$%���z��[���}�]��9�O�g&ї����Y3��S��t�2���Hx28O�������~������	�k֬!)iܸ���P�*�(�I�J��   A�׃'�q���o__�
۸��G��ی�jv;w�,]|���_����I���)�W�K��p/�PϸΛ�ٳgINbcc�I�򽼼*lspp�iӦQϞ=�	�RѵkW����̙#�  T�ހ#G�А!C�Q4������\��[s��c�g|Q��<x��*����Y]���;Wq��.+��  ��`oDBB�9�>��Sa�^N�nO��S0��p/�Pox������м�╂y���'� �� �W�'�rk9�4�!A�Ƙ�g�w ч���w�i�4��{������>�,͘1�@r�����嶖   ա�����(�F*�~�:W�L��[o�]�I*�;&��KOO'�:vV���ҡ�'vRm��.n))W���[�6���Tp	�k��&��U   �P6��������5I��q/{�:W�5�����p�M��^rv�ӧ����@orr�h�Jr�T�>�Z4t�����^"�s,Z��ڶmK��{�s���-[�L���Ӟ={��   �p:j������5rh���������@|��B>��$w~�D3^>:%N�sEno
�w��Q  �VB�=�=��̜9�~�a���Y���   �W��Y�{ �ؾ}��f����t��ͤ�Y�x15i҄   @*t�A��B��222L���   �R��%�=�x���=��_c   �Ko{�{ q���N��/˷�(   ȃ��)�jki��);WE�cn   ��]y�j�����\�3س��PQ����lZ};   @u9T��=X����>~3���7س�G�R��h�z�{   �� �,��NA�N�{ڹ�-?Ɨr�nk   �ɤ`���^�C��N������?���оj�[��駟���   �dr�g� ��Q��������T��~����   X�j{�pPs
�N    u����!���=   �ͬ`��̇`   b3;�3�{     i�Q�g� էR   ��j��=@��   �&J�g� �C�   ����=�i����}?~<�X��   @�D�L�G�C��/�=@e2��t��1;v,  �<�����s8���=�=ԊLE96>��M�/<�~;W>YUU����*����`O����p��8    .�{6xĔ�6�:4#�׈
�e�\CiI'�`_�Fe]iTz�:o�8+�ݭ4���:؋� �  ��,��=ԵK	��t���h��&k��B��@
;Y�+%�=   �͢��!�C�ѓ�vvԡS�j&-q7)�ǲS�P�c.{   �Ń=C�yQ��Yj!)�z   [�{�pu`�R�yeY��Jq�  @\���=ȁ����^e��\)   ��j5�3�{�M��r�.:��{   [�{�p�V�Ӓ���    ⪓`��A����[pT�    �:��l&�  ���4�3�{��ܖ����    �:��$E�	���   ��D�g�`	��g!�+,7��\   b�L�g� 6���vlYY��J��99٤�S�o�T�G�   �I*�3�{S���M�UB�^Q�?VR��S�--�����7��F�1y   �&�`��A4e�4<ϩގS�Pz�
��eK��J���,Y��\   "�d�g�Pm
})J�=�w��oǣ�����{MW�b �   dB���!�CM)4��v��8�e#�L�RT�_�s=   ��$��=�T�@��8���BU�5�˪TG��G�����   �M���!�C�hFޅ$_Z��_U�����
�{��o��   ��d��=�Eqg�lYk����|_R��8    #�	��޺��׾�C���/�0VQړ��즪�e��Ŕ�Qh��D�vTڊG��   �"�`��W^b6)�k콲o�$i�J� ���.�Q�C}����l=J�}��   @\����Cԅ�z�H]���8���"7j�  @l����K7L�����C{   �	�{�pUQhf�R�қ��
${   ���=C������{�
��&��[2{�`.   �>���^�f}�J�������Q����
��    &���^��n��S��wC�1Y�W�iIt;KI    b��`���)�f1�{'�v��M��   ,ɪ�=C�����b"+.;G�   K��`��AJ�  �6Xe�g� i���   P+�6�3�{�k�l�F�  �Za���!�C]�/��    )V��=    X;���    ���{�p    �ʦ�=C�    kds��!�   ����`��   ���l�g�    `-l:�3�{�����   Pl>�3�{�����i��|��g.   X�}�{�;;͙HӿH������FGGSϞ=����t��I��ӿ:|�0���   H���{�{u��9!�
mٛm��_�>-Z������瞣nݺQAAA��ӣG�3g����ȑ#)55�   @��u �׍'�x��/����������*ڼ�r#�������
���;w�����:օ��z�P�7o=��S���E    M�z �׮���1�D��;4r��>>@����̞=������y�}���TRRb���g��5k�P�f�h�ܹ����SQQ  �� ��p_;���	O���Є��"�~@�	����5f̘A���5:fBBM�8�,X@w�}7}�����믛}�    ��`o½�u��J���}��n����p�<yr��7o�]�v�r���K��;v,��Ջ�N�J3g�$   ��* ܃��?�!W�ҋ���\�裏D=>����׏���h����n�::q�  �t ؛ ��k�SRRD=f~~>:tH���o  H����A.��%ddd   H�}5 �[�	}5���eg��+ذaB�����M��  @��	��r�\�J��d��h|"���������Ua��<G;�myyyU�ӨQ#a�R���������)�  ���`o�{�pu'���g;�Wz�ù�@o,�kF��������)��H}���ڤ0�VC˖-��vvvB�{S��Je�ˇ  X{3!�ˏ�\��Y�VA����0˺��T�O�&M�?�e��eU���	   �����A�uC���/��z�*��d58؛�  @��k�^4�ޔ�xaE��IVǎi�Ν��~�V��?�z{Sxzz   H���Ae�1�*՝���(�(���0ُ9��m�FG�ջ}���F��t�"���/<f@@ �w�}�   H��H�%J3y���Jg�^���������zꩧ��͍���i֬YB���dõ��Ǐ�𘓓͝;��N�o߮tlggg�ꫯ���G�<66��  H������5:s��ҀnbJ��8NO<�,|�\:�$$$�G}D3f�>����iӦє)S���W�}�����^�{PÆ����{�B�wuu�/���ڴi#|�c�z��r   ��^d�W/{���zoK��晐x���(����>#��5;~�L%���ެ<�޵kWz衇�����/L�MIIF�۷oO~~~���Sk֬��^��E������-l��v��Qxx���СC4i�$*))!   �{:j�k��>���z�쨔��"��Bv%���Ttt4EFF
�s0ׇKtƍGǏ���Lz��ׅ�������#�T�����B	Oaa!  �4!؃�P���	�Q�z^uV����٬�,!��X�B��OQQM�8Q�lѢEt��M�9s���׮]�^x����	   ����Y�\!{��e�Y||<�3���n��9�sY���7ұc��'�j�}}}���@������-   iC���C���sH��^p��U�:��℉�    O� :�L_VcOh�   2�`V��\�%8
�<Kq   �6!���Y�
   @�t����Z    �@�    �� :x�^��z   �{�j*���>�w�������p�t   �`V-",�\�W�R�&Ö���,5�ʪJW�e
����G�U#��79���V�m߾=]�~�>���r�
  ��@����	��0O�0�>�W���,�(�(���ή4�+x�L��ԩS�G>�������OEEE   �����2�
r~��:�������CY�W�z��)��c��#�w�޽��4���s�   l�=X�	���7�9�����$�
����   �{ +�p�B�Gc�ΝO   `;����U�����ԱcGa���͛	   l�=��8t��   �	�    �
 �    X{     +�`    `�    � �=ԩ%?gR���hC?�9�JZ�5�    �dCq
���#y�Ɯd�dJ0ق��6;�N](���=�H۶m����ڬcxyy�'�|B�6m����   H�=Թ����OShٌz��d�

ա~V
9�o���ׯM�<�
�7�,X@yyy�>N�.]��Ν;Sff&�ڵ�   @��Av��Ky�*rw��`_T����w�nS��~eߛ{3n�� l(-�-��Mh!�a�e��� F�*��7��a�v�#!���ݶ>�G:ґ,����mY�u�d�9�y�9�]��>�"�·M7ݔƏ/���h}!R�p��駟���ߟn��7n}��'   �`����S�0ҙ*����5��}z��M7�x#��׋�<�w�Y���]z�4x�`�f�mhҤI"�gƌ   �����$u�.�eM���R�\t�E4d��x���t���WY���3�<SD�@�'O��;��͛G    { ��O-���Z]���i��h�=���s
N��{ٲet�嗋}4H���N˗/'    �= e����QV��Z����{��?�Y��s���?�\���9��Yg�6m    8@�>��H�)5�[�b   �`��ፏWS���������#�P��Ü��s�x�xy���?gΜ�엇�   @p�؃�p�_3��_O:�t�|h��貪w��E�.]���;577���/F���   6{P<��
Z�,I��)�,\�I��Z����𓆳�[Xi5k��&͜93�6����/    �؃���SW�M,˹���o=�+�   ��� dt��5�:뮻��xĈ��۫W/   @p��2���s�ѣG[���}Ϟ=	    �b@�8��C饗^��!�E^M��d�M|���   ��� ,Y��z�c�<�H���{=��ӟ�D��	������{,����_�Ýh.\H �?}B   �b@x�'���H����J��}���X���{��/���;w.���i�m��4a��4M��s�g��ٳ	�ba�G�l @! (������N�s�����|�馛��O��ǌCg�}�c��������z�t����������կ�n�=z���t���o�A    { B3��k��ͬ��Z��/f\������s�=Իwojll�L&i�ʕԽ{w����"8j���    �	������ԙ?��Y�����G���,�Gu�y�4h� �7o���������#    �= !c���Էo_�y�=_����NR�L�>�ƎK�\sm��6i�?��"�    �b@�����~�ȋ����E���(7�{,�9��Xc�-�3o�<���/E~=    ����c�/_�<�mX޿��;q   @��      @�     {      B �     � �      @�    @M�3��-��[�n�b  �*$�I1�  �˜9s�L�������z4B�    @m���A�Fד�i�     �0 �      @�     {      B �     � �      @�  ��v؁���  �?�-[F�?�x^�@�  ���w�Y�   ��ﾃ�     E �      � �=      ! b  �����[�r�J  P8�/�{�=  ����k��  ���      @�     {      B �     � �      @�     {      B �     � �      @�(#C��x<Ns��)��F�A����p�B    P�؃����k��;��k��>��>��#��}���׺3f̠�S��ZwԨQ���S]]M�2�n���b��=�\:�#h���4f��駟    @�a�M6��o������k���v����_��WY�k���t�]w�H�t]�	&�}�ݗs���S}}�x��f�Q�l�喤i��у����   ��=(;[o�5�z�Խ{w��t�҅���:M�#х�����F߾}}o�b}��g�mn��&!��xz��%*Y����o��d2i-�W������Σy���_n���_�B?�0M�<�   � �e��h���V�SYX��-[F+V���L�nݨw��ԳgO����Xͯ�v�m%=�m�ݖn���of�ܹ�駟�����q577�卍��q�xn���b��q㨩�����JJ$�c�������o%��w�!*���C��#�[=�����y�AѠA�跿�-�  @`�؃�q�G�9�#}ժUt���ӓO>鈦z����O��O>Yl{�)��ԓ���*�~�s�=ž�U���C�?���"�',x\p����cN-���T�   D�=(9,㧟~:{���W_}%�8*��w���H2�Qe>�`���R�G�3q�ᇋN�\y�5k�8�o������>���m�hCC��"B|ꩧ�N��x>��Â�Vp*γ�>K   @�؃����ZR��+���f�r�,h�͝h�=��C��������W<XY�9%(_�~�m:묳�t�m��F�.p�(��3g�
    �bJG�y�Ѝ7�H����<���E��Yg�u
���_t�E"O��k���������k�ђ%K����    @)�؃�p���d?�v�B.���~1<����V
�ϟo�=w�    �&{x�������R��    PM � �����1���ŋ)��6�z�`�    �&{XxH��.�̱���?�jÝoyt�^�#�����X;���L�=�pK	�j����t�R   ���fe�eN��������&uuut�����k�w�}G�<��ҳ�F��v�m7Gꓛ���_eZ��K ���&l��-i��7���P����jÁ=I>3���x8o�o�ܹ���Si~3��b�0s�5�Іnh-�1��<�̒LPU(C��������O
T���)N<��رc闿���mx��K/�T�� �]�ҟ�L8�@�����t��>%_�<_�}���3U��H󸤼�E�u���n�����ӧ��]G��NɎb�_��o�=�5�F�AÇ�5�\S<V��u�����կh�����7>�5�X�v�Y�r%�p�	��?(;찃�����O�7ޠ��
�z�1�P�޽����/}��G��O ��<d�q�ݩ���ϸN��	J���M{.=��k$�*�> Ȉr���{��Gs� b1�bZL�C�|����]��2��{�9��sKr�{P5x6�q��e]���?��**χz�5)V6N;�4��/��k���x����f�ԩt�=�P�~��s�ؿ��;���?/�}衇��7�|�����6����cb�`��D�	C�-����R�ʕ�� \�p+��E�2��x�jW X���}<7�MѧY�}�݇���O+�p!��jp$���5-�G�s�y2)��/Z��"��#�p���;�Ǐ��Y�f(-|X���;ebƌt���Ӄ>(�et��U���|����@�=�@��
���S�R�2ߑ���b�H&E�����΋{3���WI�Q����>ӑ�r��5�@�^S3D]{̖�8�R�q]�K��s�z�~c[�f��v������)S�:f�=�,no���ȥ紗��[Ot��!.U��ŭR���^zID��X����8�{�С��8��p�I'ї_~I�p8�.'#�<y��q�o��@r��裏�e� Pu�q4b�p!�	C��'M��Q{N�R��*/��t��G-���+Q{�/7ľ.)+�q˾��k�_ϼ�q�O�?��\���c�؃���n����������;ҟ��g!�οg��O*!�駟��W^��m��V�~�_X�x�Y�e�s�˙���F�����7+R_f�L����Zb �-�|��D")n��#��	�z3GH�|2�rdJ��7W$�;�
�o��z�k�\G3Rv4[��5C�㺺3�3m�#�v�B�n�阔��<aB�����? �����뮻������z�%�G̩V��| ��S:� k9����&�d{����577����#G��0Ýb�s��7���Ջ@���_��5m+��@ ����)����Z���ӌ�۷��'e�ތ����j�=����#pJ�3P�y�.So��o���转��k	#�>u]ǒ��#_���o~�უ�g�q]}�մ��{SP����/��V�Z%����Ξ����d�������O>��ϟ��{�0��r����[�G����[���?�׾�:�,Q���縘W�1�k�{d��p㍭����~##��7��uU�M���z�=(:�jv,�-��y,�Y�H��>�0�>&;ך��ܙV7�>lxQG����௺�@����oQ�=zd\�%��9�<�'��\�SN9����k_����M�\
�����ӛo�)� |���0���GH���h=��i ��>}���6I��,G���J��ݙ����0��d��=)#��q�;9b� s�ˤ����ɰ=�Õq���� ���s���\?>���c�M����̩'N�����￟�9��r����:JTTn�����d�>:::��SO�[n�E�=�~��7<�p�/N�����γ����{t�}� �t4�}����v4^F��w��c�˴1�	CY���N�q�����Y�4�UI�h�L��H=w�M$y���kqk��sժ��b�G�9�|ʔ)E���FK)�����D>�m��F�W�.j_~;�r�O��Rβȹ�<�	��{�����ȼ
���������� ��B"n�Ȇ[�y2+�{Ns����(H�_�V��
ڹ�[ՙ�/���;�;�;�ޖz�ػ�b>p&㠿,(Y�?3�ߔzcHV�^��9��s3�c����}]T�"/X�=(9�n�)]z����n+�Ӆ���b���Bָ��3��8O�>��}��֌�~�>��~:]v�e4f��afQ�m�ӟ9f��<~����_���ʺ�+F=z��袋.ʻ	r�-�̹�[�w�e�����HGj�[��w뭷Z7�l�dd��G��(�����~�̙I�L{�s�zsXK����z�1��E�%�$�^�zE�y�z]�� �2)�=���dZz���Y  ���v����O���c�=�;���H0�쳏cy�N����B�7�xc1�գ�>*���%e�s��x&M�$�+���^���ܩ���T�#���p~<G������9r�-,��W'��N		s��Ӕ8����8��}w2^k��D��dE���<����x�wO��'@�>�,���Y��3�/��])�cd��D����c]t��"�ʺ���j �\J�a�I1I�f�ZS���[�u{�'ym��u	bJΧ�~*�Y懳�q���3l����l�]y��bX�yB+7,�2
+�H?����L�Հ#�\r���se���{�8�?�0�qq
W
T8���SO���{�M7��by��Ư�k1�����irJ������~+���o�-�&���=��k�l��t/�ׁ��<�U6x���k���=��#ZPx4nq���E �?Rl�4]���N�)F��� ��b����k�Df�2{�2���*��C�AY�v)�,�G�Yι�'G�8B-�u�sN}���8�����E���	�/dmU�󞣿�Ύ,}��n`8�����E���i��i�s���H�ﾻ#��p� W
�M���%K����}x�[���p�'�xb�}j��s�J� �)S<n���^Kp�I����9��+>|^8e�+Gj�;)���9�ϝ���g�yƱΫ��*^ �57^wߒ��Tx�^ӐmʏڙV��$3�ٙ�j�2V,��C�A��xN{��
�/���^���l�2�
�Q�L����s9�x�Cr
Y��nˑb?��Lkk��'�|�
�#�K�.����o�b��RϢ��
\�#�8B���J��[o-n~�:u�H��[�U�M�&��$�Y��Q�:"�����;�>��C`�(=Y7e��b�؃���矋��W�|.������r�Z���]��K8�>�e��|k���g�N�9���������;�иq�Dk����W_��o�����<<v<���3G����+�^r��_���u  P~�tF��zZ��i@�qw��ø��z�F�(�� �e��{�Ο/������<ZG��|y�&,b\pm��F4{�l!ʹ:<r�5�����/�R����O<q�\��θ,���#��E�|r�;W���lpw~-)��w�)>���Y   �d�(=٩:�b*w|���Z
87��8
��>�j����pE�o���s� ���2��փ!�;�n�c�+O���    ��Mǌ���Qǽq�Ɛav����   y�}9J���3l�2Pw6�a/�џ��/��   ���Bg��D�Q�  5���[����)e�bB�:�,Ñ5�c�>�jt����:@��αw�T�犆؃P����N��o�YLz�����i̘1�s�~	 �U�^�V�u�q-���ˑ��   @ՁÃ0"���H��b   ����N��Aδ ���a�*    ,����YU#�kxo BO>�{   ��jD���g���PR��4�   0�#����4hР���y�|��c�$�zB*�9��  �4�F����o߾%=��������P�h���=  �H����<�+������G<�����mD��/ط�  9�,���	WGZ�?��2~=y�>+��,��  �,��L��u�1 A��R�=  �HP��VK�3�o���a@^���s�  zT!�Qm�	B.y���i��TJ�ϟ/:��%;�[gGi�<h��@L�G�����[z�  j�лwojni)X�}�	����Ƃ�[�r��|��	T�J*J�@�  D��c6�fϞS�����LK�,�>}�.�҃��7{   �%ӏ?G�L,,�Ps�����.\(Cr@X���{   �$�464P�����m
���R��\ JCm~�    �= �b   ��\r� �@�A��ի�9���ٳgO�����[lA����?�D"Aa����F�U���۷�����q����K��� ��2@ރ	�I��ȱ��=(�n�-�p�U=��cǊ[��Ŋ+(ll��Ft��wW���k/q�6��;͙3�  �$��k�
��j����b   2�U�ʕ�������;:&Tʱ.�_�^r/�o�g�b   TD�G�^y�$>�\�xM]��?:�|�xlɽ�|��Q���[@�A�H&��j�*
;�ù�Q��X�,��ݟ�(��됝�!]
}L>�{��X�\�4��烮�^��1�'�1� ��=���=��v�3�믿NQdѢE��;R��ҥ}��'@�@Ծ<�S+DY���X̸��Y��s)���/���y�O7�>�䨡��+���C�  �;Pb2��˴y�ٌcR��
�bC�+/�ħ��麙�c�}��[��kre���6�@�  ���~�XB�DjK}]�OI}�\f�h��!��ZL��G�uq������ד2'��i����C�  ��(E�!��H�ф�ץn�uu���cΨ��|���lXRoF�Eڔ�'�I���ä�	�e$:��t �     >���R�ެ\��.8�L��C�ˇ-��Ui�t��9���n{#z�GS�!�     >�beg�X<&��u�:Z�b9��ґ�4*Tztc�{   ����('TU�S�x�ȭ�R��{��4h����^���p�B�R��}(��J    (!���f��������uu�DR�����Sb��]
έ����>�羻���#E���  PS���Ѹq��/^L ��S��1�c	OT&���4F9D���>L�h���n�³�kbd ƜS�zl>2�5�s�'��u�.N��=$M�՛��h�=����1c��|���:::�f�����fGY�,YBQ�}�;;;	T�$��{�Ȍg��↎��C�E3���cKOx"���v�y7ek\^Q��gщ�����E��ݺvM_7�:���w�y���o?�K�.�L�?��s��9nO�XE��  3*�R�B��c�6-�m)��RR��D{��v�7D_,�Lձ��"�N�q���S�7+ο{�^T��G+Vo �    ��nL{J讜�~}�S}}�H��L��^�g�53�I�k��^�ٗ#���EH~�3���   B&�*-~��SQ�z���1l���Ï�G�wt�O$��v$]���J�Y͎�Q����z�b����y������!�     y ����}y��TWWgE�e�y������֜Z��kim���Vjmk���N+�^b�=ҍ[��J(?Nj��8UAH�S��	M&�@�    �b:����E�e��Ï�x]��%u�))v��ň���w��®��*��P���m��,G�;ĠF4^]��Ƶ?����8IQ9�V�	�=    @4름��p���655��b�"�,���"�<iF��M�cg%��C=��#�Fed��T9"�{L�4�w����׼��ܑ�(����    �B�xn��ɝi&��X���9��!�W7SW�H�-���-��U\y읝I1�oRw�LHԿ������n������DWQb    PFX-9�#؝�VԞ�q���Qb�uo�a�g��}�gg�JL��N�(3Q���ђeK����s{wߚMV�R�|�
N �     e�'��aX�9�<�C@�ܛkP1n߿_Z{�5�q��D���n�L���ͤe˖��$^>V�k1cr+���ѪU+i�m	8��    ���=�RRςo猓=�;��<+�k��k���G)/(�(�_S�#;�x���}��Q��aYU���9�u��K/P{{�x�+�Hb�Bc�F]�kgj�QK,�G5���u�Za��=��JJ$q�A�����C��4�O:#�F�ɹ��:ݺu�79"�����]��t�����]�И�W\��,�K/�������:{���6m���V����=����7Z��n�t5u�������;����~��'N��U�H��e	��As��o�^M�d���šZ���u1���ϧ�Xa�Ck��3�;����S"���[,.^�`�D�M����h���z�@�'��҃.:�?�j�����K�����/�Gv��/XSR��kS�it�m������4��A4rD�%&?���<�,���9�h`�I=�׎=�>�ѥ7/��~� �9�&I��c��h:F���yUWs��<���ռ�����d�ӊ��K}=566���Q�Rϰ��~Š�������۱�M�l�j�S-��.Ɣ��Ƚ�[՚�3��[��#��~���~�]D�.�����>��L�!k�Lu��b��B��q�f�!����j��%��=�W���S��״����?ݺu%��=pP�R/1�u�o���1��}-K�$��9fvݡ����\�$]�ѓ!�1)��Z�����i�F���.;�ڝs�bXu�����Kٯ�s�(�C����ԃ���7��Ǜ6�Q}����Չa<�? ���֥^�W��$|����K��}��1� ش��QkkkZ���jJ},%�����3�&uR����L����d�Κ��뎔���ٕ�R�^ePF�a�׌�iE冋�z��c���![1d��x<Nu,����߯�@� ,R/�%�a>&�܇I�%��>�瘁�\X���ȣt��{Q�=�f��۩=u���)3�)TNP%W��x�֚	��'s��9�Y)8��f�J1>��S@M����vO�I��aObe��9����Ē��T �=��K2�}�����0J����S�$�瘁�\>��qs�)fu:xPJ�����FcL93m���g�Խ\���N�r�'z)�^ϰHw�n�\�X����ߚe���m���}�	��KXh�?�N�ؐ�(��}��z�qc��=�}T�1��V�觟������v�v;+����Fz{%Rʫ%�G�-E��r���H�)�������H=�U���L�*`��@�#Lإ^ҧW�n�b0�|�R:���57�e����Sn������'�����]���s̰�?��J���V eě��Gmmm���%i��tvv��-���Ev�]�=��W:�)��c�7J����(Q�zI��q����5x��(q�nME� X�!�����<�Kcc�x̫q��Xk�FOj9#��~��Όu�]&�V8����HI= ab@�0�u4F�!�C�x��jE<?��[o���_��!��MK`�j�zЬ^	�g����S鄨}~@�#�C�:~� �di�����5޼�����1�����ۭ��5i��i��zR_ {    �"Ft�b"j��bV�X#m��1�%�9|��h�Z}mW[��>�T�{ ���B�Ɏj�  ���ec����H�#��I1��X�\�=�����)�>���/��8:��#G��4�}�@�AE(�{ǽm-	o�ʭ��7��S�*)��i�E �h�MΠ*�ni�I9ּϜ��C�3-���U�}��wA�y1�8��<C��A��r����^�B �A(���@ ���Y�oD�E���e ��=(n�p4+�S��/?�{0��`/�*��5R�b��V[%�Zn �?I6b�T3��}>��S@9�؃��I�U�u���:� �$�Z���zp��K���ˠ�̹*1~p�˽,H������� @�X#���ΰR�SR�'��qd��2 �� ��������kz���rF�ZZ�}��H�^���&����Tf�_S�d�h�̥h����8����Ĉ�k�5 P*t���#�h���=()~��^����H�HF�ގ�#z�DW�3�U��Tn�d�y
5=-z_�2��⮨���UqQ)i�����  ʃ�m�҃2�eE7#n�5���ֹДsT�mѵ�st������ev����VˬVj�侚��*am�l�Q+kծ���%����|���r?Z �/  ��bAʕח)jm?w
��n��Mhʍ�۲3�<��W[�T���d2K�s�^���J��{�=+U撵J(�1���,x�^�u~��b�ll�d  @�@�A��ZS��ʱ|����P�����ˣ 'S��r/�#(R���R�I�W+6s�{*m��D�)�퐽!������V	�m5[vŋ�i�ȔV�Uf���(W��XI  P�@�#H֔�R��[�T��&�p����V�4�h�)���{w��d�X�E�*�cR�ZBO���ߏ$m���^�QU��/�U�qW\��>(��I��Z�<��n�����ˈ�(��Z    �=(3�%CnY�D$[ț92�+|-�72���Xʽnڐ��TS�S4t��ˊLң̖��"�F��^���)�V��QݴJ���&�ʚ�*a�o��|��JpټD��6GZY��Lһ̌�JTP����
  ��bJ���$�|[�D�9���7�=xHL���:i�!	RSz4;���OP$H��,_��w?���k�t	�L��2t��I��i�=����P�+/��Z%T�����]��V������z�j�y���R/+2vK�3��Z�FMTb��'U��y  @	��G�J��X�E�h�'���f۝��>>z{2�1x:�uC� �D������Y�u�_�O�>����[��Qk~b�cV`t�����3T�,ѩ�Mw�W���FIQ���cԵ�]�r$+l2��N�^ie?-Щ3A��[})2\��t@�$5t�QLm}�����
   ��M����J�nK�����]<f�'�QzwtW����~��Q���}ﯱ�Ί��h��[eU�6�c�tD[-�����7��k���s��f�;��z�f�|�
[P�e~��Mh�-v�^��y�~����h�F˽����
   �����(FޥnG�Hg@�4�H���l?�
~Z%���ԍ6�h��]�|9}��&"ݚnG��V	^�J�?�~�z�Uޮ�fR�Ϛ���_R�e   j�}��$����2��*1�s��Zm����F�s��~^K��H�+lK-  P�@�A�)މ4�_Rv?�\vL8F�t�������-��ɛ�)V�no�Uy��(}Q�V��:�y4�H ���k8���m����rI���؞�)��z�O%ڟ�'   �<@�#�^��^1�ՠ�s̚94��-�KKy)�%�^�V�񵐗  @y�؃���et,$gh��B��]e�ր��)�#[�aj��k�3����}>�ۇf�+Hx^�%�g!�   ~��G�J�Ɉ4�� y�b��M��)�ֽ�L�:H�܇��[O(��3-�e��i��gFN6Uо<N��s	   @�AYQ%W�
��\M��'_ѤW�l-j*M��3GF���)]�)���絸�#�\�����J������b^-��   ��=(	j���D�F��[DV�")��);�$ɨn�9�M,�q,f��\.�_i�uTb<Ҭ
#U��ٕ�@S�
��l̨�i���Vf   ��Rɾ���ƨ��xGn�S��B�
Ma;����ẉ2S	2噧�Y�oys���T�J��le.�#*l1�\���b�k���::��˞�yjnn&��A$����K/�I�  �bʂ��A�Ф�M��5uk�W�u��R���4�ޱĊֻ����l���-I��Oj�b~Ԕu��x��+�ZR/_?�ԣ�u�%;����<*0A�ش��C�Wiv���bϡ��������K/u,{뭷 ����A�iӦA�){PrTٕ��H��a��>�9��Ĕrk	P��6�=?�pdm0�sb"�I��2��gE�)]��!�^�㣋�tZ�x>����][d�M����iX�NKp�s�:�ՎX�2�k�u���Y��Fy�װw��.]E[�"��V�����   @�@�#H�b{n��B�{1�)��-�Cʽ�ԫ�y=�&��
2#ښRn���A��҄>��V���RP4s�#��K��\{v֤�|*}_V�Z��Rq��xC%�*���������z}v��JEM�������:+n���  @��e#��Y*��3^i����~ ����
�%�f��n��g*�5���_w���W�^�#�V�D\�'crͼ��U"��׊�[�)���En�R�\eR�.��#~O�g^�!,YE��G�r~�#�^r/��7)�^�����mRS��I�+]�Yn��ܫ��,�W����dk��O��Z\w��
�g��2��A)+ ����;Ĕ��ZF�u;�%ˣ̾@ ���d�{㉴ߴ@n�}Y�*���T$�Un��܏�8 e��*!��i����$�Y+k�s�Yfc{-�2�� �b�i�5R���ӧ9֔i}�6zV���C-��p ��,xɽ%F���]u� �^�"g��,��G��"j������H/˧��I�2P.���;"Һ�$;b��:�dҺq?�li6�k�L���"����+��'g�od;Hd+�����|�W�L���V	+_'}{q�V�Ld�ЈYZb<��� @��y�՚��;�+�L�'	�fʽ���o5{PV�t�#�����r�˥>��*�����5F�y�Uf��kQyZ���@��U~xM�,Ch���Y,�dʽ����N�LtR�#���H<(�=��h}���a-wTZ%$^���9l�v��X�yX\#�O,��_koo�ztttPGg�������V�}TPS�@�@�#H��'���[���*��(� P ,�)A�ҥ�u�����j�H�[{G;���
�g�oO�D�ތ�g����(�b�� ���V	-1�D)2_,.Ʋ!Ƶ����	H&"�����-������-љ0��k��u�_�~.��.a�� J�ח��aMknd=pn}�:INW��o]��46t��F�K��mFn}�έף%a4-�u�C��bA�9�D�g���h>D�:Џ��uW���(���7�r�*Z��,r�Y�F���9R/��d
�Fk�<��Q�=  �P�W�y����b��ߤ�B�YHCA�����_��V	K����h�j�6jo7r�y4�3m�*�Y��H�)�}��? �?�Q%bB�j�.ԣ��V�\�ab���������ya��ƞY�� �i�dw��(���5���1	��
+�x]��>���  9.XX�R/�ӧ�����d��+�jNZ�+��u\䪜Ɋ�kr��ې-Υ��������et�U���  @�hmi-J���.&�������X��|y�Γn�GoN%����NRIi�.;���3����4k.k��<v�gx\(��C#w�#W�=F9X���G�` @�ɖְj�*q���\�}��Ґ!C|�뗷�~��M�������
�' |!ǋW��r�J��z�H��3�]\�Z8� �Q~3�^�p�<�߸o�����B�{   @!W�3K�iu�B��}�R��k�t��+�u���o�}�C���~���׻�me�hJ����py�=-a���ޞ������}"Ʉ�  %�=��n�P�b_ʙ?�D�����x%�{���s�׊f^;|K�t��$V�sJ��t��Z_�ה�d?��H��"��5������"��3q��^ �� ��\ @4�#���\g)�^�b�3�兮�GS��\��N�P׍q��cq��jb�Tz1HN��3֒�ڢY��Yr�v4�-��?y�;�,�J����k1���fc���9�FN'＝���5�c��@�b   ��jPF��b�)�M�qo���a����;�,}]<)d�%7�ԕu3����DJ�9���Q�K
��TN���=�Nf�*��ԹӘ���7n�hOI}GG����W?K��餄1޿�#�gbE� d�3��|��ɵ����޶�c��6�4��꾊�������b�)�Is`��w\�h!��?м6��%݈�;/ig��W�s_��<rߪ��p��D'}?sf�ϚU�I&i��b���#��b   ��3�O��z�g����Rҽ{w_�A�k��y�X��.TϝB�a/��|�f��ET��Z��T���-*1F*Qg2A��	����\M���]t�]��g�EY.o�ٓ�<�\�:�5�oߥKZ�hM������  �����i�=KI)%"S��j������9s���dDύ���/��O��F�x)hf� �ŷw�S[K�ͦ���J7�$���T�[c���F�E�7����S׮�Գ�=�ܳ��[n�8��
>�>��r�s/�
?��w��Q�ܻ�ϔ_��.��7('��-:�1���Sb�G���K֞j3oۙ{ݘ�-i�񲄖0�#�ʦV�V�c؞'@��D�ez�����߾{�.��NQ�C�AE����jɬI
-3��w���7�>�����-��C�ˋ��ԞtVwXyss3}���h�7��򂘒��:O5w��o ���ԣT�E�qT=�H��Ug"&'����Br�������װ��+CZ��V����}y�744��ux:E��!��"[{�E��S�\�@�(T�U�RN/���X�Hf:��w+�)>���{_�߷���a9SI���)�^��h��������b����Ǔ�Hp4����3d��u�Ҥ�Dro�׬�"����J=��"�ڽ~�
�T���/��^����r3Ş�Z�X������t��u���D�Ant3Z/o^ttv�SO?AQe뭶��/�BD�9R/;���z�B�9'��z�C����Bu"��uN<��� ����I}�O]Zv��]��߳r�Y�3(�.�wf��J��w���(�x��\��׭�p��� �n/���=!�]E޽�4&��/�����ֽ֙�ݡVM�Q�������Ip��������Ϭf6�y�n�%7c���޸�l�+#��}W�ܙ.�|/� WZܔ��^�Au��dq����.%K�.�}��ȑml���Ff�/���:#W>�GJ�α�5��"N�D_Vj�fM�+��}��H�����	E�=(9�(������9��X��3.���{I}�J�3�o�)D��?����Y��.U����w�Ž���J�ʫ��4�Z�*k 7RH�v�J#F�(i��믿���ISVu�f�G.dʌ���~�a@�:��Th�.�)m�P]��p����zF ���d�zUnu���9'�p����
�q�R�%iR����23�+��� V� ��&W��c���\��UB=��Ŗ9H�5�?��Rl���s#�Dޒ�,[�����a}�i�*?^#LeX�^�U���]��ӌ�R��B��+r+{ѫ��Cҕ@��4ۙ˭H�)�A�]��z����擴r+��I�+)���J��(����{=����л��kA�kHx�����!T�YV���	8������.�nݺ�>,�;��>c^��|�O�ñLt��я{P2�Sk��r��m�Mi������NэI˕�O�U���
��Ie&J/w,f7U�����*�E�V	�H��������٫*�e�)v�+P��s.T����nk� �䍩���7߰žĴ�������G��	�%�;�k|!�gP<N:e�O[!d>�ݤ)�^Q�jD:sUf��'����-ʩ�sA���X,]�U�D�m� r��(���W��W���ΚV�g�ŽWy�=���"��D7?�B�y(�DBo	����ի+�~r�[���C�#H%.����S��DiRd���%M�ٓUȘ�W;�>[�E�uS�~��3�����M��*s��� (D�Z%4�5ƫ���n2I�u-���l��)�q�*4 7�zTjǰ��[BORgg�@�q��V5�=(	VD3�����E�8������i�?����mꠑ�;m�5m(h��j'a)}�Vi4}V��4hN����e�n���Z�R�e��=�VXU�
�o�m����|Z%�|r�3��V����B��dR/�̢��ۧ��V�B� P�XR��]i�G��!U�T�q���!E=�H��L�'���^���"�%�1
9S>�ޗ~�����o�Ak��b#�C&)���~��\�y���1�L�ӧ��������ޚ�"��ь赮����*A�JۼE:����\!��R�q�Ƙ����Խ[LH�Xϣ����,���I�ڤQXG��'Y�!b�P���'��9*�b��V�  ��G��7ti���o7�>�RO��BIR�ſ�ca���[�ݒ��U ���׼�ד����/�}��5!P��[���V
���?�{�Ϋ��Fd?�*��9*4:yK_����ǔz0��h�-��U�WӼ����v��
[��R���tz���i�-w󽟟�ͣ���iԚfz�����i:^�0h� ����y䑊�_�D]������ٜR)a�N�#�ֽ����-��5Ro�E�'rm��c?�I*�#=�i8�ޟ�Y;�]P����d;���l�J����~�/_N�,"�
[�Ӭ��.�sۧoS^��ҕ:~6�wX�=Ӭr-�*]tuttГO>Y��z����wJ��QjX�L�BH�(�\{)�|o���~R��f�&B�s�� ���#C�B^�Tr���n�)�����Ӫ��*�yN�����鈼Ӭ�c��)�מ�bT�>�fEM�Ye����DX���:���e��|�嗋s��SO���+9�G�H��d�M�,X@�/&P�~�૽��W>����yH�7{P1
�c���Ubt��(�}P���EԎ�Q�L�Nrlyr�Ø��Jj�R�j�[o�U�a}��'[�X�ǏO����裏RTa��<yr�Գ�w�q�l�2�#��5�,��K>�Ƭ�o��Z�!�؃�BG(�Zd��Vy�Uy�����z�9)��B�gެ����#��\0�&M�������K.��(�R�7�tS�r��c�9�f̘A�x�g���N�\�_LK3��bA�U�-��L�R(�m���,������d�y���D�ro��,~~K���#����{P��
��騅��bQ3'���є�b�@؀�C꫁�w�Y�w��=(֬;��-�r_r?A�ۢˬ)"�E��PL��Z4Nkň��C꫇���|��h>��>���(<���9�xKy�w�1g�Z�\�׫��aH�&���\q*N�cf���7Y��pU@`Sض�񝃆�y����G�3��g�)X��z:餓�ea��=z@�D�<{ 2�)3�S����؃� ��,�"Ups�o�	\�^V>�N�)`v%&��Z�j�ӘEQO;�ŵ�d����5	�K9ObV+�]i�
^k��'��(�=K=i	���ԃ����� bE��=$��b4+Őܘ�B��$2�����Ȗ�*Q�@�W�B>;�)ɍ���z��F�8�X,s���/�k��}h����NX�s[�DA�!�  / ��$dK�Qs͛��ҫ/L4�?w��9(
/�\bG;]���~U���AvԾ�{'���������e&r��y�\C�h��.���_W�D��$g'p�e*g��m�kY�-
9./��X)V�pX�y\�N8�Z��/��N?�t�u�t�B]�vu,�ɧX���{ D�=(V��K��L=�a�U)9�H��)g�%r���9f4W�_LMK���	ZtSMC�`d�F�����H���i^�c�f��]���J��+�j���������AÚ:�
���b�GP�p�)H\�y?͢W_�����X�t%m5����wTڼ�;���[n�X��{��^�zQؐ�OA��6�R�@5�);WJ��53'1i�(eW�؇3��� �|O��j�8cF��L��L��E˰?w�cJ���*�W��p��}nji�4ʙԽsOet�y��&#�T�r�x�T�u<n��)a�m�Ϥ]Q3�g�r���N++�2�4��xE����裏��  ��td�\U�U�O�<#�^�7�\�[+�(�]��*��NS˞^����ڦ�Q{y>�UBkjy\��88�5!�5�5F
��b0Ω����iV���4ˬY�VK��3�9S����}X�H����  �����{)�d�l�+&d���S.P7(���B�;�^,��Η^e6��(���W+��zo��bUW˄�N��#���u\Ǻ���e�YST��h=��|p���w���ab֬Y4o�<  bA*�l/��x�[�j�����sRV ����[��})8�n��������U�����*a�4P��n�1mt1����c9��>_��9��x�2m�4 �0�%G�9)�2�I~��e=� �A�le6���.��2W�l��ʚRIӳ�W��CD���d*��(��)�j�  �6{P�DW�������H���I�2��!����j�}���*!�!�<u��sY�O��k�}�e   
bA*5S�*��e��m�OT;H�*s���؏��"-ߞQS��}iZ%����J�9��   @. ���#���B�tJ]�b�-%9ӎ�,#���G�9.�*WKL��   � ��C^{	�߆�Z��q��P�rgL�2��2QKr���.7^�^KƱ  �@�A��,�� l�u�ez����L���V��   �R � M6���]-Qhy�� �h���6h���1���^u�8�% bA�lʉ�� @Ahֿ~>VZ���;P%,���pg��*�{C�   ��G�J=�u_�A��CO�7Ѭ�۽�-�!�    �>Y�|���3=C�A��H(��y�4.�ce��"��G|  ~���������䌝o/Std�^+y>'�>�@��$Qs>� <��c?�R�%������[Roɽ�Z(�}a  ���������8�c1͜�N �:R��h|�A�:�z,Ӭ�$�9���!��%��V�!�����ܒ�k�\L׏z7�(
<��r�ku���2O���ya%M�j0���y��%��++	��FSF�є<d��\̮3l��|����{�d���}5Zo]�J�"��Pn�w	����v�Aa�#�g\��>���f��I�]1��5�;4�K��O.��?j�[.D]��]^�7Vѵ���Ӯ�O�]��<遥���+��GɴEǊtJ�R:��
��kGͯ��.+�j�}�� ����+o[L}z�i�_t���ѡӹ�R�|5��κz>�|�`���?�eB�.���u��x,����{�t���V��W߶���O�hՇ�R����'� a@SoRz�н�4��2���� �F��c�^^��:%�л	�� ?tv�;�����
\��',�w��8��E+]~�B���Y��XM~x�cٛ��u����'��0��OZ��Pg¹���[銔�_~Z�P�燞O?� �<�΅1�bIMt�Mj1�DRK��� ��ڤ��|��?�λ;��):b�'�xه�GNS9���4��!���z
��N�޲��~����Ko��H��}��+Eε�{ޯw��?�7�	������::�_��U����ǅ�<?��J�)�9�f� >���'������S5t�xyt2z��d%@��גʇ���K/���\9MUJ��u��53s����Cmi��Z�2I�|>����4��_����%�rJ޳�"<h@�qL/�u^x}M�kq�u8}�+3��Nӟ}c�U�wd�I�_+i��z:|��.7�!������5�>&"�<��N�G1cF3��/x!��A��;�`�T�s�} �� 2]7��S��{!����1���S׳����!���c�YP�/�S��o�&�Z�?܁��H!���T�����5Q��w�i��_��4ݿo��o��T�|5�]\�-m��o��ꕪ��Kmv��> �	K�c|M=%�:���3��dJ=9s�x���%��.4�k�+_�n}���.�^H|,�&��k�������;��+�Qc���8�<�/��O�~;�����F��]t�B�z��-��o���{��ެ�j��?��i��!L������S�T%�[��y�>��qg�zb4%�i�*p~�H_����.�G3�^~&�{]��e���;&�ՠ� �9��kGS���c�!�u��+Qz�fʽf��#���/�m�',���@u����������)����ҭ��-6��}��V:���N���#�9~0�?����v����+�,4���������Fgqq�',�+V�M̐]���u8oF3Ed>��$Ӣ��6���@��W�����o�	�R�q+Z�׶!�u�����!�1e�� �i��Q3��u]vڀ��T���
����G
ik7ƺ�|�`Zw����_�9f�4����ܯ�g���!�Ɛ��4={^'�x�ϴdY�R/������Ӕ�Ө5�}����\} �eZ����K�c��'4Jh	!>IM���H�1BNRF䕏��.��/�- Q���ӟ�����[I�a��)r_gF�딈=�Nf�U�?nmm-��!���M]M���)����Ó�p�x��Z�LI�:��=�y[�Nw�s����L,[����/��y>� 3oA'�t�ϴhi�R/��|�Y?Q��`���5�H==�-2SRBRg&�T�ńܧ$>��%ust�Խ9b��%��^>��+��:8�
�ؿ�o�C�cf��{���:GĞ�}wZXsK3%:���d�'����@O�HM����D��;ST�=���:g�����9�pI�R/ᖎ�U�� �0>�d��_7;��9��Ha`�O��덨��'�q��"=C�XUϰ���f�xe*9�,��1G�e�^�RrϹ��s��/~�����c��9�:���t���O:�  *�������DC������
!J&)���q�>��z�;��fB��t	���@]V���<�"o_��ѝbV����9��:���8���kE3�    U㞻/��!1i��jO�x���SG�$�'�	�xC�����t�W�"��]p���s��(��_s�˖/��{OQ��   @�x�����Hn��������4:��t��BO���@G�M�)դd����Yh����Ya�6
?�V�	�__T�Yb   ��r¸c豧������	�љVw���G&�R�x)�c#� !/��q�Vso#�l����(�c���z�!z�>l�=    �ʊ����1�ӝw�Mn���5͕Oo�:x�([gG�1���uMe�t�G�y]]��w�#���D'M�8��|gIb   ���rȁ�>��w,:�(���R㾦�ez�4-c-����蠏>�����*�a�̒#�    �᱇��ÆѦ�oA��.]�rH��PL��\c+V,���Υi~Hm��yb   �����7 � � � �F��M7ݔ�zꩂG}�i��(�HЛo�I    �} � T��ݻ��g�M={�̺���7�Ls��ɺ�u�]G믿>m���t�W�}<��?]u�Ub\�wܑ/�g�=묳h�6�{��<�=��   �� ���t�ڕ&N�H[m������b:�c��̸N}}��;v,}��"r�=z��<q���j�#Rl��֔/\>΋    �b@a��<y2m��f��2d�{�t��Gg�{ɹ�K������j�+��R�!r   T�= e���IH=��3��H�ɖ��{�<x��{��Ϛ5+��\|��t�)�P�9�s�~ȹ��_v�e"�/����#    T�= e�e{ʔ)��&���|�	�t�I�z���}��W���_9f�����iܸq4cƌ��q���{�I��׿��|��w��7��\��{ɒ%t뭷�4!��g����	    �b@`1�Rϑ�O<����}m��/�O?�D��r��ߟn��v�u�]snw��{�'����[�����n��F�g��J
W    P~ � ��>}�X�y��R/��A$$��/�̸^gg'���޽{���/Fߩ���:���۴��;���    T�= e��q��͛G�rH�uX������_.:��t�j�aw   �*@��a����O��ѣ���.��R�6m-_��     � � N���oKÇ��t��.��     � ����V��뮻D*̘1c��_�:    �{ B�����O�gX�����Cl    @��^{-m��v4h� :t(�q�4~�x   @���P%v�m7�x�s����F�&M�ϕ+W��5��cǎ��_~���}   @���Pxv�	&P<Ϲ.���{�7ޠ�^z�v�}w�o����ۏZZZ    �b@�������>e�?G��j+1Qְa��SN	    ��= U����L�X��{ٲe"���k�����?���xF[    ��= !��y�;Ｓ��������墳��    > � �ί��/I={���#G�	'�@��z+    |@�1,��n�I�i�{���k�    ������c�ў{�I��կ���������    �b@��u�.��Bz�g�k׮Էo_�i��    �b@��a����k����Z�u_*�ΝK'N���>��I�~�h���   ����̰L��P�>����9e�%�G�)%���%g��6�r�c��}��4d�   @��P�O�N[n��x̳�r��u�]W����=��ҥ�;��<�LG������W�cJ&�t���O<Q�� �[x�K�����	    �b@�ꪫh���t�'R<�=�P1����U�VQ"��^�z��MMM�c���?O�]vYɎ�S�&O�,f��äI����3�:\!8p�cٌ3�3΀��'�y��i�Ɲݹ�[�n�5�����M<���<�^��  @��pt���n��?�X��*ŗg�>|x��9u�ꫯ�'�|���v�]w�.���+~���y����  p²>b�1��gL޸b��ؘ��88�b�
0��4��͛G��=͜9ST   �b@y���i̘1"z����L��l�N�J�_=�������O����y�<{�I'	���Y�t)��Y�fф	0N> 
�9�h���m�6�5�X���p�"��[���z륽>�|�R����W_}E�~���� �	��2�l�2��KĭTp�<紳�O\�iA�����1�C ����_��V[���<�l54h��m��v�9޿�����č+� �� ��F)T�%��P8��7����bԩR�hUJ8��+|�;N�y�7���_}c  ��   �N��(�{�!$Yv�/�A���p'�R�O{�!����ٳ��_��^z��,YB ��b   ���Z��o?���~G�{�.x?ܩ�����q��+w�厰<��2��q� ��pK�s~��;t�PZs�5�q�w�=���裏���{��~�i�6m j�=   ����_�<�@��o�wԼ������k���/�o���p��B��=���[&�w�Nk����P�w7�xc0`�����=<c��5�'��T�\C� ��   � �d��_�򗾷a���g�s*��ŏyX�J��;\���6���ܩ�o[l��5>~6�Yg:���E��|P��@�.{   �ŨQ���o���g���f�#*C[�adK	�<��s��}�o w��~��E�?\)�a{9����W^yE� , �   �	竳��瞾F����^xAt8]�h�
<*���%��~����7�<k�����Kp M�8QTf  �b   ����Gyd��5O$�i6O<��\Z�k�|ni��;O�ǒ�������7�,��Y�k�R@���  �4�G~�Yg���`~�������N<���w�I<��h������3�ϩ<<o�-\� T�=  �H£�q�"o�g�;�r��n1��������C^r���C�~��y�ˑ}ο�e�]�k����� �  9�N\p�=:�z�vʔ)b��(­O=����s�����8�Ϻ{�]w��W_}�  �b   R���t�i�Qccc�uf̘A�&M��>�� �ɲz�!�r1n�8�7��d��{�0�7�t����ٺk׮���-;|�1jp��  �,$'������l�+Y�Hb;�B !d���W(�@��J��e�_ii�
eZZhٳl(6!���'�����s�+_]]IW�����Oؾ�eY������\t����O<�6e�c���*����>�%��N��;�#Ԛ�[n�E�K�;6LF��.8���� ���m8���ذ�2.�6m��7]8�K{""�x�?��jép���{��_���Rd˖-S�$����j��>(w�q�|��B�����ԩS�[���aЌKQQ��]���,X�~��6����u�DD��v�yg�ӟ��B��6>��㜥��7���ꫯ�7�����5Ci�m�ݦ6�z��'���Sؘ젃Ra�M=\�=�X�=	�����[�裏�~�{""�X�����~v�'�Dn��vY�f�P׬X�B.��B���T�L3��!g�u����Omj��S�d�������'a����.'�t�꤄���[o��͛�������2꼱K�UM0|��'r�]w��7P_�2��K����999!�����Zfb ��~�Y(�A����1cl~6�y��}�v�3��/X4�~�0hƙ��cA:�=��<��Ng���0�8����SO�E��6��}��]�`ODD�c�����ʲs��#�<�������0{;q�D��c��/��Bͼw�;�#�W�V��f�<�@U���(X�L�p��N9���$,�F�;:@��3����ڈ�c�ŨQ�T?.h�ZXXhy[���z\P��NL~��x<!{쉈(�`f���/W!�3��19q]m���3�O?��� �w�ʕ+UY���G;vl��(��FV7�t����
�f�O8��� ʞ"���9s�����{�kZab���+����X\���{�M��uV�`��o���>[�w�}�gzl`�'"�����p�3�X����X�� �fRsssUY��=o��p���=`V�EY��F@l��Qn�p�M���l9�Z�� J'����c�=&���TWWw�{����_���r��7ˌ3B���-X�yϰ�}x�Q���i0�����O�g�;�˳�>���̙3�����!�<x�:�v��'�.K���
�����2�K&�B=��z�v����Ԍu"����
��zv���@c���j�W�c��կT�{�W�ە�pv%7x�Q�m��,�e;��k����
5P
�g^x�Un���g8c��8&1@����L���������<R({""J{(���UM=f'���:�%�A5����賡�}�����FB� ���ѣG>g�ѵ��0V��ŢZ��w�q!������|�p�CW�g��l���s��fė/_.� �3�~�����{$��!�C�δi��٧�^{�lM쉈(���f~�:o ��4~�g�z�v�HP�����ΆZ�E��\rI �����S���?�|��R!@�B�����w�E(�E�^(��F��0�=�Ͻ=�4�}�?�,�~��G�z��o��F]�������]�3L�^z���~j�
nvՉ������~��U�z��c�>���]AVl���P��hݺ�:u�*��:��E9���]QRR����ֵk�Z����7�Pl�<���u�>0��a��2�X�)`=챎�裏���3�T�X��}���U��4�������Z2Z_b�^�xݙc.JxP��3Q�`ODDi
GQ*b��e��暄����f��8��1fQ��C��;U�Q�2&��	&�{ｧ�%� b�p�=��Pz�!�]�Ǉ�׆��9��3�'�xb�u���j����ٳg�����^K����J��N��4������f�ƍr�"���o����w�!��Z�z�駫Ё^�f,�m��T���)��/��6�BhB�!Ύ`�"B>:��R�Ѕ���)S�]�����E]�7zo��ڃ�E�٪U�Ծ ��r�(����^��n���t��(���ћ�H`�'"���.+ư�Cp���[�~�dC/xԖc�������^$�u�V�Xpfe�u5�v�E�瞫7��Q��a��
�5��̒�<B:�!������녋";vdEY��y�-�kQO��p�8%�0[\}���.qi�;���v�d9��r�#�!>�W|�>񹵋�'�&�x��S����]׮����ŋ���SevtP�uX�}�}�����)_Kg�DD�VrP�mm�Ri�~X������#�[o���ǀ��YN}-�8J7����Q
�7�y���L*s��=�Q�ol�	S�NU���Eco�V�L�K͚��T��S񂐞]�+9��$�,O���h�|^���)SvIp�&b�5�Ҷ�Eڶ�H{Uk\�>֣`p��$�(�,O��x؃�[UTTHo�`ODDi�81�E�f�����JP�� ��H�Ah[8x�>r�����|�}������Y�&�m��MR�qc`�m$��׃}ii��p�G,�Ca �r�Y������_�B?v��GP��3,�6�8K���T8�����A�3��������#y#$wH�������w���.�Q���}U�o��,-U��y��E0h�N�X��1}c7��g�p�g��;қ0�Q�@����Gk?��T����o��ٰ#dҔ)2q�d�e���z����TWU���_�x�,��{Y�lYH`�&E|���X���s�e��\�����<�L`a.j�q������,2�̿����Wo���}���k����Iw[;f��`׾�;��8s:�6����?�G�}8�S�z��rHް|u�4��e�6P]]/�֮�]�4���5��%��bm��%k}20�QZ@9˩��r!��v�&�=��Î<R��1CJ-��tf�q�4u���T�����#-h��g�N)��Į�z�t��Y����CKE�qt�A:t�u�Q��h0P@��I�&�|0�CyUo1l�0�Z6�zl��윝	'�([
w������
�� ��A�5;���v����h���I��~Ҵ�A�Vԩ��X�~�
���M�PƄ5
(��-���R��b�1������D�XoI�%8�V3�h#�z�jIU%��r��Ǫ@?D�=d��w_uA`G�O�K-R�Sa7R���?���[�N4��ۇ�p��/�Ÿ��{�1@��ͥ'�!���>R�_2B(�0ۋ�G`��Xʦ���]R�g���B���7���u�/�dW��^:����!?h6o��b�΅�gT�4�m��e��m�}į��ju��xVkr0XB;�Llj�`O�"�YNu갼|sh�#E������
ˍ�(��>|�ر!��ϟ��lS�@����SN����@=z�a���3�eْ%���ϫ�,.�7Ϛ<y���GA,X���	q���X�+t�y��U��#$��%;�b����0xB(���	N��](����C��Rj�Ο5�'�|�Fz98�7p�1��j��#�B���c���9���ߥH��(���5Ҵ�swd��(��nP�o��=����{��曻�\�{�����C��-[�c�P��]�ѢԆh􍞌Pr�� �VW߿�Xξ�5Cߕ���2~��E��V��?�y��x����[������983b�f�uؔ�;�	��.��O�q�pf!�݄���9ǂO#�c@痮Qt��;�D\E�3���y��}_g����p�a��wS������E�>�
���n�8�hJ��ȗ�o�b.�ihhP�������j�:1e����zĐ!C�L@���L߸$/7W,ӂ�v�{��:z��3��16�h :�${*#��z�rᥗJQ7f�{ڮ��.o�����{o�wBw���ҏ���?j�3RG�ģ-%���g���{,��}�?��c�2�i�����a18��t�te-���xP�>Co�x��Yo�����r�&����Yz��;�{��3x&?�}�|�#�r�I�ქ��*i���sPYY�ں"�K�0p]�h�|�����3ܯ�k�M\��`��L�r�e�rG�Px���C���n���n�X�i���W_}URŨ�w�kn�Q�X���Q�G˚-[d�֭2հ,ʆp�%6�x���R���p~��>�z��SO=%[���.L��P�o���ź��6�`�^��4B�8f�c�`ɑ�T��yC�g����?�{��x��s��ƙ���o��olN���Tpi�\wܗ�_����ǣ6��z:2��}�~�L~�B^}����{�� �.k���U�څA?��0@�_��Z������N9�D)���@�YUU͙{z�O�N(�=��5�8�aO��kԯ_z�U���S��Y|��we�q�dԨQ��Pߎ�\ ��(�[\�P2�I�x�@y�w[�`�)b�X+��l:������s�����%���v���7�x�Ǧ@�z��C}V�K��lq�qZaF����i� ���$�Y�mn�Mn��s�3�S����q�_��{C�=�,Dv����B|m��/_�v8ƢZւ��&>3�|���(���,g�x��z����6~�xUk�Yd�NO6�˯�F���~��8��	A�����B�S@��lUo��1x�Y�r����kr�	'|���PW��>/��13�M��0�M�0�	0+o^,��㏫�@����T���Y������z ��PC&��9����唸т�3ץ.�7WrOs�x����v����:�s˙{������Ϸ��vamւa�=�bZl����[2�}/�3��Hu���l5Q�d.Q �^�EL6����;dwm���mmRW[�zl#�����w�3�}������Y�E�k�Сҿ�D.��r)����Ps_�3C��fb�mOl ���0x3.΅��>Z����/��1c��!��{�E΀\�7�L�C������{�}vq��s%�(֕���wC�x��T�NǕ�Y|�l���7��� ���Z��O��p�}���>�{b�T�m^S�}/��fx��<�iӦ	�.�}s�ԩ!��}�ݸ�rw�X�v�]2b��.}>&Wj���B���d�;&3|>C}�>6�{�@�Z�/\ gJ�ʤL���ځ������ܣ-��+6�B�u@���eɒ%=>I��1p0�Y
�x@�ʟ���{�E,�ivq���^�%9	�����Yv��<Jo���٥}�U��@g��rD
��]�.��V�[��4'B��wI񁃤ꓭ�m����8�{�m��C=��Ǡ?�SM��Z��`ODD)'���%N�aZ����{��k,�֭�U�k{�BD���5V���p�6`ئ}��~��N��1vF�c���kU z��7T�2.��x�b5�m�a���ƺ�4U`a��kFb�5��&��g齡���d�H���8������kZ���@��h�O��(՟V���^�_�f�ڧ��3��XC��N������R
B�r����Kj	���+�P���i�F�R^2#��z�i�F��=����U�q�E�u�L?�up{<��g�?�`?r�(���m�����+���E>О�dy��'C�=f��;�8y�g$�`A0v�5���F�r�i�v�A��u��z��|��F����Ajal���Y8��ijO]�:�`'ܻ�fK�����Β�(01p�a�-��կ~%s��͘V��DD�RN8ᄐ�k�_~Y����y�4lxcJn֮^�gA���;4�W̎cA���^��'�Z#��Xt(���W����}o��I~X�T�ጃ�uK���^�f����kI�ڣ�;!أ]-0N#���`�37�,�L{���.8�]�ۍ���x��@��Bվ2�aЁ:|Ou�z�v½�W�<{���|���w�8�>�h���#�H&`��^��{���Vl���G$/7/hC��̲��s#Q�C�9sf�q�Q߰a�$B�� ��.���D6�[��n�\n��q�Y�os��$[{��{\ol`�\3c=��_;�?Hhӂ�[� �TUV������#���=�M��"�_y��^�J���_�[��`�z����O-�M�hϻy�JC���(أ�
����ު�+�����`�U������0�ʜ.�_�G�5-�=���Za�(���i^�h�k|�R�A�qS��?^mʖ	`2�S��Y8,2�c[�6[=o���}�R_I���Ƕ��!�_{�5I��/�@��sO۷���+���s�L}a,B{���FoY�0������i8c�0܇Q ��i�����}��*ط��u|���+e���K��,���]$����S<}��g��\��^���Ѫ��3Ă��{�����#c�v���,c��՜2��W)éz���ݣ��RY�_vf5��;�D�k��x����XD�A�~f�q쓀үt�`ODD)a�����{I�}�?�'�j�#i��Wu��$�����9�𞓛��W��1{��h��>�a�_�{��G�{�_�o���s���ذ�5�(ͱc�a�,�?�AtCB�q#��c�;��:,b>蠃�����K��h��N�wi�����E��	.�q�ϕ��ػ"����*��XT��Q�0��k1�1��`0�o�R5gk�s:k�ե�� J �31���=��h�.fo��vR��(+�kn��vM:��W._�@ָ0V�X��5�X0�@��aW��׍�x�xfm1��������~�@��h_]e�����#m}�r�,�?_���%������n2�]���!�cJ����������cx��,G�3��ު�^�ԧs�7� %�1�����%9XL�gL�4���-	gK�i��s���X���t�`ODD)!�j���ٳ��x~u�j#*;P�n���z�УG�
��[������f�1���|���c��-�?���?m���6�k�ڵ���Ѷ���.�H���+�L�,����U�����;�������|����+��b��)�4WՑ���HP��;�]�Y~Zb�,G��pJ`wZ���q��uS�xl��ǚ�y|���cؔ���(ۈ����R�Й-\�Pmޓh{�L�h�i�7˗-
�z8׃�
�}�j���=p�^��ݳ�E��:�������0�P��B����rUnM~A��{�r���$�6gΜ�`���P{��;��uml_�͒^}�U[��.8�W,Jp�3��mnY�wNY���+�U-�޾c`�쒃�?EK�f�v[w���(��gJKKUC�o��F��=%�p��c�������M;���������O�����g��{�-B��s���X]���֫��ה��e8C���3�3����C�<R��]U��H�d���v�����nPNs���>����Zy#�U��9[/�%8��ˢO}ajl<��R�����\�c�;��:��^}�?�(˴A��ߞ#��7�=Q7`&�X�˟~�i��q'�hkQ)�1:̘w����f�f�1S�矵Wa�����e6]h��ru|=U��FЅ�*�oW3�vZa�{�Er��'t�ʆ������o���v�Iƌt�ni~n�c��g��=�ko�K��37K2�?_��nu�}������}��+{���y����:�%�T<0�QҡÉ�����W��??�$[��n���6|�(���7vz���{�Pֿ�����ܣ�nз��"P�zN��VN�@cw��Z��ƌ+{k?�ys�J"a�Ps�ǂk<�v;�$�O~򓠏Q2�M����/�������Y�a�,~���k�_�����y:��@��i�>�]�#��mQ�g/���� ��"ܣS:b�'"��B�4�NC2N��<�h[��Q������j����F@�,�Koe�
����ew�}�Ytc��3f��� �--���B�Rͬ3�Hx��zM�y�4iRʕO�96���ݳ�uV����ݠ������I3^�Nm��mh���ֵ���k_��&�"oα�q-��0�u��#,7��7o^B��ɳfٺ��ի�,�,��s�����P�{c���ii�����xx�x<�`� s$��/'O�EH�lݺUu39rd��=��3���;��������>�ˢ}��l��(����3�wE9|��fwǂ���ڣ|�����|��zJճ@���W��	&�C}�+�8�<8��P�^�_���z�}�
��֖z��+J<�l�YGz����Я�ڱC�ku�1	��NI�`o�J��S�}�q�Fٴi����3����j��短�&d��7���OC[���VXH�7<_�V�G��o��6ha6�"��x�a�'"���
e?Xt��i�yd�� L���U�z��ꍡ;�5�:��^=~<>�c��]i����:�H�?� y�����5��{lбq�Ʃ�ܸ�9�Pd��� H�a��N8���?[���gNf/�Ǒ�%�fG�	��]��{���ߜ�'�M�2�����(V�En�t�҄>t��ӷ���J�!��B���^�z�s盠�C%�,'��8v���k�m7Qo�҂=��d���=������#��d��ǁҗ�+WJ*������{[��38O9�]f��g�����z�%9���8��hhQ�䮋>�����v�N�DD�4�Ç9�ٳD������6,���+��Y�aUO��2cliid�z�\��x�
���O��Z�C?<��u�555!�2R)؏;V
��E	�����������oy�����j��T�|�;b9�ʳ��:��ǻ��644H:�ݯ
""J*��v�B��Y�&��c�EW3��KN�P��_ �����<n�>j����=a���&������8Q���DY�v�*�0=z��
��_�^���m}n�@�L���o�
{G{ˈ�z�v��cql�ߣ��<iZ��	(����F���	��������f(ٱ#z��x�h
�V�o�ho	���߳>P��>����2;�6��V��>��8���������t��=~��D�C��~�]v�T1´��d�u�t���;S�%9ǰ-u��{�<�'\�}΀\�nA�� �30�`����`O�FP�[YYi�؍��݊�
Y�pQ̏���E�z�aÆ��ll"��x��]_��[a�X
�Ne�;��3�N��7�w�M��1ܛ7�
G��˿;m��c�f��c�g�ɓ�׭[r�굔,�=h�i���7�Oc���.�8\�sѬ�3[�_�u���r�ϖ���g��s2�t�`O�Z��m?��
�
-k��2ِ!CB����a�i���[Ԝ��o�Z4믭w���e8� ��;�:��W����5z������͛C���������d3B����=����J��Yy�n�]�����楞]�k+؛N�Z:ૃ���f�E��m۶%�1�5*�m�kk��}�]�2��	ǿ�4�>E�},�u�u����Q;�$���fx��l�"Ʉ=�Sٝ@�*�e�u��Yy,�1B���y*��K�`���m�DD�49��`6�Ƭ\�C*�Km��e8jWY\aQl��8���c0`l����%E���0oެ�㉾sgQ߾ҷ_?�3�z�;7��P��=f��;�?�3V�lPt��N���#��NV���k���)�v�e�'"��)..9�腳�m{�����S���ްH6����};�>��6�~|�nC�N$X��,A�����Jt��6�H6�k�g;g9���OVh�=�&�� Kj��D\@ku&Ċy ���}Ity`w0�QR`A�y�У<Q���,������b��i�ݎT~c숓������|��U���g�u��`?t�pYf�yTO�Y�T�}��	���0(��V�D{G��:ўt��kiPzfl�۷o_{""�h���,��^z�+9f\-��E-.�I��{��b<���z���(�j-�$�1X1{�Nő����n��6����tF��3m�_��_G�0X��=%E�`__}3�x�3�0+z�5֢�f��;���Mm��HV@�n��RPP���{;%6�u&xZ:W[��;���cc5Č��Ύԩ����:���e��1q��9}&�����}��ײ�bW�:c�=�q���BCf���K魬�p ��#�K��0j5��s�x��'C��og��`�j��hm9���8N�����}i�(���Eny�P�o���gX���Je��ԩSd��]�~�۷�`��3a��}���v��/���m�Aa�p����}�D� �;ci����AZz0���u6�}~�g�����d�r)g����b��	��T,�"��DD�+Y��D�փ���$�ȑ�>*�_,�e<X�VR!�����}Ecc�D�a��5��I�뺻쉈()��&������p�݃>U���얜ċU�[*��σ�3>w�׾���1�[��D|~�k$=��]�DD�Ve7��gm�f���2S�����f�]�e�<X�����n#�{3�u�e6�:[ϯ��R��k*�DD��P#m'���B����0������Ot��z�X-�M4s��cc�<�etQ�黩v>�>��M��YO��]�p¿R��؛ϰ$�KW<0�QR����H���	��h�ٹyy�b
lƚ{��La���6�ıl"��}WKq�m��y�n9���~]�z����Ot,����k>Ò�}5������"\};j\5K�D��M����o�g�!��8��lڰA�\�����������M@�;��{$��{^���6��O{N;ą�ip������?��'""��j�P@J�S�h�!���:�
z���{�(E��;/H���%����r,�k*�***�>����Y?O���W�i����?ԛ�$��G���L<�W;��1�*n߾]�	_������0��Woٔ�Y"JM:���nGڞ�i�ƨ�)��Di�A�8�c�ۦ�,�vh᧵�Uɸ;�.�&�l٢�q!����e���Q?�S���UՌ4ڪ��۪��$��g��MP��a~����:ی�I�6Xe�K�U�˵_�����ܱM�����Њ���8���c�����_@BN�Jp|"Qgo,/;���<��f�:I��	u�b�f5jT���`�npK.�	���x�Oڣ�����F�L�vf��7���{""J�;v��!C�$�1,Z���́�naQ���g��E�^��h�a6߸`VT���N�_���ݙ�gu�j��e0ɂ]�����i��<�h�:�v���Lm��V��P�b1���h��w6�������n�*�M��J�c@X_�n]�:�ee�`��lt`iokS�����d�8{o,��[gZ��t7�w�~̏�?�{r�[}F�(��~������zJ�@h����h�8��Y_��j|�nq�2�I{�2O�[-��c�ȑA3�� ��f�������G��Ⱥ5k�쾺h����z��jA8++˲$�%���8c��v��F�d�A}��#M��3=&L��x�����Ź%9�8�}�ξ�]��� 'z�O����Cs�߰!���UADDIc5�jwv3����+��I'E�;�}�*�������B;;�8\�OF�7�N�������.��^#V��dY�pa��%%%*4�_�>��mo�������G-��x�Ӭ���wL��V���������M�<9��SW�Z%������f͚5!ǆ�v���',^�@�WTH���o7d�0��J{-��ǥ��v�}�tŪf?Ҍm�����
�����z�	d����gϖDmqve]��D�m�65h5�M�2�V�o-o�����?z�v�6�#qc�^{����j(�	�+��ߺ�޿#�F�-J��bՋ_DD�lV�ar��v�~�!a�A��?��g͊x;�"�9�i�:t��6- ���Ņ���V���\c�P��?kuv*ԣ��_f�g�8�g/0(J4�`o�ZJ�����O��������z��k�nU]\��������@��.N�xZ{o��u��G�)���-�k�w6	/�Ix]�C/}EQ*��B���RZZt|�]wMh��<G�0b�(���Q�#�?G��K��c�SG�Z{0����U�?�����؝�����	/���ʼ��Z�G04{<�v����R�G��r���`/����.�>ѻeo���k�_����7���s}��	^/�DD�T�c5{,6|��7�86�['�ϗ�S�F��,<X�mݪ�q;f�`ߞ�+Y�BZgd�p!>��>\���h��Oaa��D����3�q�ƅ:��LB/�H���3�1�M��&)߿3�:o��8(�o��^��&��E����`��m����<0�w�W�^-������j�ҥ2mڴ�c�����F�0|�H���T�݃��.�����ŦXH+�Zw�����̽��ܦ�;A���"ݗ�u�@�Jp���=[�-	�%��sϐchK��?�g�V�X!��[�ؑGi+أEc��&��o1k����w{���.Y�'����;g�#��4��W5�v��b4w�ܴ�qV�`ODDI�dɒ�cXt8`� ��U"a�~��x�GX ��3FV._��ꊓ�%������A���{c�7�z���z��	Ww�:�x:f?q���ΆT��_z�yI�`o�J�k�c�?������0�ay]G��f�;��w}�8�\���-r<>�AW�D}��v����B�]�q�hv���=%�r-����Zq���w�}7��g��[�3���Jr0�ݦ�{��6]����[�Y��t�	'���ǿX��o�Yh�>�3Gʓ�yO^^��ٜŋK*�����/����������~���MZ�5K�>�����:Kr�c������G2���M��T��k�ks��̙3�>�dB�.�{""J���VU�3iҤ����_R���_-_���7cF��b!mSc���׫0ݦ�z�}�;�#���>\Y�~]O2���m-�P�E�vJp���䱇�d�:u���Tb(��od��t�QG�
���C]G�cI���������OS�d�gnIJp|��%8��o\Ug�>�z7���g��e8�`ODDI�����~���R%,z�H"��d�"1�	���q�T�NkK����CA�d�/��Vj�%:=��V���6@�h���ٌ
�}�I��2��g��c�_���
�8�`��	�u����^�*-%oDg���&fN�-�grv��{P���$��$Ӡ����W�utͱ�ft?�t�`ODDI7o�<������,�����ۄ?�
-(���srƹ�F�-��nZ��a�R�z����:��Ӽ�6]q�^�hk����'?_����A�7_}U��"���aP�ʾ��K������������/)��v��ϯ_\#9���Ю����m���P�||�iWI�8���yI��gS�FQ�Jp<ni\io�^�9���ڵk%�1�Q�a����ٳC9$)��8t�i�d����6G����C�k� �*��P�|}���͝q����!3�������\[����㎤�ƉE�XPm�&����/�,�~��>����O4�}n��V�&w���-�rv}Ύf9��n�l-�c���}?���.8G�P�����1}�t3fLб��|�c�'"��C���O�SN	:�S���_;ZH&읷�*>����������U˗��{ii�(��ܫ۠LG�G�b[s��x����>��,=~~A�������W��d9��B�UUU���Y�7�xCN=�T)**R�g>k�,�뮻l}>��Q �b���8s/3��CgG�o��b����>|��֖Q�lhT���eڌ%]_}���;{���c�����,,�̶���KN��?�D��*�#����_$�1�$�;�[��G[a��k�~�M���\��-��3!3�Z���v�]s�B���S�L����b�b����s�g���K�`��Ar��?N����������q��cGq�<��3�y�樟��[��)=l�8r�ڦ�{Gg�=���,����O;���k�z;%8u���	�����=�쳒΋fu�ԫa6;�,]��wDS\\,�w�c��_�ڵ�D=	m/�nݪz���g?KZ��o��J���ee� `1B

eݚ5�l��?+��o�҂*�*µ��=���#o����o�t}�.��f��u�5��R,����W��w�-Ʉ����r��t��+��I'��*�W^y��p��>�V�~W)���uWs��M�T�H�}:��cӭ����-ԋ��k���;p�%���
��L�`ODD)a���ޓ��:+�8:���>��O�~�1����N��9�s?a�$��]d���{�l���(�Qi�V��q���`�N9��y�s}����ӻ
�^$�C���j�-=��c�	9�0��SY���S%9��vZ�^�p�|����uK�j�X���4�b�^��pL���fq�M�R��E�jۡ^S��Z���gG�t��'�LJ�����?e""�5�y�U�`,{������G%���ߤ��D8�`۟��>j�e����<���I�{�[�v=�=f��~`��-��q�^zC_z=�#ܣ���/+���%��ħ��V~{��RUY)Ʉ6y���o��V����7�C=4h��e�]&�}����h�aI�d�$ϼ+���Kuc�!��:Za�ڼZ��G
V��m�[|nKK�AFy���k�y]�����	�C��
�{
k��&K��1"���f"D�\��%6�2:��T�
��'`���?�I�����b�|��vS��[7o���UڇP���`6#Ԩ�w�BZ}�9��a^���Ko0�Y��.z@�G�ߔ��e�N>�����t�7���?��O��[�j�>fy�{w�����U���9�,���s�g�}mnqWy�U���Rh����阥��l���6,���kaeܛ����?�����O�RNAQ���'�VPX$DD�\�챈;v�������&�B�%W^)?��B��e�]Ռ}uU��TW��
f�s��=B���7�ԋ�9z���P�0����.��mݲEn��:��7ٰfɼ3(|��gR��3	]�u�o|�c���,v;�`1m��;������o�Y��zi�a�^���u-Lg!໒W{�k����c1w,��к�I��W����>��}^}�U[��{""J)=�ׯ�Q�FGm,�/��G]��������i��ޥq�ݔ�.�5�~KS��i����gg�	�(�Qe<Z���|n^��c#Y�|��r��{K�V-9_z�%Ig�����k������7߬6i���{۽R�Y���^&9L��,f��=[�GX�ZӪ:�8�h?;q�\}��������,=��7IͼJ���a��v�+��"�Z�>��S�i쉈(�`��\s�5A��-�'?��
�Ɇǈ��V���n�!П�+������ż(�=�{b��9�/�s���_����8��"�-R;�����r�A�q�岲2�馛��ni�
��o����\c�=�g��9��ٞ�֎uyNq�z��=zҷy��ڹ�#��5����R��:��U(����~����}�ݧJ�2�=��O�}��RZZt���OW�s��a���_|!�_p�ܨ;;��.��D��N�h���9s$����P{����?��L��c	2cƌ�1�W�FV/����;�rr�J)l�H�h��U�׻Ψ|Am�x��;jr��{�訷���:��襏Ű�v��ZQv!�#�c�pӪ��
Z�b���l�ۓ쉈(�`�7,����˃�c������0�
lbuï-'kA�풓�>��͛;W��_U[�T��%�9�a����c��w�}���_����w�y�a����/�ߗ�'�����M�N.т�Eb6|�y��������y���_���腯8�����:ڬ�<�����y�c�����.;���Eb�}�6�g{���K�b�'"�����^"��y�jF?U��g�{�I�3{�\|���i���W�	-P~�=�Tt�EY����`�����.��sO`'`�E��u�]g{1��b��m�o���m}#=T��g�}˳յ(���{�G�o���&4��ka^׶�E�����c�����/�8�ֲ�v�m)sƯ'0�QJ��g�yF������(�s�Qm�R:�����T���@v7NR	��k/�$o��r��қ��r��^�7�V��k0`9����0�A ���-�֭������R��V)�O���#\ͼ����s[���0�d:�� ���^i��V��K�q{ｷ\��A�a`@��?�Y�n��쉈(eaêO<1�FV�+VH*�f�\u�C�'͚%�M����SSS#o�������^0��>�^b^K�P���C2���?���u��۷�
�x>b�u�0�I��M(�	�w��i��^ߝ0�������Ե�W�ﾻ��P{B����u�F��_�������-�����ZA�5�_��㘉C�N�'��e$K/V��������#�>Zv�I8�1��o��?�ϴ�-�:�4�e�]B�Ϟ=;�;�D���@����l:���7ܠ��c�ipK���7�@
v�+���b[�w�m�lUN����&M���t`�e#,FN�u9=����Z�q��%�����BBc�=z�����g%�mX�N��.�?��L�{oU�3i��㩮�V-X ���|��'R_W'�b���j��YSS�<�裒�?��'�N�8���<����7���K�v�[66J˦F��G
v�+�Ź�*�W֩�����X�`^����ʽ�=��|P&O���AZ��㏒޾��u���G�#ô`;|�H2t��ͦ� v�j�X/\(�׮U_#�`��7�h�`��������,���{�c�x�e9蠃��vb��(s��9y#$oX�8�<5�����MҼ�Aګ�&��c�Um-�5��Jw�uWF-�������Rj�����K/:�:�����S%9�PjbV]U%����r�� �r,�f��1�Ʒ47K�v��|�.~�
��[����_]ztn��l��e�=��FK蠃A����n}���-2s���>#
${@n��|��۷�H�Fi�֢Ztv~W����N���?�;�#�K�z�=���^{M;�0g�4����\rIJv��
�+���V��`�ĉ��_�2�8f���"�@tW]]�\{�r�-��4C�T�ɹꪫT���c�>�W����s�Kr$�,O�|W�q�8��<�nq׶������i���yqq�*O2�-�0�ڜ���a��^#������mq��ή����+=rs�rCv�$�N���,�#�<R�s�qǩ�]�JK����o)� ��Y�v��V8#��A��c�	�����w�Yn��ָ��a�M��9Y�U�%��lq�f�#ǩf��δ.�jKٱìW��[o�G<���nhW�{ʔ)ST�/))	�e�oDo�`O���L��م�B!��6oެ�֡T�h͚5�j�*�ԇ2
�Hw]ա���/�(����{�jW��_�"hr	��1+�]Tq6gz����<��mSʑ�>�l9��C&�0���vh�ۛ1�QZy��e�}���:(�8Ϊaq!�rRiWZ�v�嗫23����Lo,����tZ�l�j{���:���z?ꨣT��jלt��7x��h�588{��-Q�b�'"���N�F�R�!C��s��o͠ť���Q>e��|ܾ}�P0��^p��<����Zb��#�ha�?S�w�޸�����?W����쉈(��9v������v��馛�g}S6`���-�{��'��α���ꫯV�`082�M@iʑG)�����+�<���k�	�sa�
��k�]�0�y�7�:1�QZZ�n�����oRo�2�ڣ>�7��Nu����V�e�	Y:l6�l����P4@�vs�(��s�9�$�͟�y����t�R�Ї����߫3�ׯ
�`ODDi���=�ܐ��I�z��Mɇ>�8˂�̰��u��Y�r�*Q�����|AAA��8�u�'�O�S��}�ݔ]X���[�z�ja���x衇�O>��`ODDi�g�����P`v�	'�n?�0g�5᨝7�M>boQl0z��W� ��a���t���.8�5{�lU��
���9R�q���bu�FiJ��:�������:k�?m  �IDAT�����;�"#P����p��^r�m���i��EX�N�"����J��{�9��*�6s�����?_��?�*kY�|y���4Cḯ	ԦR(�;vl��c�[o��Z�rA�=�DD���m<Z]"�X�Dy�Ǫp����l G]���HȪ����Q�o�,2��K�<��2k�,�9s��s��?y�du̂#�/\�Pm
�q�Fٺuk����C��#F��ѣզR(ǲz<fX�E�/��RFu�I{""����BZ���c�=B���~��c ���B�Δ`v�j渥�E�ߠN����s�=���O��G�^�Æ{{z�M����*�#\c ���A .����H�����RXX�6C�Gy\�Z�p�����W;H�}e�0�Q�@��,0bN�4)�z�棛f��l�".�K.��R9���-�G D�_�x�PϪ��Pu鸠�3��~����/��bf�;��$����*̯����`ODD��7�x�������\���v�w�y�|��B����&V�P�YX�l�Ch���.XH������[Y�U�)(�������_�d	׾��=e,�C�D�D�<3�D�ꩧTW��C�<�(Ű��7X(˚��B�6�7C�{��B��y��n�������B'*�5@I,P��(Ţ��`ODD	���o�6�Yg�r=f)�>�l5�����tꨱ��@��5k֨P��&����N>��3uѡVu�6Agcp5�Ɵ3�X߂G�/��.ӦM�-C|b1�Q�!�Q�{�WXv�@�����9s��C�C`�sʝ0pb�KX\�r�L��^�㎳�9MUh�ED�]o�����㏪#��F8��q��7��r�e#f���y�gٟ0����#����Y�D� �����Յ���Y�b������Nm_o��D�}��Џ�a�!��3fL�۠$���:n"J{""�5�C��W_�z���	��Z�]�?���ꫯ�D-����TOt���v˖-Sk��%�=�*(y�Tw��2d����jÿ��;y��zm�1MbS����䄽�n<������7D��`��`�ٳgK�8�sT�]"�x����矯f�O8ᄰ����k/u�;w��ɳ�|tB9餓�s�]E#�s��N���������A��^{M���~�3{"�1ة�����s�ת>��L�6M]�c*f��3qfg*о򨣎�8Cx�0K�ꫯ
g鉒�����z=�8_x�r��G�N/(?	1႞�~��Zd��]t�t�}�Q]�<���;���� �M�6v"J�D�Q�Y
f�����z�1}m<VJ�G�z�-X���Z��ו���i���f���壏>Rm% ���jg^\"f��.]*=�����D)����2ʳ�>�|�(�j|����_�3�<SfΜqp��O��.؁s޼y�La?�vZ��͕I�&������_N�B)'�n���k!���`ODDd%&w�}�<��srꩧ��mЈ��q��k�ʂ�,7j���yv���<z���(ց�%KԚ�/��R��"���`ODDAyy��{ｪ�%Z>bot���qqAgرc�
��W��u����͛U�w���|<x�j�9j�(�k7.#F��]Jf����?�\��`�Q�`�'""����F�H�r�3f�1�#S�N�����<ႅ�F(�A����U�@�`:�455�۠��4�
��}�JQQ��������w�yG�{�n6�(�쉈�b���.�|�4H-<=�Cd�ر]�O��:T]���Z-��_��܆(}1�u��-.ÆS����L�0!bG�d[�~�Z܋��X��D������(P���t\�S�)S�bU�|��'3�oڴ)�����c�y��`ODDg�� ]dp��`m\��u��vR;�������xA}��cF~͚5�j�*UnCD��������aq,�˘;�`�lp�Q�`!,.�f��Ѳ�nw`4x,��"[,��BWt���D�{1�S�v���zX;p*����v2�l`̏��-^$D�{`!�ƍՅ����W�L��6q^�W͘E��w]i=��\"""��b�'""""� �DDDDD�������(0�e {""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD������(	&N�(���Bɳl�2����L�`Oa�\.qee��~��n�x<BDDԛ�x�2i�$��9��d�ܹ�)�)���U���5����'����%DDDD?�DDDDD������(���JKK�P�)++��)����z��ʖ-[l�6??_�l�9(�T.���6����n""���^y�嗅zΧ�~*������Wۺu����¢B>|�u�=Q`�'""""� �DDDDD�����z����#)��+DDDD_�ֲ��J��"����;!"""��b�'""""� �DDDD��l��v�mQo��w����d���d���os�%���`�������(�de�dȐ!QoWZZ"O���فM��<F��=Q`�'Ja�55RW['���IQQ����1�����:������W��BDD��1�����z���V�"+A��x���Y���z3{���� ����yPV&�+*���E���z+{����$;vT2���W���R�m�Q슋��W^��3�y晲nݺ����O��g����믗-[���O?-�x�D)���HE�v�>�R�0s߬���(6���r�g������n��&]tQ�P�R�C9D
��f@K�K{�������""�]yy�lذA$�W��z�.�@��fJ�DDDDd�o��9묳�����)�������l�Y�;�C�9�9�sd�ܹ�����j�����_�~A��Y���v���`ODDDDQ���ʃ>({�̚5K-Z�n�]v���{O-�E�=f�}�Y��o~#Գ쉈��(",��׿�%#G��SN9%���~r����p����M���������R��1�QXEEE��SO�p�I'�v�V*++eǎ�t:e޼yr���P��˲e˄z�=�>}�,^�X��D�z��v�i*�G3p�@y����/�K����������&N�(��~�*���;j�/��B[�0(ظq���5k�%�=`c*̴#�������n�M.���ۢ��q�0ӏc���������,�}�ᇥ��F}���&3gΔ���ۛ7�B+LlZ�%�=�է�H�9E���!""�ԃ�f���TTT%�=��˸�$oȮ�߱�/�{_��=Q`�'""""� �DDDDD�������(0�e {"""�������9��ZZZ��pH2�k�y�{"""��m�69�Y�n[RR"�p�=�
��=��~�:��͋��n�T.DDDD_��_���Qz`�'""""� �DDDDD�������(0�����"<x�P�q:���쉈��R���^�.D]�`ODDDD�쉈���2 �=Q`�'"""J�s�=W\.F�djnn�L�WQ���Q<1�e {""""��`ODDDD�쉈���2 �=Q�����'�un�[|^�e
{�4TZZ*uuu�a0����ү_?!""��Dij���q�&�2������B��ۅ��(�0���aÆʦM��cY�-x��o�.����p8���(�0��1��)#0s�a�0�G�P�C�����2�=Q��̳^�C��P�i[�1��2&L�3�<S�Ő!C������!����Z(Ԏ�J�z""�x��̴i�ԅ2�}~~�P(���BDD��쉈���2 �=Q`��e���eÆ�.Ə�M�����l`��e�y����$]<��\@DDDd�=�M`�Y����������K;�b��v7wN%""�N�D6M�>]JKK�� -]���}�>nw)).���̙3G6o�,DDDD:{""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD�������(0�e {""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD�������(0�ٴa�����z;��+.��_��wHMuM̏���Q������lz�W$U:T���+DDDD:{""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD������.2h�������ec�V!J&��!Ç��}b����<[�mjjR{؅=��녈�({
�ϓ!#w���~��l���	Q2!�_|��q�Ϫ�*Y�n��ێ�u�پ�ٳg˧�~*DDD�0�e {""""��`ODDI7d��kz��z�ҥKcZ3Փ쉈(�n��V)++��-DD�"??_N<�Diii�T�`ODDIWXX(+V���۷Q��1c��?^�ϟ/�������*''Gub�'�tSWW'�w�=�}����ODii��ղ�>����L�:{{
���V<-u��F�'�}������g�x�b!"J7���j��뮻N���?'��0�Sxk�/C
�����6	{�����R�����(-Z�H8� �7o�̙3'��������$~�a��Ζo��V���U[[�,Y�D���j�q2�=�=%�̙3��.���*Y�p��;�y���UW]%S�L�{�')���������������C監�:J���d���RQQ!DD��_��L�6M^z�%Uj�駟&�10�Q�\~����x�%��'[�l���r!"�Dب
�~���r�5�ȯ~�+y��7U�O�|�DD�m�j���(DD$�i�&u2d��p�	�_�B�m�&_}�����S�=�������� ��.`Æ��?\�?�xq8�M&�`nܸQ�&�_�^��Ÿ����X1�� �� ��0`�Z�4y�d�7�?:�a�+�[\�z�)y�l}{""""�۱c��D2u�T��b�'""""� �DDDDD�������(0�e {""""��`ODDDD�쉈���2 �=Q`�'""""� �D6͚5K����v�Gj�jm�gaA��F:V.��j!"""�1��4x�`)--�z����Q�C��_�_J�Kb~,+W�d�'"�A�C(�|>�P�1�Q���z���5$T:�Π��a�|��	w;�)�3�ǆ���*.*��!���2!""J���v���U�>??_���%˙%�G]���_ !�4�nw�}�q�e�f���}��ʲ��4��?�c	w���Jzz��?��8���`��`Oa5VrJ���~G�""�djll�ښZqe�����YNq:��pj!��o���3�iq4�k�z�}^�jG�q�9�O���?V!R��>	��_� �۩��g|L��D\^��x����`.d��^���=�a5�п��:���%�(������q�j�g�'""�^���Y���T�mhhPA�T�ػ���*����V�a�aZ��D�����*H�Ɂ���q�&���D�9B>6��Àϑ��Vg �o�lDH��?n���:��Z���������}8��G��yPb|VgI��k��P���\���i��г��쉈���@�����ֶV�.g �a?ۥ�u�T�CE�7���y�+,����#��A_�j"�u �Z�W�>���Qn� ����>ogP|�3a��(�Τk?��Ƴ���y��Q����-����B @1@�v�+ED�"^l*͊�� ��U�+^A�"Mi
��A:*A��JH%�'����g�ϻ�ξ����ٳ���o>�ݝ�}gvϞ=����}^G��T:����'�V�^'�iqG0�k���Rss3����w���C�   P5���
�ejG�Y�e���a�g���N��22�W1�YX]�W]m�����˥n�#↚$�0H�K4������d�o���o��z@}�R�S3���}�#3���������0a�!���|"�{    T}��l��z#d^I�	C"z/So,���@ �c�i�Rp<B���@�9�٢���)�"R���H�Q�I=f>Q�Bq�j�p�C??��h�j�XD��$��Mvfv��!�iii��.5{    TRPy�FD��4,�"�FF�q����r������F!������V��z�Lw\'�W;R�Ћ��_�i-'�O|����.���Z	�#���c���=�oq'��s���J��ollL6Ub���   �*`Yc1���9@L�؈�Χ���F�V|!���5�օB������ܫ
-�Uq�U,�w��tn��R���8�S_+�?��gBVO�c��x:RWW�H��ϕ��=    ���"�b�ٖ"���Ȉ�zQ:шwԒ�j���H_>"\H��\s�L%��L�޶���;2O�J/�LJ��ׯN�+8c�+7��#?�BG�Y�y0vGGGN�R�b\y������ힷ��+� P9��������?v\ZpժU��  ㍌���Ԋ�8&�D��*��z-�D��\Sb��p�|�_=�l�����u;I���K�^�N�幊R�<9��b�zQ	(0&��{YƓ��y�������=p��"  �ħ?����K�_����O��[��[o�E �7\�p���}b������ѱ��fY�x��W��H�U�3�$����f�C��9�����8�6�6m�g}�����g,���+���(	��FĠ���	~}]]ɣ�{   �G�n��fz����o��Ҋ+�񤩩I�:[_��!!�r�%9�N��U ��E��mVT��cU�Ѫ�):n)/r�z�-Md��1��}�}�̫�r>V��k��g@oC�=�Ā���5�5־�b  `\ٵk}�s���ﾛ��cZ�~=0^�����GGF���c�$L�H�@+����	�i9��닜�5��WI��|]��"���|$;]��?��x���Λ5`���C��r1�R�  0�p��/��~�_��Y~���qX�X��Em{9�̝�p"�5aQ`,^
S�g/k���=7��n���	T&�R�)>N).����C���I�IR��������Y3`���������>�ԝ�= Y���RCCC���@��./��r^���� ��ڵk���'��>��k� �	���j�>�Q�Mq�4G�GFG��<>D�]��D^bE��U5�VMG���yN�wu�Ufd�}�Y�S��ZI������{!��r�cf{�n�QE_��TE_8����R� K^~�e�ӧO��������Nw�u�,�.�x�����e
��Ɂ��g��WEI���Z�2�Z�Lk�Eߖ�!'�JLp�F�-���wJ��Sz�+��ؿ@4�&�4(VO����:�+nc��٦C9�?�3��)�z�M�  �:���u�hΜ9�& ��E���J�u�YfY踬!K>߲���s�����gُ���"��[����D�|�<��[�b�j��ӟ���S���yn}�$��jC�}��3���j�}}����\s��˟��r�Z� �   Jʣ�>Jg�q0�8U�QYϓ����q'@K���˨��~.�908`��Ev ԫ <��\(WD'#!��s �>�.�����+~���T�<=گn�����vl��k�}�~>��\�
�o5�Lϱ:��W��  ()�<��{�@)��X��j:�^��mB"^'s��N:d�_ʾ|�^��|nV �r��3��W ���r�y�筞���̨+� ����H�S���q�����:m�l�>��[�����_r�  PR8�Y���4�.t��TYe����evʹ�eVv �I�lK}��:���d
��
 e��] ş�
��`(9�n������GF���3�Z�(�J@�ye�c��q��ŭ#��|"������~b  ��p����f���" J������Xy�9�k����)*z^x:Q�{���F6W�vٱP������8�P�tԚ�2eH��u�� ]��s�"�Շ�)�+'^�ϸk��O�C�  ���_��8�~�3a�#���m=r��M3ɑM��نz+���:'�X� )�|@�VүH��J�|�����4��YPS���QS|��!��f����v���sQ$ �   JWQ�XP*���1=%t�T��6iw{��?_�X�r�M[ʺ�9��������F���u,�}y@��)@��9V��=���)���J�D۩C�G �   J���	7)�7�Ct�65]�R%�N���g[�àQ�:��Ls
P���U YT
��Ȁ�s�����%AE�Č����<5�F�z���P+�����$ܭ�_�={    �4x���Q��|s�+
ٞ�R�=J��K�w:o������NW<�����`N�SS�d��
Sm]-575SCc����9� n[�pT쉢�6��    `(f�&�F�E�3R��w��8\)Х^J�:����.�����@��l�?�}M�0!.��Q#j��S��g{5��u�^�/��    g
�|��B�F���S��"�ߤ�����t��2���������nھc;�޽��M�f�,�#+�T{    �2$���ٴ��@T��Ƚ�|��w�j#%]���qyٶm�߰�f͜%��T u�m.��6�����[e� �    (c�J�a��
�V�'�Fl�AR�����N�J�v��n�=��A���"5��q��     ��
���L)�I�}f�L�1�u���8<`6�~�ĉ�ώ�;(\���tzm�C�S�^�S$ߏ@�    ��B�թ�~�{�����,��-nW)u9i�$Z�v-M�0њ)W�ܪPr)�YJ �     �s��F�m[n|e�ι�����xE3J3�����;�*��c����ޛʅ}�ݗ    P�x�W�^���ί���!3/�ɷ�a޻r��t@쫌Y�f�    �\p��71i�\x�Z9�{�I��y *�=     (�轜����&��������s�b     ��j;�ƽ�'�m5H=��py�z뭷�Rx��	    Ս-r�X���c��z�O��5+"���p�}�Y�     Tz}|�3g��r�!� ��$��m���i�<!J]]]V��X�����Y  �)��^�Q��L�� � �����׬YC   �Y!'�n�y�����     e���U2XVb     *
���4�JH��@�    @šNd%#�z$_�J��C�    @E��>kVA={�=     �xt��Dɇ�    ��AI�gy7��H�     �S^}���@�Ȓ#�8�3��_�pv�Z��H^#�l�B�#�   T;Fb1�	��Z����7n@�Ȓ%K�P{{{�����h��+�js����&�|.O=�m޲�   �j�)�n��6']��rb     ����m�ܧң��     ��ԛd�@  �q�6]�^Ͻ� �     ��b���266F�`ȖO_-���=     (�(���S\�#��B!�A+b�>�Q%�Ҫ�@�    @Y�J���z�x``����(LH} U�+�=     �5zT�ŝ���6!����4{�l����jb     |�S
��o$�ސK�qOO��ajjl{!��]�MT�     ��8ɼӭ\�	��A�;w�9s�PMM�|5b�&�f�B�     �eϧۭ�F�J��r�y�fjkk�֖V+�^�:I�� �Jb     �"]�]��K{R���2X��s�~�ƍ"J?k�x5�`�&���    �
ѥ��(;Ɉ���cj�yu�bmN�@�-[���	i֬YB��i�l�Ԝ��1��K�    ���&�=���x5}&�\��v�u,��O����{̥��V[�\'��f?n/�:��'�=�    �L(V�[��D���}@��5�s�}Y�GFF�����'����z�������ԛPPLF���{�[.���B�    ƙ��^(�(��B��)4��R�
:��[�>o������Ԅk��7�7�ׄ����jkk��`@��T��#=ƭ�xڑ�$b    PD
��;>_X*sгi�)�ީ��I�����S���r�v^Xڥ��%[�񁯢c�Hoڜ���m2�>�ԛlp{���o�{�= Y�f�ھ}{����/fÖ�[h��m9�K__  ?
�ty카�4Q�[:M.��f�'��tU��(;â�r.�Ǉ�T[SK��V�;��H�	"��ٗ�)S��Ɋ���r��̯�c���@�Ȓ|�����ө���   /�7���DƳmOʤ^)Fo'� U�
㶨�nE�c��b�����`=��)�(�"�V�q[8B/f�5(�=����~&^�ثB�G��(�{     �L�Y�iKOu�#ιT�1��Qw�cgd��Ŝ�ZX�y@*G�嬭R�9®^�vz_�&�J����鲯�%�s�\V��ePo1f��m����{T�    �!�`�E��q�+NR�����Ք]���H�	�X�1���"���ɛdjK� �$�#�j����HQ��;���kr�z5
�֡ϥCU����}#qy=�    @�$��s�o.�J1Ts�������+��\uta��d�y���c>W��ޒy-%(�vt����T�/uʋ��4�J�    U��Ȫ�uQV%W�a���S#�I�c�.#�R�mr�E���g��mB����y�V*�ID�C٣����W��}I����qj'ݱ��Z��+	�L�AU     �$����-]��3rЩ*�Rإ�˔y���Y�nyjn����îW�qJ-Q[��?�&���<�wjo<#�z�D��8�����!�    �N���<�)߲���c��(c�M�N�	�X�Qw9(U�
#��tlF�D�Ψ4����>�kR�qw��s��ug#�~HkQ�+���q�gA,�1�saFK�*{    T%e���R�3���Oc�^WW'"�,�|�N�$��9�]�8�)M�M���2�&Q�]��&�z���^.i0N�m�K�v����\7����U^%��M���fF]_K���   �����.1 U��X��ZW[g�ͨ�2B�% ��OS"�J�[�^Oyѷ;��S4ܵ��8��o��M���2/�^���V���O�QӖJ�3��   ���ݻw�2o	{0`E��."�ʀV���LR.�%5%�A��䥻�KN��<�+��0d�!�"mH?��O�*��܏ERRsFFG��]~ b@����G===R���#  `X溺�Dn���pr�Ә$�u�Y�e�߲��uR�꼫�I�8��ӽ��{��`KA��M&�ש_��Km�6єIVꍌާD�G#"ukhx�FGFE����L�81��+&{ * zH�;\�b�)�}�6 T7}}}B����uV�=`����"�^���%]�E�y����g��S���4�+�����)P)�5Ȫf�y�r���H���1�d��z���P�QHG�+ � �9�}��յ�@zx0ܤI�h�Ν �^8�:K�ۮ���$�٦}d��L�x��,����S�Ո7#��I���9�[����~<X�p�2P6:&��2b�2ϑz�|QQ)��ɓ&ۣ�ȱ �C?�ܵ�@v446R{�w�3 �!g�#�1��(=����BA{�r�T��N@�Yu�VkΫ�\3�T�P���,K4�s����\"������L�|���1��yN��3 ۢ���b{d4��k���MD��+ �b@�280H;v��ݬw~���I|��9 @u�R�B&ēR�}�
�3R+�Xbo���4Lk5J�����8ɹ�߭���!�+�#�ЫeJ���>�i��Kt�����,�C��ف9z?��#F����Ԋ�}��vjnn���?/�= e��uvuA�󤹥%����� ��"��A6e=rq����Q+�oe>��c/��K�I�g�J�C��+j�?_
��KKNӄ�4d4���P���|(�o�ӹj)W)Q�Ĭ���*߈�B�g��+x^�Yhz�t_E�%{ ���
�'�1}0�	 0~H��������Ǆ��N������uR�ժ8������X��GM[
�:�m��N6�<We\��SSV�����HA����ի-No�i=�kd�7�X2/>\�]��R�PdJ�O � �!Q)  ��K�([����RHE��H���`(H�� FS'��MJ�T]I=�������M�0ʒ��y!O������ٰ^���[��l�e� �>������+�Jm�&����K�u?j�ҳdǎ#��g�y�FM���3{    T������)�)�q��x5�c��6F!�r�*N���\�6c*�&�� S����r�ت�©,J���)�5�	96�dj�^쓸���.�꫶c�W��@�!{�՗�����`b"1"k��d)�O.>�'#�ߪ�Y�5�-Ԫ��n�{    Ty�(,OB���+,���s�Qc�81m��	�z_��\��e>7#��4��6�o'���X�:D*QBZm�j��I�~JD�iЯL[��k�[�@�@o�mN�z��`e3�2%r�����a,m�N�~b   ��b�ĉ�}�vjnj���>�Ds��@$!�FrSYIE�0[��T߶��\�>"۷Uj1�����$����Rf�4M+]$�_:�VZ�huW���K:L��n�W/Ȧڌx�y�>��y�n�{    T,��'O)9B�x��(mh$��Ydc�e�{!�A��g�"�)�/�p�*��E���l���t�)$R��b�\�1��YI��Zk���=S��է�t���ǺD��.��   @���˳Qs���O�l�.�,��<��-�D�w�<|5�EY�1���<�[�~}&Y��_�tFf�˼
�  @�a!��0�p�}}}��/SZ��;WZI��L���1�4�
-~��\��S�@�  ���QS J�>C�LCQ���ڧ�TIE�7�4Ą̗{   %�'& J����.cVQ~7(={   %�k���� ~@��Be2��=  ��"'��{�y ���{   %e��Őz  � �=  ��r�q��g   P{   %eɒ%�b�
  P{   %��SO����	  @a@�  ��P(D��~:���[  �p �   J�c��;w  ��  w.��"�k�����'   � �  0nL�0AD�'O�L/���ȯ  �{   q�%��̙33���� �~ǎ�t�RH=  x�  @Ar�!�m۶��Lq�z(� �� �  P0[�l���~  P: �      T {      * �=       �     �
 b     @ �     ���     P@�     �  �      T {      * �=       �     �
 b     @ �     ���     P@�     �  �      T {      * �=       �     �
 b     @ �  P0s�̡��Ѵ�����;�C�H�   x�  @A���4s�̌������N�w秊+WB� �c �   
�'?�I��644ЕW^I�z(���K400@   �b  `�`��袋�_�"�t�I�t�R!   ��  0��v�m4y�dz���'Ry   �  @I��{f̘A�6m"   ��  P2���:��w��  ��  (���?hpp��M�F[�l!   ��  PR�y�:�# �  P {   %塇��;�   �  @I���@ @   
b  ��p-���f���% J�a��Aq1M3�c�{   %����!���H��[�����q:���g�  @��P�@iЅ^]����.^�ϔ�g����;�  PrX�gJ�[�exx���h�L��KU���|_�����K׆*��`0�����+������ĭZ?G}�߀�  (9�R< �K��]�hll�F@,��Մk(��bK hfK�yc$�4֦վ���u���ĭ�O>���}Ƣc�4�mD"�9�y�����$���P;j'BoO�/�c����XR�ն�6����W�\M�K�Cb   ����xǎB����B�Á��������a�`\�����
�4����;*	w����t	���QT��1��P���Vd�ꔨW7�-�ޔ��<[��JiCtn���z~*n��LWF��rd��">����T^��_b   ���#�����2ǋ�pH,2b�b/"���域c	�aX2�M>��=۫T�
�[[������#��,�ra�6��աI�ܿ��Ԕ� N�%/_p��Q�i�΋lO<?�������i������ZZZ���N|��}\@���   �jB680��������h}�&.���%��WSr�"��䞅נ�R���:�s�mkB�Z�
�����������Oy(_�ڑ����SWg�FF��������@M��{    T,�2ם}�#��1��0|k�z��R6D��0l)R�3�k�H��_$���mɽ"�"�m&�>l�-�uz-��*Ÿ�B�J������>_������:!����b�:uj���K���B�   P5p��ёѤ�J�������,�$��y7�wJ��D&	N'͙�eJ�ѥ�JWQ�Ѧ{����Qa����ʆ��	xPu0`�-�-i[|�St�}�]�>}���t�=    ��5��E�l��`O!~�sJJ�)��/ɥ��7���|�*E �͟y�F~.8]����5��u�V�1s�չ���M1��   �*�M�.)lb`�r+#�R�eN������U�3��d{>�"����tU�%ls�Z��� E�d�qe&�>;��G�T���H|�F������Zr�g �    �
dE$��{���2���~4/�hD��2�Z�[�tk]������[]ݖ�|;٤��\��/d�t��"���r��E�%�g�?C�o�i9===B�)�NV���߰��Z��A����ϭ��F�L�����K�����?>�C   JK�+�"#Jm���	�b��}$^�Rԧ�΀��5W��ʭ^S]�8����~�5����l�f�_hdYp+�܉��&�n8�6,��keQ#�9�aSTLb���cTZ ��7,YPO��r�3=��x��C{  �MMM���i	���s��h�N�%���沖��bN�h�>�VNb����i �ڱH'�j�_�xd#����Q�B�t5C/Yj�6��$?��V[Wk�}���=    ����Z��������=�|2l'w4���hM�t���m�Y���Du���3��Rc�D={]�3��Ѩ�8���SI�u�!�މlR�2]9���W�^��9uK)yYJ �    �*&L�@;w�ƆF�7b�Q���Y�y�鄂���+r/��'��[)��i�r��S��u��;��l[�G.�m�����D��6�����S�9� T U�]  e�WGG��d������쪼p�{9��J
	N|�Kq�Є.n�VG 
Z3֪�[9���c�ꀞ߯�~�J9��ZeӤ������v�R}��Gp�i/݀_����r�ܙ�)U�=��?N@�("S&��W����-ZD�V���NL�<Y�aˇ5kֈ(  �3\ɤ��Y�F�9�r�Q������L�s!�	��y��Wኈ}B�j
����̥VG��4��?w*�m�0X���]�d*P��#��c�H�Q���}Q�;E����g���+�z�%�f���?S3^)Iv�,��Χ�@�("Z���SZ��������t뭷����O�6m��?^̐������?Q[[[^�8��hŊ  ��rKKKJd�c��	�Xb���߫|˲�F��"�FG�<����`H��'���'G���ʙp�"��׊t�@�64��}�mu /�mp'H�VrjC_'ѣ��.)E�ґl�?�)@�(2�>�������-���K��k�Rϸ��?B� �jǩl����ɇ�Ɉ��v"�Oʾ.��Xv �>##�"�G�z掀lOD�U�5���,�����\r��R��4ly,3y�8 +
Mڠ�ĺL�
��YPR���zj�S@m�m o&\;7Z��/�4���a����8�wǥ�L���1zj�@Q�u�y�ёG)�s��s�9G\^�ٽ{7=��Ct��'  T;��ˀk�Ny�PDl�"��Y�Ul �{���Jv �����J �����4��UzBA0�S�PSjgEޗ{X��* ��c �&�rJY�S{�Ы篿N��:�}WS|+e ��*Ӥ@ٱל:��T�c_r?�Vu�l�WV'7������>�z�ӟ��֯_����N'�t���v����?��G?�Q���  *�
��URM�(��~���U �i�+�� j��[3�ڪ�$D_D�#�ȿ3���p��s��5a����P�r&���O�<����ɩ�9':
�����@r��^H��v%@��U����̗J���@�Aə==L�
���{V�B�	���L��\��V�!/�	W���j�K�^���/�s֮]+�;����Z��ͣ?��Ϯ�c�, �P�^}�X��|�"�6�]!��nXҎv���oY�m�@�dG���6�� ��d�}Y��I��&jod����x U����צ�N��L⨿^MȺ2�G���K����g��J(�	�%eִ�����ޖ���hl�u�M���}m����O?��M�&��4K~6�u�]��sZ΍7�(�� ��ѥ>E�lWD�)��u�L�W�Qoe:O m�5�m)@#��}5J.nɰj��J@< v_���Ubb�-:!\(�����Z�{m�D�e����n��/���Y\��9��f�*C��ګ	�=()'�L�C�%�z?��&��ݞ��$?����g�s�=G[�n��S�����詧�"   q�f_ͷ-�ԞldT=����K�E�ՈxL��55�� F\���i����jl��y2/����� ��	����0	��ui��d����2�k"����c���EIt�h��A(��= F.b�_�<��t˜r�){  p�+�s�|��ip�L���lO�q����·*����e8b]��Zx�|}YH�1�~�4�� �U )�r�s���b� >?_L
�NN������= W���g��/������۷  ���U�v�-׈�+z^��U ����t�^�*�}Iiw��$�ȫOL�œ��(��E� ���/&�
�'�b����P�#"g�u*Q��>TH���
#�A��7o�W_}�8� ����8��?  (>�J���P��f0�=ΦDe���q �$V2����-����vxd����������phX�=w�uVGBͷw�WM깚H� �	}��l��_�*Ğ�4i  (�D49ud�����I�O�*��U�	�����<OKWW���Sccc<-g,>����0����+'~b@��O��۶m���$  �� ���`+J���Ċ�mQ�j�>VC���� 8�/�r&r��BcV>�א� f�����rA����1   P9��v�_�<��$&�J��'*�� �9s戔���AjlHD�r�1�LdUn@��0��s���'�   � ]� �+ b0�2@�Ysƌ�a���å.���:p�-�F_��DV~b@�q�1�г�>��s;�0�>L   �����VZ����˔)SD䞯Z�"'��}>�L9�\3ߏe2!� T���'iݺut�-�d�?װ?�裭��    �@:qfigX�D*���5�5Y�8r�+��[U!I:��mA�(��I���F�a��-��?��$ejk��H�g�m�����=���ė�m�������_/'���ر�    ��N#s�9uh0^�ٚ��t���T ��b`�k<&f�������J�=��R��w�o㋜V����1����س����t�GX���oӱ�K/��"uww[_�,����b2�������C=D��?�C   �_Q_���i{zz�|Ӿ�q��J�~�=�x^~������~�]����~�/��cאi���\����ϧK/��N?�tk�Œ	�b����n�r4  ��P�krN=Wő�z!���LmT{P�f &��T�}ǻ��/�Q��_fW_}5�^������]�̗��s��ӟ�����\FƄ�  (!)���c�WMF���Z��؃���$����=���K���~�ZZZ�����I��z��$��Gy��Ν+.u���   �)�)�{�˾�쳕�Tn���כ��k��������=m�'����   ���;S<[h[e�T.��Qʃ2K�   ������+�g�	�=�x
��6a�   @E�i2�rb*��SqL��=    *k6�
�{�=�xL$�>�`��W��I[O>�$�}��   �!�F�.�\b@����~��_�T�3��/�  @Y���WB�b@�3g�1��WR�<��c   ��JK����
����n��f�8q���{��/�Pp����   ���c5�Ưi�{P�T��t�hjj�_���4c����k�E�  @�c�w��"�jν�=]t_-�i��{P�Bz���SMMؾ����Vt��Qփkjjj�n����O<���H��~;   ���b���:h6��;���]v�<�؃���Ɍ>c�h&��4�g��~A�m ~+b���}͊`0H�\s-Y�D<����NW]u   ���3͢m[�H}�m��=H�w��}ԤYQ��i�
��]Q�*`����6�����}Y���{��s�1���իE^}$!   �R�E�))�L����[5Z�$���rb�1,�#=���g��z#�����1���FSa��K�g��/��Aeg�_����SN�w��M_��W����   �J���η	i�	}��/����u�L���>�t��{����B�����.���'?��o�w��y���?mM@5<<L�{.m܈�%  ��B͝����&��Y상`b}��	��G�ԇ��_��t�H����f�#o}$6�h=)�z����������~���cN�Y�l   ��*�R���3K}(�G�FE����� ��& ��S�ϨQy5R/��0ʧT&��ɨ�Ν;	   �$�"����������("!ש�,%f�ľ@ �>�%�n�ث�[iy��'�)'�g������>�1��/�K�o�t�R   �}��L�QoY�9���AD�Y�e:N5�/ H�����9����1����> �`���LɣW��H����7��}N��SS����?L�gϦ��?_<nhh�_��Wt饗bR*   e�[�5Z�z����m���4}�t+b/;NQ�Jb�'�z�1��hp�`��6���zW��?T��c?؂Ω!�+��@��|}}=�y��1OR�����Z[[��   �A!�����z	G�GFFhB���Q_����H}ya8��8�ۄ�L���k��8�]q����D��z+   ^��|���$�*�Vn��}���4m�4
�C"'��W*��ԗ�dӆ�^y\�B�r��׋��_|�����o�E�=   �Rh�Z�q�6���c�^x5J/o�}Q0"�'~֬Y"G�gV��A�s R_�X�fn"�1����������N��(*0�s�Ƚ��k���  @�L����%E\��C�y�CoPj:�J=���e����fb��[#������,����_�O��Bu��W�l����1����g�ݵk����z���<-X�@�/�|��y�  P�;��(�w����4ٶ�v�TK�)^�~˖-448D�-���&!���YŒ��H}�x��!��U��˧P}	�c��pX�/�z������]��szδi�ĺ%K��.w �  0�xewKy1\��Cqu0���G���H9m=�<��Z�\��s�8K=�Ȕ�#��ү+�y��ק��!�����o�`�v�$*���~ɝ�R���Kz�Ûo�I��v����'R��*  ��(t`���B���~�vd�He[��o��N�v��~.�cy���Q��̏�������������߇���S�5�9���Iͱ�����=�@�� �?X�9=�}T��J�%�z�e0eԾPv��A   2�V�݋6�D:[���\��J��i_y��z:�~N,�r��η,��N����c�jjk������9OTzS߃t�,s����Q3*n�^���ػ ����D���zA��^�_���.�G��,(
Xj{��q���e<10U{�t�t����\�i����>����΂�H�\�#��3����ۘ�775��b�I|M�F�̫��5]�����=���K��x&��{b� �x�� ����?��lq+��϶-!����|v���\�Kc)�rG�U��e�`���)�r���yMS�-�.��;n�3�:u:��N��٢w�� ۮ��,�b��^22jB���  JM���Txɶ-� &nU��'O�jW{�� Q=�iQ�]F�9�^Ә�pMX����d��9�N�C�~N皩�.=&�Ύ��c�(h�y#`�.Z�@� ��k�Q|� �700@ �]����L�B�V���ɔ�v\=��$�z��o�=���������+����¡��w���y�N��������X�ڒ�y+-GI���Y�� ������. (�d���"�������)}�-b�N�ݢ��:�躚ù�c���\��ƺx�=�D���į*p�P ��TM'��V����n)8���v�1��Ye�uJL��%�z  ({� J�.�R���z�=]���I읤^nS��n�0a�J1VzL춮��&�*�D�ӭ˕l�/�}��+��TB3�sRSq��4�?����z�jI��z��� @i9���ń3 �
U�墊�S�7���y###�z�z�]氇B!+��b�%ET=�r�y�S$]��W��G}n&a�$�ْ�S�_���j��>����8�+B5��B��/EĞ���z  (=�~8�_�� o��^�z��Dʞ.�jv����΂�b��IԔ���8�Տ��J��~��Hw�v�>��7��V�s����?wqL�����V�!�  Pz�>�h!;���
=��v�u�g�SbD
Lc�-®�ĨQ�l�<�W
2�.�=��m��1�+ר�ɖb��g�|��tyl�~Ñ�H2R/;pb���^F���k_�b� ��Ñ�s�9�֮]K �7R>���C��(��Qt���z+=FT�ID�e��U۔�K�$���i�m�ҵ�UU�b��}օ^{����ԏi��"�ruJ�>T��C� �\u�U��-[��?{�v��&��^H��w^��
����}^� T��������)b��oZ�S�]`����X������i�lȥ�|��U���k=:o-�yK�m�d?2�/��`esN�EU�=��7~�� ���o|���Z�t)0ް�q������2{���.n)��/��N�1��Eϗl��=G?�t�_�:!�c�΁S��J$d��_IX�����z���"oFmm�>oS�W�>R�9:�y������5<2L��DjV"UGΦ[j����ԃR�sz�6���_� (����L�B���?�J ƛ��N!r}�}"�F��V�2���d�w�\v�H���9��E�3	�-��A��0��<�(��)Pnǔ�82b/Rp"I��|u�/���b�s�����?Pb����T~u�T:�{P�pJ͌32����'�H)G��V�T,ai���b�Q��1�����٪Ȓg���w���r�� ]ĝ��Qp9ϙB�Hʧ��_��>�U�ƌ�Ȫ���ؖ��1X�9}��=o*^�!��C(X�i+���@�AE�)5۶m����-[F ����~1��-�=j:��.}"��TJQ�᳭P�&�N������d�kG
1G����B�[���&~2�JM�4>o3~��#��5<��Ɗ�8�2N��H�����q�������R_>46hɢZ��a�D �����,L ��6!S�dTYF�Ձ����ɔ�Vk>ƀi�l�E���v�|JJga�<��x�z�S�^V�����F=�����7��������X����-��� u,�|/�-�D��Y�쿶�L	�X��ԗ,��_1�ښ�-���g���?�h@� ����$-Af�z��Z5�Y���y�r�l�I"��T�2���nz�]=H�e�)?�t
\�(�"�7��"'n�`*'����&S�u�M�)�਽mfY}�E�!��9�<n�/R�T��C��)�����n������� ���&�U�^`$S2d������a�<n���n�^�t���j�L��"g[\%����>�����Ӛ�5�9bY���k���R6S�x�t�#	���ȷmmmV�Od���R_^|�S�q�/"�"�����K�Y������w  ��#�2Z���"�B��T�Ϫ]$#��oD����7#���
���ш���UWde���o�������ێa���E?2���@��	L���v������X�yP�I���gI���*J�!��GM8P�cĿ؜?�����&�'_¡�(  ~��3��Y����1G`)q�؊�#B�E�?�O0���J��S5w^KM�I�E�<`Ӄ?B�H���T�6�c$��l�ɫ
�.%���N��Y��S_�A�Ι-��tu���Qccc��g�Q1b�n�t�~y���z   ��S(X�m/q�}쟸���H`$�����-�>C$]s}Q�L-i����e
���ɫS$<�R�|�x+��Uu��8$�ܪt�Ll�jd&KX�}�ف�����i1�2�B�W*B�!� -	��?⊪zy1!�R�!�  Pyp%���3��ur�5��Cn�N.�ێ����6_���7/*�1�8K��n�IR+�0R��q�H�ܦ�So���m��3z�L�%C�2̲{H=�D�%b����ddFF��|�  ��@����Eu�u44<d�.#���E������Hp"�D�n�(�<G��0jU ]�����D�3Eĝ��u�;�\�J���R�!���r�E�����擉�  T �/�r�{�njnn������O�6`T�u�9W��6�N��X9ކ"ݦR��t�J�YgՊ<�,��-�Yb�r
I6bn�s^���)B���\�U�G�l�R_yBT?�)���>�CJ>�Dx�^Y2�jcX)7��y��3��S4h�   ��k�9����T[W+��ZF�fg�`Z��c"",'��G��b�:�i��\���+&����<��Hw�P�b��P�Tߒ�ˡ�s]��s�ޒw�bS<$��"�'v�~J}��4ʽ��  �?X�'M�$ĝg�f���Q!{4>����"�E~v)�B_����C�A��#��5�ΐ�F͸�Gq��X	�-T�  P�p�JCC�m�S��I��D>�: �AY�=���ؘI)3j������X�crϱ�{3a���  Չ[�|��xQ6b��ۮh�ԃ4�����+S���c��q��r/Rp�N   �H:(�B�ԇj�K���z���炫��b/ʇ%r�9G>7ȗU�DG �z    ���T��Ճ���3��m��	G�@Y�Y<�>�X�\�=g:�    (|-��z�o�o�����̲��Csg�D�=    �ߊ=�xO�1}�tjll��9o�&    �rb����    � ߉=�     ����C�AQ@�<    � ߈=�f   �2#
�Y�sz� H=(&F ��P�&    @1hnn���Q࣮��jkk��3�ã���iӦ��+��C�A����d�    �[&O�,���&!�,�7o��+W��իi������o��~I�R<��č<��z    x��3hڴiB�{{{�Ŀ����s���Ȉ��*��C�׸�8�(�W{��   �3�N3�|�f�2����<@�=.� H=O�<k��ĳ�p��L��I[۶m���p���F����O�֭��� �Jd�����3gҚ5k��+��6�۱�]�!�`�	�1x�#��rt�UWщ'��I{O=�}�ߤ��1 g�u���_�>餓�����aq9�E  *�<�������=�\ڸq㸟ø�=��ԙ��Qz��;(N_2J}�@�6�/�R�_|�gR�y����~Wt HGWWW����'?�u��կ~�>����b��. @93a�z�{�K=��t�M%;�q{H=(6n
~�~�t����s�6���F�M��>�l���?�y���v�H�)��<8%����'���������-  ����Z�h��W��Gy���2.b��$�a��G���K�/���O>�����������-[VP����_�R��s{�v��￟ ��_�.����OJ���H� �%<ƈ��z��b��E0`PM��4�����G>��*ö��^��}����'GA/��R��_�Zp���\@�]w��������M�?�8�%o��=���t�A��/�L  PNL�8Q����/~A~��b��I(&��#�n���|F���Y�fѵ�^k�P����}�Q��������_.��87��7�D��n�A\��{� @�0{�lz��'�/M�!� ���v1�4�]�s�=���{北�>�=�Pq,>&�x��А(ɑ��;w  ���K/�_(��C�_˲m $�_������* ����o��6���R   W���/  ���T�!�      ���R     @��D�!�      ����R     @�)H�!�      ����R@���~�     �$/����ؾ3B��o����y���v�߻�����i����%�&�w:&    �E�b�^����MS:Bt�q�T��n��ݞ��b�
z����c������[�3��uvvz�~kk+�x㍢m�駟��+W    �INb�^���޼K�?�cmTɰ�_��.���:/��b���iɒ%4{�l�կ~Eg�y&�v]]�hk޼y��k��F^x!E"�w�   (�{H=(R���[GG�D���R/��}�kt�w����E���~�;ڰaCA�Ι3���w_qժUt�9����   ��d%��zPl�#����W��K�%===t�Ygѝw�i	���Bٲe�w�y�    �7�R@���=VT��p^��g�Mw�u���{���ݻ��_���{    ���b��0�����7
�?��<i��G�u��    �W���P~���b   @��(��zP
�Z?L���nۺ���Ҟ�k��X�n�V��O@�q&�   ���"��zP*^\9(��� ��LjmP9��t�owҳ/Vn     Wlb�OOMM]}�մh�"�+�=���G?���]C}�~q����z&2�?.젋��A�'��/����u�]GӦM#��eJ��   �/��C���R��ґGI~���O���Z����O�h�ʕpؠk.�{�R�����:�?�N�\>HŢ���n���1c���{/�v�mTnL�8�n��V�{���\z�d�|    ��C��â|����a�F���'�,f%�ꪫ��gt�7'����\��1��ߝL_�j��zq&v�	�>�`/Z[[�����[n�ŚA�ϰ�_r�%�w�{   �z������K�/�ԧRWW'���r���ԧ(�]�>�6t�9����ܩ�5�?�3��z�6Z�����X�����f���CSS�M �ƤI��7��MYH����{   ��7�-_��'No����~��_Ӓ%K�)����>?�>qL3U
M���S��m�7�z[!��_���ޟg����(�Z��n��ƌ��tWRnL�>]��̚5��D�  �K(��#�u['�^�#�7�t-^�8e���(]~����+��_��G>B��ַR�s�)�?��V��'Z��hr?�ξl+����v��{,�~--����1��~��{���n�{�i�&��{.}������{r   [BRhnn�����v�~322B]t=���'8� ��s�)����?�D�}fU*\���WM����~æQŁe���I=�̻|�r��]v�i��f[��   ����%G�ݤ��.���~��G)'��Ər���7�e緋��Jfb[�n����w�Җ�޲�{���)S��l��줳�:K� ������@�w�{N�a �   2�W��_�pa�6N���K�M�߷�����
RU0eR(&�����vt���=��ST��<yr�6N;:��3i����W �   � b� ]�롡!:����^�r�����SZ(\e��Y�Bt�Q�t�}�	W�a��Җ:;w��z?K�r  �P�L��iooy�Ne��_�j�H���2���\釥�g��ٲe��Կ��;T.@�  BՋ=׺v�������Σ_|��Ƚ������Ġq���6o�,�~�ƍTn@�  �KU�=W�`��={vʶ��^��W�B˖-�rr�OJ!�۷o�˟�W_}��Ã�ݤ��3��UI�\��  ȇ��SN9�Q�w��-���̞� �=���^����;76l�j �R���R�=W��z�S�N�5k�P9ÿ�N�7�ׯ9�[�n�r����?�!���:ֹ���{   *U-�N���K_�7�x�hǨ	����A��葑Q������M^�c'��t
��K}��2^�������^�����R�cǎ���&L�-���D#�c��3@C���O�W�x2<F�{   @b��0����6L��I{͝B�gN���F���br��NZ�n+�xs#��yz,�<Y��U�J�M���j]��y^�=r���?�yQ������;��܃�cR��_o� mܴ�V�������<ꨳ����{   ���k��R'Ml�#ݗ޻p��(���XG�Ο.�����|{=������N���,U�x�F�MJ�>�rU����{���ɓZ��-��̢`0�q��zZ��L������6���-�
/kZ��   
�,Şs��ϟ���/��a�\mm����B:d�^d'�y��!�e+ߡG�|�zz	����:U�3z����¨~!	��/���.�%�wg�;�!X��,ze�:z��ר`�   �bR�b�ᇋK�:?��Ϭ\�R1c�D��'��	M����=�i�^��O�H+�|�@v�Boɼ���Dz�X/�NJ�&���=�ޟ̜�N��~'�5�����Esi������������  �/e)�~e��3�d�v�+������<��u�R1��&�fr�i{^�Gg�T�����	�7�m��B��@��wp��I'�?���\il��ϝ�z豗��^����   J��#����?���	��G���� =���	$q�z'�g�7����V��|k$�� %�ox'��?�޹����_ԟ#7|��%
i���"   �k �0w�d:�ă�*�*G}p�o��u��R�tYu��XG���$���D�zPgL��o�	����5�S.���z�����p��������'>�d�~&<0�+�p�   �K ��?��CD.�v��n�������k���z#jAs�����'�.��RKO������[;i��nI�Qy+dO]��t�Ǿ�SO<����2@�%sr�(=?0��s��D�#����T�tZip��S?~Hփ�c��#[��~yphtYdll�A��X�~^]]x��I-����ej��}���j9�:{	   �
�}��p쁢�]&�n�ݳ�������nL��>s��ӧ�ݼ��i���<�O��~���'(��Rx�+���^��DN����q���92�^?^N�^&b_�pjW��Ħ͝]����������;��cN�9}��f�w�ۏ'�����[�|�d��  �<|+�'�p-^��q�ܹs�u�Q4c��m۶m��o����'��A�ɞxr�e+߹�׷<�oٴy�]��o�f��>���-�sYL \�+�,Y<�^|y5��h}���m��h=7���Gc�2	����J;{�զ�16��Vn��M��i����/vs�W����-��p��J^��N��3�^[��    /��v�a��<��p�bqb��՞����_��,��ʚKn��krm�7�}�{�9�C�\r�^j��u���a��K���ql����� ~;l�QC�}4&�AY!G��\{T�)=:bA��#�zeٺs3]es�o{�g���/�������_ ��T   ���b�w�Nn�t��lݭ�H����~�����K��z����1���׫s ^�Yf��7��i&+��R�f�� t�pz^��{���;�3gΤ���7ߤe˖Q%0{�$q���Y��l���z��w���3C����{]�6��g��{ϩ�j�   
b�'����v������>����:746~������A�}��v����&�?eI�h̾3!�B��W'���(�1o�<�馛��8W��W������ݾz��7o�ݟ/(�8�����45������ÿ�{   ^ �ϓt����uK��:��������676�9�^s�Q(�H�8j�>U��L���T�>��8^����b���q�J�K\���і�]���X�v�<uάIk�k��]����  �0 �y�%.;�[\�oܴs���>��Wǻ�ާ�M����}fⴝ�~��vZ���fL�H����l�P%7[y����,\�y@�9�C�gϦl�2e�؟�N���m�A�w�}�����Hm����7lܹ�?<�^����n�䎕��=}������2��;   �o���[n�|�q�GAg�qF��?����c�9>�'��
�#���vu��/yLw��-��Cܶs�n���W�y3a�f��7I�ʱ�Ē,�R�/_N_�җ2>�����.]J�����o::�����1�������m;��B�  �o�~͚5bq­��;３��G��1<y��c��l�m4:�f�����x��x{Z�EqJF�������{}̡H�vJ#���	   (ߊ���K�i���1������{�XsS�cy���̓���O�1Q��¨��n�3�zjVz}LN�;쀽��Z�y)jk�U  �p��$�w��t��	�v�#���i��gFFFr�_͸�NϷ�r�\g`��2#r�4jtt�|��G��q��H4&���	�  @��I�F�\���L�'vw���m��qˏ���S5��������������"2�fbFٸR�;3�}HT)1(>x6 ��|AI�ɻ붚�����3��;���1���5�=��Q   
b���z�1�}�؟z�3���g���"� �A#Rh���9ӻ):f�ҕ\R0^U0^^�txj@��F����)䞋�#��td������t �ڷ�z��Cܯ���"  �*b�;w����������m^�����t�wu�Q5b�8��a�}���� =[{B�A#1���G/�7��(�:���p�8oPvv���m���rA��}}}�7�mߕ�   �l������b�`�9�}��C�>f����m߼���='��#�f\��7M�*_�5��� ��r/��r�B��sgx2+���Ɩm]�ΜƔ��#�>f�Ė��۾�.  x@Y�����7:��S֯]�v\��3S���N�;g����I-�g~�#?��w�~ǋ�}N�3��u�޾Aڱ������'����]��,=(��p��6���#�>�s�.䥘y6W�~�m���+頃�n�����������S'8n�:����~������ϼ8��>}�f͜�ᶝ� t�x7�  ��,Şg�䥔�|�]W�g�ϛ������=�<����|��Ť��@�J<+�|�1�Z��qJD�)�3���	��o���F�I)3��h=9H��/��KO��K�ÿ3nb���c�U'�x�M>�|A92��ߺ��N��t?o>   ��R������G�\�ZfrB[S��)S^��
�s�1�̓E��>5k��t���l=�8��'�ݒ{� +�L�O&�F����,�ȓ/_^[�����{�m·ɓZ���3�������L|�� �m�����   ��<��8//[G�?p��>{�1y��'�8��K~���������=��f�n�5�Ѧ-ȯׅ�-�L����n�|��yV{Zꍡow���	(!���i�����3޴��q�'^ڼsա<A\.�sy��-'>������U�h�N��  ��}<���iqLj��9�i�56�njkj�ԝ����l��짎Y8c����uf�ۏ�����N�)�M���ےےcfS#�y�%Pj���JZ��,�A�̂}f��T������w���ٴ{��:h�g��tLM�_4�'�]N   �W@���=�������oƴ�mS'��e򤦕;vv�t�}���Sz�>}��-��Ο7�p�('�����Zzw3��nXUr�F��'��=Qk��O�AO����9?���7{ƤI3�N�ۄ�O��kW��~��'�v��s�}҄	Mϟ7��pؽf���W���   xľ@���U���i4o�)i���>{MOl���o�-߽��kd8�m��XMm����~��p�����~�Uv�0��ט��m�l3����8��y��7���i�����DZ�]����������ݱ���pxBkkÄ֖��ޝ�EU�a �eSVEA�}�J3�4�3KTDDMm_-Ss-�4�J��TD����45-�ܗ�}c�E@����=8��02w`fx��H�w@��s��:�{��x��   9{=q9L�փ4ilr����8:�Y*^���U�9�]_�w(77�@7e��~\9���U���ؤ����uq����89�[*^*|�r{Z�~��+��  @-{	�B�u��ф�^:�����Υ�Q����3���������H���ˣ��l������Y������n���+��n߹G   RC����^��ƌx��x��9�����?̪.w�_��c+{��`k
�9�T����i���,>|8��ݛ6l�@��|��|�[]�9RogR�"��T   ��`/!���j�.طun�'i <�&m�v��g�9�vGM��Jd0��¾��r��Y
�?�E��wt��]����\����w�mIz��gc��G)''�   �^����^�u�?*~��3��'ﺵ�:w�ر���w�/.����3�-;�^���`�p����ax�~�'����zKЁ?۹y����t���T;�����]�E$�u[[[  (���q���ѣG����z�'&.��\����yѣ�Pc?O��,����n$�ѓ��s1TX�G��O�Nu��!c����u�xɭR�}eA�7���{�.^�(����m�7�R�&��S{_j��q�ZU�s�����B|���*�,�/&  ��T�`��_��ό�X��^~�e��=�:~������ɧ�y�;��S�/lk1k���/:e��fPl\*]��H���.T�2e
�=�$����3r��bd�Ku����E�h�a�z���N����i͚54~�xI�=�q�S�/��6���I�]��͙��ׯ��0sy���J��Ч�UE��E�R�P�l�2�֭[�c�r� ����~�ڵԥK�ܹs��s���/���_�}��I�\��F*!!!j�-]��n޼I���?�yo�G���+��G����L͚5#oo�R��p�n�:q��ʕ+�=��={>V�TkkkZ�d	��ѣ�1�|�  ��j��ǋ/�(B�j��_��~����*���+4i�$��>��3Z�z5�]����{Ӵ�=B���`��;�Uý���x���2YZZRhh(��ի̱���6m�ٳ�   J�����s�饗�צ�ʕ+髯�"c�� �����7������=���>I6��7��\�=���������S���۷  ��j�9�{.��u�p��#0v��>7�}<Ճ�M�'���[����\��z^ ���?  �:&�˜�}pp0���;j����ѢE��T�q�>��Q-T�{k㟹W�� �Ws	������W깳�|@۶m#   M�K0�pϻ����j�������8���ɴ�=�����:�~Ĉe�q��7om޼�   �A�Wa��~ذa4{�lT}�����:}!�b�ɯ�5���|:vV�6��;S��=&F�Y���?�����	  �<�j�b�:t(͝;Wm�߲e�8��F9Uű�}>�˨C=�oM_��W�$QzFA�3�p��oj�c�7����$   ] �k��[E�Z��ڶm[��{��.�&V��\��U�3���/f��m�c
�,�YԲ���f�6�b�'�<'Q�M����)�����������o��l+}���[4a���x-/t  ������◮��{ClbU�����Յ�;vЬY�L6Ի8Y��<���i�z�G�~�\/zi6�}U�pϋ����j����B=�1�P  ��<s�e,<�meU���g�n���t�ΝJ��x6��_��b��p��y�����Ǎ}���F������ˊp�Jp������?/s�g�����U���k׮��8s挸S  ���Q�n]��]]x�m�y�[U�z��� :i�������������޽{dJ\]�~���Y7e"�+���f>�7nܘ����ĉ^KaccC���t��y2�Z�w��IMM�)S�T�ݬ������Tպuk1�0g����  U�^��z\���5����ě���Y��F5�w�ؑ���Kz�L&�{�Y)°'5�cڡ^�ICZ5ߋ^��D�ws��gϞ�l�2q�[�Y��B��0���/�@�2.Sƥs< �Y�f�c< ~�������T��/_.�]�>U=�����wS��  ��^???�����ӳ̱������ɓdxӚ��\ѣ��@I:tuƓ&M��;��r�]e����ǲQ}�V��E���'����|ă?^��`��RՃ֊z�'D�:��Q��9�p666���	ݿ_,�U5d�qe�ԩ���O   �1�%��͛�P_�V�2����E�?}�4��;wRNN����0PR˖-��ó���#/wK��/��i�?����{qV"�ܖ&�;;;� koo/�޳g�^.���K� �ˋKϞ=K��W�^�dɒ2� �.8'N���D2&|W�g�����wx�ś�q�  �6晢����\��G��r�K�.�1��<����e���gv�D�?c����a%Bo]���q�6�-3������K�ũ��cJJ
͜9S�{��1c����������ƍd
('�w���˗���֭[d�x@��}�=T݋�;_�݇7�xCܙ  ����N�:�ʕ+����-|�r����_��wUK�5k&z{s�7��Ӡ��(S�p5�����W�qR}�ʙ�[i������O�>�o�)l|ׇg�y��ڵk�;=�G�&c�JÇ]�Ե}�<So�w�����ğ\W��u���C�y��p  � �?н{w�����\.K���#S�7����nԨQ��1^;�5�\g���LU��I����y~���^�R�|�z�4q��~�Z�s��	J���(Œʵk�D�E���������ȑ#ŝu��رc��K/�=)L�{�s�n���F�`^��0   U�TT��=�����\��OJJ"Sr��Q�<y�(�P�ѨQ#�y澪�--*^:Ru�^S���~� _� @WV���D9`���Jm˖-"�3ueiƂ��-<e�����8Քl޼Y������Ҳ�1�σ.n�ij_  ^���R���;wN�T޾}�L�������W_}E��5lؐ���)$$����ɜ����o�I���L��cK�y�½�D������\�Ã��|�j�L<������ӛo�i�e+��g�C��M\2�״)�� ��Q��}߾}飏>R{����/Nc��-���;<������y��̾{�.�M�^�Kה�e�}Lq����|[]�
��|�bj^\��鳳��}<w`�au�M���P�{;pi��w���_ğ��=���R���`  P�����Z������e6���W�{ղ
�������P_&���>�_-��K��?L&/����$6�l�K7���>其��tc�|���w߉���eS'�<@Y�hQ�RA��  PR���p].� C.N���!�dgkM�����G�Yt7C��V���nذ�̂ZsT&��K���FN�ºL��_���)O"+5s/3�j�b�+{�0ȥ ��k�9����S5kؒ�S�U\�\����~��ާ�{��	��]�v�u��  �6�*8�K�k(�|������wo��!6>��\O�3��ҝti�\�pA�ds�rsSj^M�/���%:T�eF�Ɋ�pJ|1�/{pn#	��6bR��I�&������|nc���d���	�5�����ȓx�*�_[����Υ�8��#�@�;  ��ހ<ݝ�ɮͩeso�R�n�� r��~����I���z�q�7&��d�/,���*V~̃�.¼�(�[XȊ�s�p�<U�֫.�V�7�R>�K�x�Ey�W܍��ё���^��G��Լi=�%{���l�i�:����m��围��sb�  P��Km��lM���U����e��/�/ޤm;�ѝt��S�Lm=�K�������D�/I�\0++
��x@��5�%?���������um���K��wlx݅6<��B��p�M�>�]�������g��vҠ�v   �^b��h�3��\�4kZ�����mG���X��/��R�^�`�^�9��v��)��kx���BM�7�֗��w���b5��J0`@���cǎT�6����=���IvNQ��ȋ���o1�  `(�j�����߶X��vԳ]鏃���=��+9[/ޖ�K�z���.T^�������5�E3�������r�����k�9�3ދ��~S������EkĒƌCG���{��=���7͛7O��_sDDU<C?̿�Ne7���tW\�'��C  ��%Ү�=;�Q��/t��h��۾4+5[O����`/+��/^fˡ�̾+�Ǉ,G
������/�C�
���N7nnn��ٳg�Y���������C����x�b��СC��yyy��իETƏۺu+��.�hp�N������7��   RC�� w�xfP�J�I��DK���M��_��Nm���g.נ���{��R��%>���.5Өc�po!*(�m��½ʷ�2�rx7d�_~�����E�_���{�]�8��=�T�s�I�\��%<��7n�K�.�����'�?�ڵkŋ��:���;V���_�����~O�s�   ��`�''G{
�{�M������G�����\V��|+����u;ww��^�.΢���������t3�6A���*a=�=���u��ϣ�»da)+Ȫ��^.��0�O�F�i܍5&&F<�g��cx ��?$$D����{1[o�j�Ԥa�u��@rJ���[�gg�+((����(����������������Cy���CvT\�i����p  `<L"؇��QӦM˼�Krss�*�?�Qt�(OL|JJḼW£vGi{ܘQ�����޷�G#m��?J+��ir	�\��M�[�+k蕳��R����&�tO��ƛqoze��:�w�ĉ)--M�p�����5�g�g�Q�c荞��Ё�E���܈MI���:iæ]?i{\��~}�븬i���[�τ��=�߅V���  P9L"�s�=��!r	N�G�i}LAA!�r_�j�/u9g����oHP�)m[�,�ao�1xy8S�����1��B�b�?gF6[�ă��ӧS\\�h{�NTT�8�t��U1b��a��G�9VVVt��=:~�8͚5�������bw�����+��w���o�r��;w)��?>���Z7�ikk���~=Wj�ʇN��N   R0�`o�zuo��x~~=~�����x�s�۰�#�:Ѧ��N����|x��'��H��_M=a��V˖-{����Ƞ�Ru���ߜ�<��cWƆG����_����cF�9ޡ���54�{=тN���`!7  �~�+��W-jX�]�q�'���yEB�RX�o�C����ܾ�:++�ٞ��lV_��Fqw����h�0�C��(��:�.��]��n̯H�W
��������4�T��ڎ�ԯ.��O   �B�����j=~�z�կ�mM��Y�qWXM{��6�|���n��`/!�2��3�Pofڕs�^����ڍ;f��<߄��ËCG�x��1M��r{  ��}5���x��b�neK�\i�����Ntt��Tw��Ǔ��,E�Ou&{���(���0^�<^����y��_��E���MPS�:��������z�[I�#��w���$�������8  �/�
����\�4��O���~@��۴i_��.�Z6��M�q.��x�n$SuU��U�鑑D����E�����(&ɵ��hS�Il|�刈��H�|[����r>ݼ�w[uǹ+O�Z��F   �@�� O7g��S��jm�W��d~������nN�2ؗ
�*��l��X�cQb���E�91so�ݝ�OI��V��L�s�k��j:���`  z�R���:^���Mm��ɣ�R?gLB�����u��ծ�@PD����+Kˢ�e��[���ԗ��q���xAAA��ϙ�%�`����]p� ���ls,��i�;��nm��?p��|v�lh#˵8-�s�۷/����N��j���l���+Z�*+ڨJ��z*�-d%f�eŵ���L�����\�~?/�_��s��]ɝ��i�ko��&Y   ���Ԍ��y���pl|�ӵ�	�YZhNs<Sl[+)�ϛ�_�����x��RW�Sj��a��`�^9C/f�e�R���>�����M!!!b�;w��bA7�Z��������d;����BE���  #���̺� ����.�$KO�$�,7Os�x�wݛ+^�|־����i��\��)T���>�wi�����>�r�غ9��o�^�_�/9[_��px��M�6Q�ڵ�ۃ�)S�����	ʗ��Z������ذa��Vz��aU��������G   �*�'0f�����e!A�\��wTP��L5�w?[�q��N$q������Fc�̼��s2w����֗-gQK���|�hWYy�c���+�,�N�����~��݋C��СC�ut�~���<�����=��kڤ��s���/  H�T���wλ�_A��?�c��	�KI��zܱ���k�|���S�OM��9U'���<�k�|?�O^��¸\%��2[�\�@_���߅�P͠��
�t�Rε��\s"I��nV�����  ��Ri�W����G����XLlR�c'.��t+]l��.����c�g��ܹ$�mwW��ڎ�'ܦ�䬽j�grR������f�e�ߧ.�WE��믿(--�Ԭ��m�t��x[,��аV��ݹ�������_��hu	  �+3�8#)2�����b��h�u�&�w���K%߆j���:�;9p!�/Zg�u<��s>�ݽ5O�{�RR�h	������<ůk����Y�;w���ѣ��Y��w烈~�|�����'��w]�m~�<\�?=}��_C�x�	���_��M��䔻t7#�   ������1��^���q�?_�4����$¤�9�1�3ű���I��_�y���[�4l�J�%E�=G����^*��ڷ�-�Xc肣*&&��͛GP1�����Ycϙ�������Y�[a��k4��T��˿�c	  @
s��/���?��?��ݳ:��\,|�=Y��^G�\��zg��ѣG}�A_�����zuk�������V2З|[�>]6��������T�Vde����n��f��=��SR״��a/OͻO��gn  �������y�MK�6}{w�s�a��de�ґW�k������+������S6o�-�a��5��7�m٬~m��x%�������}E��K_N)u�v�Ӹ�g��������y۶c���|���k��4��R����� �T��q��foZ���A�?��z�b��<G�6Һ�kc_O_���q���l���.��l�Gs3<�o���K��x�o��!�Nu��"�g��R��>ﺱG��m��`�b�2j���;t9�QO�hP���n���_P@{���   �Rn��Q�]�^?TH����FX���"M���lڵ�4��Q���V����VO�ZWn��]��vm��U�i���
rws~��_����Dy��e���n8a���S���ԯW���W������vw��i�>;{1u��c�J�(5|8Y�Z�q���z��^�5���t����   ��S����"ׇ�>�֒ϣD�G(�ẉ_j֤���qk���u�/K�g5Zܥ]��쬼t�\^`ooS�������^�}���ݧ *��C��|zj}o.լI�f�WW�k��|P�G2�����= {;g'{G�������i�w�Y  ��λڜ��3�Ec�N�#�\�Q�;ҒY�n�����]h��ri�w?�M�����:}L{Y��N�W�*�����b��'.g��z�&��C��u���5�,/�~�=���R   )���Ν[�q゠.��|%��C�W�m�=�y!�M�h����Z���:�w?��"�S�m�ة�Z\>ujM�ε8�Z�ZZZҫ��J�jբ�?��RRR*t��M�����8G^^U|M��;!��8�4�s��0�sq�  ��C�C?z�����x������j܈ѫE�Y�_ث�vSP@wj��F���3£��3ꢱxu9;XP��T�$����{�j�g̘A#F��T���̙3�C����IӦM3�;b����{��o]�Zd��zŠ�k�  ᡂ=�q:r}����o�x�Fʼ���g��7�Rߞ��k�G4nY_���A?�8F99�5�ZP(�ٟ�����zt�A��ݙ���vs��g���g����
�k�ڵԺuk1k���F�1U'E��ߨ�v�h��$�h�5��?u���<����  硃=<}cdxh�q�_\��Q�
E


Ţ�Sgch�S���#19���v��\K"s��/�i�ܢ��q�';�o��e�=�pe
I5ޱcGz��7��^�x1;v���۳g����裏(88�RSSi���T���� ~��4�o{���'�)�ߓt=�  Z��=K���z�&����>����\<��s�{�n�|��^�IH�-f�}�Q�~���Z�e�ă�KW��ɫt�R�d��P�z������E�h���D'��{ݧ>�.�;88�u+��K�СC�a�����YZ�jEAAA��o�p�u�V2'N�S�N��Y_ܵ�Ks�zR��~Լi=�ߵnMo���p9����L���_�haaA���:  ����~���y�k�W��q�uN��D�nݺ�q�F�2e
���z��Fl�x��������N�NT˥�X[�r���|J��%j�o�ݢ1)��-��J<�;~�x2f���8�>��I];ؓ�8x"�f,N&)�����T�N�znn./nW �����?N~~~4g��s��ݻ��]�6m(**�^|�E�tI���\O/66V�Pq�6�v%w7'rv�)���:|��͸O�R3(6.��ݸ�x�4%svvv�p�B�ӧ  ������{71r���A#��MLJ�NH��v�2���%[[��9�gCW�X!fD9�K�kk����KjlmmEiE�~��� $��T��.L��3<�Sk���ʦ)���%���f����nWh(,]���/_.����KF�=J�z�*Sσ��|����=_�"�_�� ^*����X�9x�   ��W�g#�f�Z:�����-��l	g�m߾}4v�X��O�O>��>}:5nܘBCCM�������ڸ[.��r��L�j���#�7�'ӧ3=�CK;2U'���;�(7�pkP8����K~^}j�+CXX%%%�k��%լYS�O?�����2E���_|!� ����҇~H   %��Y��i���t3����~��&�2���Q�h�ʕ◩*�K�_�>���[t���l�ޠA6l����-[D[Dc�p��$�t�'�oaz��̅z]��g��bHNN�2R����3y�k�v��A7o�!^����Y�8 ������wL������V�o�   ��$��d2yt��	mZ���ݣc�ݿ�l����x
��={�,s��###EI�����صk�N�����9fJ��C�[�ɴ\�[6�%Sq�j.��a2��2|x��������-ZD�Ν+���s�wr���1;}��|��{�f��������b��)̇J�g�&�2�xp�w��  PG�`��fn
6dP��1�IΗ�đ)�w����k�� �|||(""Bt�8r�����ӂ4w۶m#S�y��^��D��xR����/�ȥ��$������Iי�I�&ѣ�>J/��2���+:}�����>س��D3f�����8��k�v�#^+��~y�@]����t�};~�8  h"Y�g��N��)l��qcn]�l�����!�K8_�rE��l%��!�믿3j?��7S�NU�\�.�^;�N�"ܿ���z����?��J�]@S$Qz����ڼys�'���ʘ�pT� ��y�=a2�y`��@y�����dLx��������/��ݸq�   ��<%�;����'����lE4���N���Ѣv���q���������e˖z���R�Νi���j�q��J�9���Q��I�����ԨQ~���U����"���P����j��̗,YB			��{��siڪU�諯�2�NP��N�:�=ƃ^��3�   �1���˹�[4�j7�=���n��?���F���3ψ�1S�3����*���rtt,�1M�4)�<;���!�W���quS�i�&1�偹��rt-E�j?����;ȝ�   ta�`?w�����فݻ�=�����d�xF��}��ggԌٯ��JӦM�������.K�<yR�c�u�V�m��{S������4b��H\Sg(c�\�Γ
rSj1  U�`�s�"�<;����o޲��K&S�3ݼU��Xc��_�6��I�h��j����a�(;;��������]�,��@��ې���׹~�qM:/��ڷoO��g�g͚E?��  <,��D;�D��oL7䫏o�{����/[�ٽx�w�0e����EЋ��"0_<p�և���N����)�̳�%�m�V�G~Q7�2d�ظ�q-:?�Tݾ}�ƍ'�l�˘�$��bl�{ �t��H@�U��]���r�*,4�d@��%��v�ڕ����l,�7n�ڻwo�ʑ�9R�a��?�P���}��Q��<��V�ŃA�����S�����O�<�仱(���={������/ܵ��ի  PQ��;0+?�fM�����N��z�Lٮ]��@U� ��'x�Z�j� �}ܹW;���N�^^^�>����r�=��<���5�C>/W��o�k]6�2��  `�*%؏77;:�g��r,&6���s� S���Lo���h��]l�Ｆi ,]�T<��O?��ݻ��s�W p�ȷ�~%!   &��v�	�^̦��#ǌz��E�6Y����"��8|Ϝ9S��hZ��w�^�T%f��C�{�����nfƏ�3g��c�mj  ��J��sԘ���CgO?�CE����| �l۶M얬�E�'J���뼨�?�K�.bq-w�ᅦǏ{8   ���`φM�ް�C`@�aa� �"�𼘔_   �<Tz���d��Wҹ�#ͯ]��|��S     ���`φ>?5�ۍ���p|B�㕫�     W%��=7z�����'M;h��K"(==�     �b�,س��3"#ׇ>��X�ח�����B    ��W���y�ϙ"#��C=����     <�*��z�͏��лg�c7b�?y�     ��Ty�g��3���B�����̈́T�ĤT     �E�gc��Z�Τ�C>]�4���s     tc4�����Y����>=��?�\N     ��
������6�|���ݹ���G     �gt�> ��Mk���h\�-��_'     ���=5n��MBC���a��Դ�     �e�g���o�\?��qCf.�,����	     �3�`��]ɝ��Ͻ�sC{ش�7     ��:�ϝ;�p����>����$߿�!     (˨�==z�����<�����j܈I$     (��=<�TT���Ϗ��x�Fʼ�E     ���lĘ"��w<��_}G��ؽ
    @�d�=K���Z�Ʋ���v���     EL*�O�<9���?ի˱���:'O_"     0�`Ϟ�~B����F�ۙ��f���J     ՝�{62h�����O7x�e���K     ՙI{6<h�'�B;������~"9��   @5f��^&�ɣ�g�oӪq�^Ovh�g�q    ��L6س������B����#�q�N���    @ud����;�⦰���ܺpi��Nz&    T7&�٨��~�\���!��Y�"���    �:1�`�,�Ok�@���!O�ۼe/    T'f�
����x����ؤ����K     Յ�{6l��Ԉ��#G�/>!�66.�     ��
�,0x��Qa�oL��E䷻I^��    `��m�"��{6b��/�����I�t'     s'��a�?���    IEND�B`�PK
     t$v[F���9  �9  /   images/915d9337-ea3e-4fec-8caa-7acd53f715e1.png�PNG

   IHDR   d   �   ,�*�   	pHYs  \F  \F�CA  9�IDATx��]|TU�?o�d���B�RD�4�b�]�k]e-k�om����mVY]�  *-� Az��������̝�Lf�	�Ā{�Ef����#|2�z���ԡCkJo�r��m��N�N!����I���R|����ޛ��7��YCzS���;��|���'J�����H��A��xs���;���o0`����%�x� B�嬡�6)������������].�X,��jyr ����J�.ϫ� ��S{hm�����36�R�w<_��Qs�K̃|_����p2kS�9�;����P���t�O���;_=�w|�\�6��&O�L�ƍ���2�$�������^z��v{���^��5����������n�;�xI��a��z=������$�b�O�Bqqq���?��ٳ�X��ЫW/����C�ѱcǨ_�~<�v�"��ɟ�>�:u���r:~�8_��	�hC�n���?��7�ֵ]4i�훶���r���_~9�y�4m�cd�+Ծ]*��Vѡ����.��~��}�Y�o@D�Rt��í�[�A|�cD @+&r���9�DL�����ٓ'~РAt��AZ�jU��������g��ى	:t�P �%�=������qM�?v�Xߘ1cxq	����ڽ{7�o2��[�fQqqqDH�M���;a8��H���ת�l�&qLs�Υ��:��O�N�1Z���1��丵B�w]�|K�'�Φ!C�P�6mx�h?���6�L6�G�� d��W#���$ھ�N+�*�Sf;��̤_~��'?5550h 	/�������1���qg3�u�����ϧ+����Ow�_|AM&iժS������A�� �ĉ���@1w��ѣG�#A��w�LpF���������h��j�F&L`6a�Z�-���1��]F�c�]�d�k���ge��}	UUU5o(dDz�N��X�^r8�B���hp

�ɨPj���&/WRR�+,0XI���RjJ<�է,�d�h4�s�f����{y�Ϲ�.�@%���ԱcG3&�cbbx1��O8�� ,X@�&M���Fh}����WڡC�x���Ly�����W��ŋ馛nb�-&�|gi���^�^Wn4�j���bA �N��I�K���e�Q��x1�!P���h���L%x6^<)�9�]jˬ6�^��Iq��f���ur"�a��=�����g�M{�졽{������e�<P	۶m�a8."�5v�Yo:\pV,���CVV�s��&n!S6m�Gݻd�c6f*e���v'J�1��uE�~@��������j>����=y����c��-H�gӖ�YJ��;H�,��*&��/���A!�.�����w����y�6|�]w$��mN�ۿ�|������!X���[�x��������rZ�n�8W#�%�xy��_Q2��LYBU[-�Ҳz���z���Ç�̙3Y8l!11Q�}��:�Wt�`_���}�6l�C}����yU�>��fJII�X������v�Xqn 2�`��7�D���*mں�6�`���!Pw��AG����[wکow#O�Ɉ�}Ǵ�{Q���v��k�����E]��5Xؚ5kz~^^���S�~����a����o׎n��V<�Hۻ����s��)�� �`����+ڳ{��C� #��	�2q�Dz��H�+��P:���sS�\����3o
����g[�P���@��-��T@��X�{<
O8�Zi��W5��Z޷�~+�}�i��? ��|�7o_�\6J}���"!ན�)��+/� ���[����������9�5WЎ]���'=�����O�
��;/��b�����U�ӧ����L�7Y	l,���'��!y�z���Yh��ўR�b)w>}�駔��F��v�<�.��%��Ӓ��2&H�r������׵kWz��Q�i�C���b�ݞ�����oW�J��� �I�*���)Ե���v<����r�U	�y��䖖�ȑ#Y��z�[�n���}��K�ѥ��w�V��.+�^����s��zwHY!_�)�{CA*iY�?��{�b��d�J�b�F��]�θ�.��v�w۴f��TWc��I!� 1�؝&r��L�r�,�`wD1&���k�e�_)��_��pR�D6�k���\��!A%7�>����?��k[:4�[!�hU�G"��4�C��j����v�ø׿(a��x�'}ʵ�)~����=�~��B[�lawWþ}�B
a�x���8�no�G�/�N[������m�B&G�i$f]B�\�au���Ua �:L�!m
���	l�8��l��B�R�@)� �ڷo���J��$Rv��w6��o3bh�����.��MY�~7�K9��!$c �b:��:�oG?���JK+�t�� ��},t�Ff:�"׳�Y`t������A�n�'�A��Bp[b,4����kϑ��{o>ӨQ#��p��TA!^��J���U)}J@ȇ~(�?Q�Ν�&T��k�V�:�fv��?���Z��h{���w6����!PÜE�wt蘓��u0Ҁ0���j����e�~�K�/_N��Ӵl�2���է-9��,�S� �tIIq?��W��2"�"_���g����ǋU���`4�^�:���r��;�6�h�y�>��Z��=f�.c;$�$&�W:�3�G�	v��~`c�{��N$<���t�ȑ*���_{����ya�����O5O�˂��R�lx�
��PB��ܶ�*�V���qq4wI�����P����B��W<Tp8�֮][����z:��V��䙫&��y�
)2�R����Jۧ�@��돂@��CQ�ֽ���1���NA1fK� � �b���o� TK]YY=���U_�}~�%W?:����H��R�u�]ד����^�O���)��b�|��� ��$�ӯ���Ks�-�iO�[�`�W\p�C@ʤF!��CnMU/ ���bm(5���-�Z�r��'��]�4��gi�ܥ����m]��˓Ͻ䁓G��V�#P_5��?�)���^R<!'�����L�F�?|���[F�?�u���&���ϟ	�\�p�(T�o�2�����dI�9�uTt�E��Fκ�������~�uӘR�|���>����%o^9z�ݟh RpN�ЬV����5�BZ�%�Vo!<�N�q��V��B�	5\'J��������'{�ra�H�����0"��$��8��=6�͊3W�$�R�U~�P˗%)���w�`��yƕCG�1b�`�;d�������`��v�7�B�s\�+�N�#[ۈU�u_��͛ӚV�xS�)����-+�+��q�@�Eu��p�dP���X2�r�;�DN��<.;�����R�d��n��U��1���{����E���o�$R>�/�r��lY�]5���ˏ�V�F�|^����cȥ1P^�P��&�ٲ���8�*����ĳv��q����;w�{�$R������u霑#�1�޻��<>K�m�Gns�`W?����"E �ů�����p��ɨ����� �5�=N�;���V��Б�}��؞'�-���UGH��[�	�4�ӧ{reB�o��z \#�V�!dp���q5~d�B���@"��}�S�W$!��[FJT�yDb��+iH�1�@���yI/>�]XF��T�N���ֲ�����Lh\�B@�:� ����%�pu%�k�Sm�b.{9�1/S|XW]u�f!�!ZȐY-�2�4�:B�X$��?��C�#�����LD�
�ѿNʋ���m)�rXX|�A�d�a⑟E�+RI�yK�B47hq�Q�_����}�b�_=��)Ox��C�r����B�.�7'gU�G!`92�3�o���P� � @&l#4|* ����RyYQt��ONN�J#$HD �yW��C���`+��"���oC����(	� ))�	�C�D� ^֨�2F�����ZEj4*�E��b+�J�/|\@޺u��|T#���.�R��͑"Tf����I�8����%j��!��<HX �9^�m��4l�0Nj��SWf:<�����$�F$��HY�v��!�`�*�IG��W��`a�8���٣�����&eo�D볲��!D�Y�#s��-��09�f�d##/J���+V��B���??@}�S��������(;;;0�`��������'��(����z�,�Id���E��V)���V^FW^z)y�8�ʲ��v�y��F=�p|��
+erK�,��wL���R���; ��(�jR��#�֬Y<ѐo�_=˴p���K.���Xdi�GL���|_�,�(:�_Sb~�RL�Y����!�._ٌ`1HxC-7 �L����8��*B�{Af�� �{}��G<q'S���aL�g&��{�;V+��X��,2�J!���S�$��jYxQ\��]�mۖ�/�*y��z�#E�0L�"'�VncTe�\P
X�,����������)�v&���Цd�	 2��,���z�|�0��� *I�s�	��q/����V͛YU���C��F�jY����{�Z׃l��`Y���"y=V6���#b*	85
�AD���4pȆ\���L�� (L�����_��A:�����U
��!�!�0�ËJ5���c��Q��$9|��!��o7�t3�2z�����`�P�Q�d�J��P);�8~ٺ�>��	��R
j'�J�]���Æsi_EE99��Z�tOQAz�8�3ʧ?�#f �gZ2���܊8�C����r@^>�j]�8߁�t��y!�G	���3g��5�Nz�C�\��^��T%"Ҥn�z$V�y�'�9�脄�})�¦g�6P&khN���n̪�ލF\��zi���XP�F�p����M��ә}Mt��XBfV6:@`K��4sn)uH7����9�W��{��{h��et�@3]61�wNE����<Θ]Bǋ�ܔ ����Ȃ�(
��>��lNV@ +�	5]� �p���B��҅�
�&j"
e��f�7�hM��������U�0syB�t}��uN�pFO�k�����ZT�c7�L3��j���z&}5�:Z�j�g
H]�� �WYe�7�y�Λ0��R�XA(�������s�1�r

�)-=�������X���dUV�x�O�ts�5&|�����8>|��'Z^(�U|K���b��*����k8~�g#4�j��ۑ�'x��:?�����	�ӊ�q@+��,�Z�|<��f"�+�L�B�5U]*�W�c��)�`�q�59H]/ʈ��9�c�1����$�ǰ�c�s�$�1j~���pWX��/�Et�/��&}Y�A�*R���8$�ͽd=�Y��	�U �+��G���B��h�7�å��؇�@-#��E2�������װ�e��B��ؐQs����Q9�K�:n�d+�������8�4Ν�f
�����!�Y+�z����4JPCᦁ����{F�OR�p�x
��-��(�3���P�wt����b�}\��P��ֈ�z�h���P��?!�<Y���d��t������n��Z�u4<7n��_�-
�d�(e�G?�D[E[G�T�:�kuu�����-LɊ wJ�y��4fM�L8<]�0@��j|�`�r�5d2ǒUhX�.~wE���o�˾.��gE�e�d@���"���[(&��ý��	�~���|�dw8�cy\��&�-dbUe%�Ξ={��dj^�	�W���US�2�w�-�;�|Me��{�.���Cj�P�a�z+B�f�?��%����X,p�~q1�s�I-�;y������g�+.��bcL4��+h����RaTe�2[k�i�$�c#%�����x��-Y��d������ǡB�ڻ	�"d�~�#�e�ތ�8C��9�kD2�������8ʉ�~Z�gР���jel������'�"���ӛ�Bj�^L�SiO���ș��x�R�s�.�O����2����tP{��׋%�@��B�<��A�u��䊿C��%�x�ۙ��rbB�}r�9���_�뀌O?�4p�ψh��6��D��jס#ev�R��ɥH.��l�ѓE��l�������1�M��)VwT�~��h�������Ψ���=!t:a'����S���-_�o}�7r&L��Ƞ�;��.�&��X|�@��,���ԘEX�U�����
��z<r�	/�KY>���dS�o��715�%����:��`Ih������8�ٳC�QQأ+c�tL��:���$adpFC��&��1��St�� |�h��I)�Z!5�ז���78 �#�����dpL~�5	u�LAT�DU�DlFQjPz��	�~e%͚_JW_�N����do�a�?�=�.K�\�hA�;Ĉ'��렇_8N�]OS.M�u}�n;M}*�F6�]Hb^�qq�>+=��	�h�6`�,�/�lvG����q�BV��m4�@f���"�lay+C=zq�����
>���?��M��gҼE%�Z`��>�9.�/��_\A߯����&V;/��,Q����ŉr�5�!@��M�3k�����9�qLa����?�f��u�ӻ�޽�z$&Pv�&�5u�ؙ������C�z�����z@yEm��WoBM�!�C��Gi�ZQ��N
e��B,��hY��KC���8��A�sZ��cƌ����yw���[�F����4#��{��n��o���ڐ���Fx�����ģ-, y�HF �"�9J���K��pU�2��A��Y� �d4J�M4��ǰ�Offf����X&^`�JX�' /@�X��'����
[�Ȟ&��n跈|_4WFb@�������~,P$r�1��%r��J`쬀s�%Ly�E
͊��:�J� �i�E���F�λ�%bQ qBv ��C����u�V�i�R^���<l�g���lv
	œ%b��5�ѥK����y����mi��6�������l���o֛@6� ��uz�?��kI5
%f�.�CI�W׽�4\3|�(�C6E}a0`U�Ș1cO:��1�sƌ�Bl��w�#��������t��W��7��~�p�hq>z��ݛ|����$%NCZ��<��]��J�.�D=z���>������ɾ,^/���}D@X؂�B)�z �j(Vw����l�}�Nyx.jAP��FF��Ub�i���E �+�+�@��#�~�=����D���?Ε_X��H2�I��IoO�N��J�NZ�����x��:PN��]<�"n� os8�u��C�
]V�\x &���SO=��!��ܖ�q�d��� )V�>���wЉt|}���q�*J��AP�S�?O�۴�cyy�C&|z�v��n��.�!�(���"֮�jP�-��JIl�D��G�YG�?	��顸X�M���o��nddoڴ)$RŲ�A`�����%B�K�O�Ǟ��9l�e�-6�g6�-��Wd��I&��?�HXø|�1.U�-�1FP���U'
���R�x'l E M��f3���0r9:e��X#CՃ����Ř�PR�Z���|�d��P�h�.����W�EY`k}ړVS��%G�*��d�-��}0��ΑBn��|{Ne
!������Lv��k�L���/�mGF?4/i?!�j����)~x��x]Md�I�h�
��ӱy!BCk�`E&jZV��x��B�~��A+^�H4ǘ#ҪԈ	~F]Ȕa[���KSyY�
�F���PQ%~k#&��0P�	`��M +��{���$��E�8�@�0�v� �f-�|Z���}������˃a�����3f��%�J��T����Y�1I�����Z�);%�%ԥsV!!�Bir�=!�T5!˸{�9�%�ɖ�V$���xj#Q֪p%�X��c�v]�K�9�^Cv���;�!*1u���LՐI�l���A��U�[Bjr�#��7��bk�:UV�28������IF�@a����3;�ז��.�{��s�$�͋M�AƉ���wԹ�܌���E��e�H@<�-X��� yMz����zW����]�ԉ����ߺ41�D�[y�F�eW^I'��+:X��m�5�����Pi��
b ���5+B{+q0���3Iq�&��.s	�؆�d�	�0�#C	��Zv^��� �wNj��d	4Մ�����f��'�uA�C�EM��_Y�F�G|`S?�
@�)�п_�ڶ�Z��"�)�5�k�)�n*�QD�t�,J$T�b��gY����;f�_���oǱ����ۯ/���ճ�ԪWUV5Y'kL.�9c���:_{�%�#xR%k����W_���n�HP�Z��3��B�/�>AI�P��3
�Z~6�6�;Kȶ��.��zZ�pA�qG!b����Rz���ŋ�;(��J|ը>�t9��M�:ұ3Ti�B�zJ�"�ǎ�1b��@t��M-��k�%�d�ʀ,X�?����j���W�8n��F���,:��%�M%C���d���!(��<yN���h���\�����Ι=��c��Y�XI��=���W��+2>!��}Y�t���;X��U���-����}�tr����\V��@ T���t�M�.keoȦbw�8���7x�Գkws�9��P�k��F;�>T��Uj%r�ei2��M	���Y�/�����NB�`�^�� ���,ul��z���\8\"-��	,�)¨t���Bn�Xbد��*X���ȢO{ �չ�x9�&�B��^Mâq���ip�e���pxq�@Y�.A.$�\z�̢^|�E����tP
�G0<�.��@uP,pLvC��<�lAM!��]��"X�R]�D�7�/��#�
W��7Ae����4֍������r���S�2�G�	��'�,pb��EA�������G��r!5d'�F�e)�@M!��" � �#l��Mk��A��}�Tf/�s��4!X��޷҂n���U�{͙3�����?ƈP4؊l/	���|��qG��I�` �9��eoΦ�}���P�c=2� ��a 8#Q{r�� ��)`>`#��Q�eed����L�U�/7W���M(���yMG�^���>�h*�Vj���;�d�/��a��.�A�>�� ��A;�z< <�!Էc�O�T��p���ǆ#P��D���@~��7�	Ra���単	��'�;�]-41�������&�AT|Y.��*���$���õ|Yj�)�!�%ży}}���&�e�����駟x ��;�C���?�˟����>V��T\\Q�<: ��+�g �< _�NE
Q�e	��d��g��}Y���p��8�!5)n�$d*Tl�!�ٛiܸ��WJ��(�N*)-�ٟ/fѰ�v��$ �
����/I�tU�^��λ֫n��~�;��?����J�D\���YM	?�9d��۠U�i#���2�"�z^�zP�}��.$?4�dٲ����8�;��޿&@m���!�w	�v7
!��PS�� P�㪮R4�T�IJNb�����!�Ы�ɭ�ɔ�f���]h�/>�#�Ӏ�����L*Cj����h��m!��-g[�Y�D�SF�j,4ڗ%�&�2)@�t8�T^Q�Ã�r8SSG�Tf��ہ�u����`cN�� & ���o`�6�I�K|��䲁��<@]N��&T47�����B���+�����;����#@�Ipn,�@�M�{��c�@�A��B��`��T4p�(w 2#x�F�,��Y��sG��7�歿В%��:O]���}.'�4H��Klٺ����|
.��l2 ��f�DJ�}X�ֳ�AA�}Y`W�**=�IX�*�?6G:8B��,K�x��'Z����w�dܷ�=ڑ/�T$�H���?E_�lBXGF���I�va�\�*@�M�UQ����Yh(����@��a�3�(�u7_���[˿�����ܽ,�;v��	l��l��wbC!�������ڮ��V�{���K��man@�������lm�U��r���Z�!Q$��(<�joz�t� ���D:����pђ�7�OQdԮ�/��B���2|��b�ڬ�4Ҩԇ������[���&΁f���
Ë�,���E��F
2�����p��W���e�7<؏
���ܨ{Q4���@��P*Ԋ�Lܖ�79p�@���T�uP+I��e94�H����c2K ܣ�pd�c!�lx�;����4J`#2T�a�H9N�lB0�؛v��e2/K��~�jo`���&�a�{ե�+ j,����{6@RF�be���w���4B0AH^X�pa��`��*Wg�KA'��Ϫ�����<TC��E�Et�o������yY�����"�V�(2r�M����Y$�H�'�t`�NZ�[><4q�0Ҭ<�d_�%�7c�ԣ{F�իX��2ޢ�c~��0'r�6���!����o/�����Zu
���Pk��oO �Iŷ!����TC�
͂�f�����k!����\;�<�Z�{�N�dS��_�J�Ӝ�*�kS�	.���T�қ�� !�bb`�A��U���|�h��15����/�B���X�|t�
l�d�anRPX�N���3�?#�=�O��n4Y"���n�އ�#)�,� ��i�2�f�#�Mф4{{&5D��O�3�f��t����N�+0�p!�PI�jc�I��[��@��V'��&�В"��P�������b���
f��?�
pZ!DB}�-N;�H��}���$8�"�#���I�&E={>҈��B� �>��r�)�	��P��*��!���\ ��T0�,�7�M��x�Av��wA�G��Pz��Qj&cu5�i(HgjEyw#B�+)^�޲�-����e�eL�M��L���k΍���֊7/V�Q 鳥e�׷
�d��>X&�~Ԏ��x4�D�i��kD�6l������ J7	�|US�U�.�69B��w��:t0r�TWV����%���Oe�1���ۤ�v��C��,���D Bx�v8d�����[���#����ǡI"�� �c��̶⡂59=�E�E���S+oԐ���l/';`�pC���v|-�'W~(6�ܧ��v6�߮mF��G�Hb�H��u�Sד��.&��A�R[�q��wxF���A��سn�:j鹸�>�('��UA�ο���<�>q��g]��@@9<Z�x5�}��Չ �XP���!Э�%g6ԉ�w�5��{�5�8~8��ݩ���VO�/����aW5��<zY�?���s2�Ɛ�J�Y��������袋�qC����C]#"��9�����4jD��3��wK�.*,*k_�)��]I��.��T��c*��rZ���N��M���^�H��+EN�"�4�E��#A�_�rd +1!��"�@�=���F�@�zf�^�4k��%��K"�BH��j�2�,�?Fn$����
Z���Lz>��PZ �mD2^�'Z�����O6E�Cu4Q�YH�H�J�j!d�@Ɵ�}��=�z���d�E���B��R�7�V����.B����K#��;\�Ѵ�a����TR�� `r��2��������Yp�B�y�Q�c�K4��3��z/^�nщ �46�,4)G``��9q/�n�s��i��JV��J�����/�<��wY�UR\«_�\n���+������LFŗ�(=�����#t�ԗi��3�W��}2�h e ��&�L��c��h�b�B�2-�'(1Y ʤPr|5����w�ۛ���Hp����}�� �׷�}m#��s}�Y��!�E?v#cɲ��N��;���Vׂ�
�-�]ag�%g�hr��"c|��xٿ	�:m���X`R&E��:C��"ɢe���?V�tF�C���Oj�o���2Ae��:���s,"��l�ᾺXy`/�PO�ْM�%,\�%-5P%����DJ.W2���c����/2J���|ֵ��i��G�X�z65Z�!�Nv��ZG{=xP��B�ʓ�E���h�"f!�
\K� ��aWo좐�G�q�����M����`�"A�sj�k�����D㲒	��Ѐ/���M�:�8�ju@c���+�	5��X��\�MFK��g����u�q��������*Xu�7;x� ;���&�J�ݹ�4���h��/�}�� T޷�Ӫ�V2�t��{�rkV�lT�#��-\+�n��Fe]���ء3ڠ[��/��(m���S}����5�����{o�>㭷���u)ر!5UC��]�9�	d�ꩧ�V:*,v1k¶@6c+;u�{P�a�4��/���r$p̘1��o�-UV4tV�=98�VR���C�#Jְ�qFz2��UQޱ"�۷#�'�`ׇ�l<a�L�,�bL�څN%�+�T�*4jH�=�L_~_���!䊲����������{�9ڽ{��I���:�WD�Uv��_�BR4�T��8�A0ţ�(�	V�+���^���}��.��\3��*5~�����ݲ-��Vl����}n_3_\�C��.��&Q���Lz��e�uu[PV<��N����77��1�t޸�'�F���'����t�/�K/��Eˉ�B&+�Ġ+�ĉy�d��Q��R���5��UV���w��}q�*���x<N���'�9�*��2������X�2P�����e_ 7%9�ƍ�[.(����F���ȸ���ۺ�4���t���h@�(��#�<«�"ؕ��l�:�$x��b�Q���lJk��l�+ɢ�$ߦ>�F�e� %q����(�^��=L&�`����*��*�����ٱ�o���j�!r��^x!���F�9� ����%�Ř�Q����_��� ?�b��?��%����d>ߏN��>� D�hQ�ۏz,8��x)��w���~��-q8]`<����@X�PzI1a���?�l�ݳ[��E�b�6JJJ��`7 ̍���~UFݖ��C�F��0��5�VZ���iBj�����fzl�8��U��_rmjrܵ;v��Y�yN����a"[?`�����ӆ�}\���OO>�o�k;���I�4���.���χ��gѡ<'Y�r�*R��I
u���|��/�~kr��Q��~����tѰ �ZN2kN5ɳ5~da"��n�*�&����+A��ݙB�=�/�b�Ç12��3|�p�ī��g�c~��O'�);�/�ͣ�ؼy�]�4�l�FE%��'7�)+��`7��rR'�!n�Pu]B�茌���MtV3�;d�40�u���\�"��@�%L�6��X]:�Sr���:A�	�ش{�����B-�`�����kX��֭��]��u׌�LL�|�ry�.�)��7�ֱ�_Ε����!PmK����iE1�Uoq��K�(08��'� ���H�q �d�8QH�?����W��攔VM������ul��N�]��G���Q�t�R�l��⨳zQ�Ԅ��������~��]ɾ�VU��z]�1�!��C����/>;�,�	�H�lֺ:��oJM��g�(�j5�j��ܴ�����5}�b:Us��]�V/��U>�P�&�j;�����MP`����S(&ǦӆJH�Vk�B�5;?'W�Ai�Փ��&r	rrð�� |IuZ���r�u�%�X����tSy�~r�Y���;2�Wl�M�Y�R���
#�����k6��8VP�//P%{ 7�c8g�#�y意Kț���@u*���P�4�wr�J6��|q��*��dm�Cw�i�T�����t��qw������~��12��w��4c�L*��j׳[�'
�iݦ=,�� �9�x�/����GZQJ�Vh]~1��쐯����5U���"^�A��;�H.�1<��'�~���q�)q�v�>J{���ԩ��9��-��ߚ[>fԀ)�������<Q� g���t��wӋ/����&�x�n�W0�Ҡ��Z��J�>v����~�u�F���ak�wL6�Y�hMj�?B����вe����fZ�3��U�4V�g̘qZe;ꮽj]�t栾9g��|ۺ�;�X��@.�����*��cp���O,�m��e��VkX�`[`k0A��ݜ�R�,�5 9V�]`8��O���� M;���2w���n߹�'X�L}�}�8% !����x��ѻV�+T��G _k�`D�>�7������o��������ǆ>�����.�'I7J�!ҍ�}�T��,�ؕ�,ʢ�\B7����ߞ�ŏ��E=NGղ%�/��F���}<�z㭹t,����=nۘ�k���4!7��M
�UR���FG���    IEND�B`�PK
     t$v[���HT T /   images/00941d67-c746-454a-b945-4fddefc776b2.png�PNG

   IHDR  Y  x   ��H   gAMA  ���a   	pHYs  %  %IR$�  ��IDATx��w�%�y'�;�}��oބ70�0D"�D��DR�"�i����z�ZU��r��Z����Uk��Ү�Z��%
L	 9q�3�	��_~7v�����{�(�5�>�77t���~_<��o]o]o]o]o]������������uٮ�@������2^��{O<��ߍ�c���ҋ��X�'MS���#?��E��d������5����]�g�]	B I���z� @B�N��R�R	ˋKԌT���O�D��o����r�,��?=�����C���^^^�r����k���R��
�����#�{��-�0�{�a(��z���鿹�����ȵ����I�.��2F�)�N�#��P����#���^1�E/���<�2�i*�lnO>�2�<�2����A�}�^�-m�~����/0�F6��L�<c\�铟w��;��+����<�>?g�'+c)����X�WJ4�ܟ��'��D��朗����?�m�&���ٺ��hx�Y?��f6n}�)�t}|66�MK��>4�|_}]ǃ��Z;{�+Vג��7�����j_ܼ��G�ͷ�x��=^�����+t%�wk�J{�}җl�i^]���)�K���{_d��}�x|#��kL�>�9�Zly��s�1J��UyT���䳡�7��%Yǲ�P{Sjr�}skO������_�v�����g
3���~��R�G7�������o��\��/����=�9a�� e�`�a�K�n�@�>�:�a��a�t�J[�+B'��9[t0��n��[�I�:��h#v�]zF,����o8�@?��u�<�p�H���������H�b��.}.� �g��d���=3q��ZY�Obdq�M��N�bl�H=(�QYz�#������L��<��NG6�f�o62�yȽ�F��c������0���O�j�B�E�w����a�7�����}�	�l��\�x,���_��+���&�#���I����P'�V��/m��>����LH(�o��[H ���\vV@��u�}�}_U�)(��:��f��d�Ʌ��������8�|�8���}��L�`1ֵ�	����ݫ�Д�@�	u�'��p��Y�����T���>�<���^�	�^ڕ�%3�"jK,c$�r���L�%�}�pB��L�$ ��w�݄7m�d<��;C�$܂#{�pM�Ix�vd���D������zAI�醹�k�Y1�8l���������SO�������쁥��g��9f�s�A),I�z��܄?����闲Ƅ�����kP����I��C#�"�i�0pk�;���L��ɗ�H�E���7�mHӞ��5�!�,2�lS���\�`��y��$��I`�y�s��H
�"SvhS��L��
���6�I	�L��
��¿�='���הIXG�l��� Ne���5d&M��:�i�5�_����S�~`���I�=�m�'�l+�> �>{�
:��`3u���A����m�g�b�$�S�߳�\`f��t�9�rڇU�$;�n?S��b�:�i
�3g��s��tN]t��D�;��︬[���|%�@���$d���o.����q����<j��[\�~/z,,O?,c�ڎl�<�=�6�$�
�P�[X6s\�� =�+p*1��,<B�?#r�WCH m�H��g�H�b���W���ҩ~�����`��-U6z~�����J*� %���%�@�'@wz���H��H�^�!H��C�{$І3s�&�����|�<$�����j��/�gЏe9{s�L��Y��&F�-�-
���/�S� \�o����|f��8�jK������~P�*�og��bQ�ʚQ�`�����|�]0������p�4�A��gRx6�5\�#o.)�D?ÛP���{i���Uty�׃�5m���m�&)��Y����Z��f��W�$t�RGX<h) e{� ����l-ًLB����/�@���X��
�<f��$�F_k=sQ�j�x1��U��0�E�:!( J*��9$��k[��:?gNc@���&�*P ��b��2P��ʾ{r����p�y^�x411G���11�&\�:V�#~��5k��j���,�$��I#��AY�n�Ma^2�qLC��UI�ZU5��'h8��6�c��>3��L����Ŗ/�d����t`	��	o��XB6>�îk�J��c�L�,�S�L$���i����b�>s�-�����d��9��=�'}m�螅Ϻ���.R3�����+�^?��d���L�X����c��IVbg��+���h^(ڊ��-f$���%g��5�K��B�黇ߠ�oʰ���T���ڮ���5(8��������̙®�͂7Cr��^���\�=���2?̈́㌷��F���2YƲ�i�D#��0c�b�6�j�b�L3S&�^�AI�l� ^�?���$���{�� ���B��0b�z���)?��<��Ξ=��R;_H�jx�F!�:�
JN�Y���Aԉ��:XU���6��Sv�
Ӕ-��d�W*c�TSπx@;���@�4V+�[�͙_`�rس�oq\0艱KEGjs�	�~����g���$SoC6~����2����ĉ�����Y��tQdRn0���f��t�~g�G�_^������	A���� ��A(:i=�,���g�< Yx��dU���K���|\��U 6P�.�[����Y���z[+��M1}߿x�]�s���f��M7�\��5����XRy�
�@}�p!3='(SS�l4c��.�y{��8��q�5k�lŏ��75�^Nx�����W�����0� N����/�{��#�Z<'���N#�j�J�TBA��/(��lH�M�C�VXMH�j"�� &j��n�Ƀ�_0}����`C�S�z�J'�h�rO�UGJ��f�����]���bs�v�7��?�7�pf���[|�_E嘃1�Q�/e�
�"勎\�e��ſ���8X�y4�S?/��:͝z�~;w���#�Ȩz�c�Ne k�l�'�3!�rWZ�G�2T�����
֙t�G��9�&�q��l��ɭ�Af�~b���`à�YO��'�E�q�x��� 9��Ƥ6s�2�J�Ӵ�<�r���o����$��ǥx��F�@���|�_��+!0���mx����@oIN=��j��h6D%����F�^F 6ߒ':�|_1+Su��Q�	/&�ٔ��%��Z���X��3�B��2G.��s�;�2�]�]�⮆Mx���Vf�z%v�&E�bɏeVL�ժ�CXRb�}٦nc�0���;�8Js��xM�}$vw1x�v��p���6-�>�l�
8��=� ��5: �?S�p���}-g����@Ș�
O�����N޽(tG�)k^��>�����9��*��T�a�S�p�o���[is��l`)��c`�l�^܏�o���0Ꙁ+2:������en�,�p�)^�T�XX�B?qB�����ڢYH�<�5�~�3�Ǫ�%I
�z�bS���p�K��%�_����W&�ݚfU_C�rpO3�Q��n�e�q�8����&,�����(�J��w�ơ7yX�?��'1��OKo^	kĠ9�0�;���)bƓ�d8�W����P��h8�Q/9��8�6����U�8t�� l��d��$FD�^戅 %v	��"�Y
Xz=!�cCU�S1/�����qI#d�bd��l��s��F3�h=�F��0	�q,"c�^�{�ڵh��XZ\�XI�%VV�"
���D�������C�u�n�V�(d�⿷��Xl�9�ɕ��m~��0�8��~�:�˰������M�~/�
|@��"9��b?��rG��ץ.��gk��X[K�B
}�Y��$�� ��>�H������9��!�q���(b_�#;�,Y�_�,/��8�5߭���͑�-�
&��������1�]�-�PG��D�/�T�©��wD�m����R���P��y4�.i�jf�dS(v������N�+�8?~]�X1c���ygFy���H,�,P�QX*���;r�V���#B���q���� ������0�\±�fI��q�:�r���L�q(��D"���Aq7�񯜅y��X�/u좨�ɪ�1waF���N�2	���'�O&���u��m���~��M�����f��Q��B�
�(����,N�3�$o��Uë虇߁��f���N8)�v�wN�F��	#	�	\�2r�x�uL����k���>�1n�9�������[W�Ⱥ.��[�4�;�Y�$?6|�T�S�oh�9h=P��×��%ոo�����Hx�h`����{'�P����B[uLP���=#��	���r��8��
���͜�^���Z�-2��s!�����u���{;!���`���Ee�k�zp� kY	����}K��|f���!�����]��>\&��S�a]e�&�vhCQE�B��|���N�KM��l���&aQ9�*iL;�*��6MLa�6�o��}��˞�,?����i%�2u�Xbޙs��Pn��H� �tFsb4��J��ë�FXV��Z�hT�z�Ȏ�:�7F���3i�v	���Ҡ��plaG��X\�Y����,Q��-��F��X��G @W�<q;S���Κ��9q�Y���I��y�ۭV���^�mI��y�~ �e���6����'p�����D7|��@h�A�Q�1��j�62G��sD[[#C�ω
��Jh�J�$��j���f�cU0�{�CehTcK��㨓fG@�PM���#
��u��S)�#	��P��	4N�%�9[/�ą����0Q�Ӱ?U�u�B��4���>�<�@��gp&!*���zG�)����%�F˲�Y����c���̅�V7t'B��]�D�玧C, ��T\Щu4ih�qBS��{/��?����p�\�q)Q&����ҿi9V��E�)�'�$�\e�6�B�8;�X&i�}���.a3`�X�Th4�N��������ve������2���P4I��ơx�v}��B�m���	x�gY��
S��aD�WX��4�>`�G�~@7����W��bd�L����*§Q����Yab;.E��Хuݦv�_�Ǒ�sXUo�xo'ZsX4]Y�B*��KI��a"d>"Z�aa��L=cs���gXZ#-�VF�ZuX�l�e�$�L�*F���S����5c밾>�ut����}�����Ή�f�$�nK��+�G17�G��g�4�-��=�k;�l	�K]�0%	.IhW,�`�$ˊT[�ʛ�JG�s���
���K�H��+I�L]�o/௞Kd*�u�W�Ձ |uRyA��K��m�b�M!�5�9qq{lJ�EyfÿK
�(��O�Fw���L(�a����P����{-�<�ޞ����.8ƪ0I��i>/y6�[N8��X7)���:�ui����ת��	UM�U�� f�l#?/��MYiO"a�u6]�y�W�l�K!�AC�!�f:����~�{3��ܘ|��y%���}��2_ �T�ؿt�j�L��i�t����:�B�w�G�P�ב,�رbq�}^�M�F)�P,H8V��c��G�S��nf��4?�P������&.nO�*TUq7)�#~'�ᗲqh�t3�k���J�|� �b�b��?b˘6ul��;6]��S�I�b�T'l*��*�EYRM%�aUu��Q\՛Ʊ�^�p{�O�|Bk��\ԯ.��CX��J��,�P�B���#�#2�N	7J�%���p��f:y�y9-a"�ccT�-6���75��!�IZT@��Z�C/�;d��$��Y��6Q/�09QƎ�I�����ϡ4cq&�`��$	��h�4b�XS��ifL��Zr9ۜ���Ev ��2k�nvi�����;U���y������}|�o1�#�a)�f�c�6j�*B�"3fI�����g�ϔh����	�н��,L�&�];��j$�XJԞI���g�Oʴĉ��r�نŠyP����)*��a��Q�X����l�L���a�=�����_PV��%�3�x�8��C6Ѱ��4a6Dmh��n����|��ʬ���)q)��s+�7�
����S땷�+��q����x>8+1,�M��|��Q-)uc�����5�2�������Z���HB�b��ȍ�xL�Ar�zs�@�^{ڢ@�Vn5(��<�ٷ��u�j^�cӂ���	�'a�b�9Ml3MG��e�H��K5'��H��/P.UQ��`�eߡ��f�wM���SW����h�j����&lT�K��Y�2=�N�=JZ������1�i�c݅q�v���a�f�><��C�W���4��]� C��N�$�B�p��'+Ɔ]S*��_�%��+��>�;�]�-$1*4���j�Q���N �U���B�J4;q��Y��gp���o^��pϜ}��bnV����{]Z��V�[��y�z>�n��j�6f?���^��M��q෷��\���u���^��2��#*ԛ��u�a����9��.�]V�̀��[����XW��4gU>g��s=o��$|����xV;	�]VQcM,�Fhq��gb�n	��m��l";KBhؤ�����d��:'`��v�	b�J:1qH�;�,��/�Za�:&N��V�	B�v�ռ����Mng��S�X��
�pTg��yZ��P�R"�OU�g�F`���
v�m��=RWKhF=Ǿ\ё\=R��@1���uz^��Q��|�ۢ{������$J|�+uR{Kb�Y�[hQ��pf4��i�����-�MeR���ch�14�ϟB�qV�M]�U=g������o�;���r�������]f]�=���@����lF�Y1��"5_d�1��5é6��c�N�xsJ�XH��@�\�P�r�R�Ѡ>_Al���W㎍Wc�6�0��="���V�-d{��>+�\D=2�U"�Ul��c��:<t�U�8wH-�ؔ4��0�E2"yt��H+�X
�iW&˦��`�$�ڼ���L�
��X�o�S+�{ltu޸JXrf`ctO5v���V)�2U�x������û������&N�d�[L�tmiNp�J��IX�	jZ�.�4u�6똅�}2��a�T�X��͐���=����K�Ь;ي󋰨^�7*f�֙���8�N���[�����=/������W���P�j%�~�g�����'���O�{����D*;�
s�'x�PHQg����mۯ�:�P����C��f���ZE�j�Z���$�W7l݉����^�3���$j�8�T��ڎ�>֕m���n^�/~��X5��~?��O�y'w�vא��B#n7^���Ч�n��W_Ʒ��X�J�z�c�kO@�����z�����غL���#�}� ���;��;p� }�]x�5o����{�Q�>��6p"�n�֘u�p�τ3�p�!M����4��ۊŹe|�[_���Ӱ��cW���u�>;AL�7?�_��Q������)^:~ I�mS�5�D�J���l�.wR|�ӟŮM���3~�̣��w�	ӈ�RW�D�X��~��{���Ƨ�?��w�G�^��e�QJ.��簃���yx5>������a��=x��~�]�\2ˣq*�hL�ٲW]q%!J	{N�����t�U�t� �Q}�snC�D�-*ב�,Q���q�����-��M�bUi��MB�3�_	(��0(@k�
\��;ilF�@=	1�Q�Z�=�*�k�`���B2��-1� 	Ϥ]0U��L	<�&��&�ъ6�	&��\Żhq2��Ҭ�5V3��}�5�"]j^OD&<���D!=��Re��;�8v��xwnފN��Gg�@�u��]�L���sꆳ�|T�asN���,�g4d#��?t����_�u�m�����&X;�[˰47	x �oc�Ċ��ۭ��o�@j�M4����[�µ�qd��{�Y�4$0�]W���0Vg�U�6M�fm�m�v�*�w�R��;�=\7���?����f�Y����+��(j����t�� �c�&���|	��:�kx��$��Fj������P�nHر��-x�U7Q�G0��q���8�<+Ql��,X8�}�m���ke�*$����ô����:�l>�����{1o�׬ߌ��x�6���N;�E�䡕�s.�VKh�O��g��e�]-	63�=<��%BC�8�-�3<�Φ�κ�z�4o�U޸~;��=<?��@DL������z�.ܲn'FH]��Օ1�$Z��������1���)�vSHC�<��GV�=���ľ�_�Lk��G%(�����'p�밺>I K$j�5x��g�xE�ئ�o�Ud��Y�YPr(��v�w�z�Է����?��s'�L@+fF�x�X�h���ny?��I�=�g7^>x���Ʈ$"k�c��� [�u��dJ" ���� v��Fe�ܐh'6}h�<��aX/���r*"���Z-�ar: �۴��^A�=C�#��^Y��M�&-e��-�N|�<��Ӌ�B�;�j�Jx��\��
5��ư0��F)���D(�� �Y�_yy��� U��7l�^Z�g����o��e<t� �s�`c��lӲb����o�����gC�#|}Sv�y��������9���_�iܹ�~�6cEY+�!�&Z4Uv����L�����X �G�X��P�T�vY��]a�+�>��l�����`/3��ՍQRoiA�ʴ���g��v��ZKs2�aCF ��M�Q	��U�T��{������X�ٲ�(|�_bK��E�&fU���k�}�F����?�bkmfA�.F���v;�y	�6l���)s�8�{��0�E��<���s�+0���K��ǾAj��7܆�k6�p Qé������Y)U1N������Ĥ8n{<�>�m`<��Ȝ@��5��i|���0�1GRs���/���n�I��fg�m)�_��e�i(f���I�޳��^x�_N��L��9������qb�z	����m���#Z-��8)��#�F��	���Z��o/v�aO $���BsR�uS��[]ç��%?�>ӑ��%Ly���\�][�VbDkz��,+�RF��$(B���"591q�hڀ�X���L��y�.�ad�B/�R�xg��Y�i��e�q]]6�0ь�5�����pۺ�X8�@!�B�N�����9�u'���*fI��v�)j�*[���r�$���U�q�vl�M!�Lh�;���A�<��-�Flk1p�n�:�m�;o@���1A��{�^K�}�;�"���}F�V&C�m���q�b��A">�+u`�+��9d���g���ŊW�<3�o8&���-�� ��{���Y������ ���<o^|Õ
	:����=X�҈��F=��c���jb:۫�"����X�D�)�Q%l�\6�������w�p;ݣ��+���6D���v�^K�\���8���y�Ώ�N6V�9�̠�=7�� ��w;,�����T�2���!�\���)8~NcqS�ý�����(6n�@L�4�R5�w�NC��6�~�q��A�bK&P��#�	�l��s��%�O�Ƿ����M�o#Cc�qE��u��*%������=2<���zH��hE���!�Si,y͔YO��a'��:��ʂ%�~N���OȼqV���A3�l�kY^x�]=����(��.�ûn�]<�e���u[��d�>56Id��4�I?�(4�X"1�%M0���L6軫	n_�;6\�1;&�Ĉ�N4'��Ma׮��[`H�����^��q"Ji�_Mk���4��IK�.�h�-"�Ȋ�;�5ལ�%����OT��1�&Ӥ�ݺn;1�����DC�oL���&�ę�t�%�Q$��hc��n�rg�Ԟ.n_�O�}g�hF�,$�xv���kq1�ƃ��8o��m2�i�54���m$α��
l��]���q����3�<�-�*Y�9����ׁ�U{��)�av�a+��,-��%����qU����^h�ToN	Er��{ZSxi�����"1�f{����j����9��&����
�7�i+{z���lm;��7۪�^b�u��1�v���X�3k艹J|!1Ł���VᰲJ��=��ĊΞ;C��I���TSre3}��/W��MF\���F�6%�{�\М�����+$����x����;߰v51g��vN$�ܹ�aX�+ ��R�	۲9|��T�׊�/�}�Ez"�F�=�u�^ZV3@�<��)���,I)^���N0���_\ą�XG�'Ǡ�����Q��e^Q�ƤIs��m��vq�!H4�ZD���-��V7�b��5V�U�&
ͻd|r|{�����9	
��uCX�qd��5@��q�\���LI��Yj׎�ոy�j�ZGMM�)�W,Ɖ�,t��ҥX�ɫϐ�V�$���7�Ds���n�求������V�+�4�	�^�@m�Fr[c
��h��K%	�?:,�j��^�3��0-8���F]j͑�RŖ��8��A+��ܖ0�x*�6o q`���Ϗ�AC&��\��c99'�QhH|��S<h^d�-��A�u����N���8�L�o/X��GZ�B���z�{�#�/D�>u� ?�$*��ĎV�I�҄-C�$�}J\F�X�$
�2�r	���j�!b�=U�͝�"���[򘇑T9Z\Z���]W�F���mW�B�&e�C�Z�9T��4���ʚJ��< �np6��B�J�����[��sq���ӷ�~�L�=�jJy�R���6`N �Z�,�bHԆ8b"HZcg�g5�6�u�í�4;wi���g/̢M�Î6�D<F6u	&����r6b����0��9&r�ըq$�E�V�H���9�,,/ӽ!��&�V��e��S���NzB$D���Ks�G	�i��.1DC��s�ª<iN��S���B*�>4��c�a��c����"Z�!`Dwj�j?�S+dO)�"d��i��h���*vMm���5�fNQ
Q*�L�	�7���t��(�Q�bM}�'����
�2��W�>��ׯ4�����ԌR�F�\$��	���W�u�N��`�����	�z{���ۯ���xa�1�4;h&]�ʂ����$��4����r�={4^��<�P�o��Û]E�6Ww�l��Ίb�����¥�_��N�%����������i�v��j�-��'����w�;7_)�!'�����,�N8Y�d]�u�K���)Q�����08z�JI6��0ݻB���1\v�*��%��f�W��:��
��1�,ժ��+��:}���=X�>41J�j�''�!�(�W�坸��a�굱�m��]�cc����s�T���Z��:y���\�$T�~q7���ӨՄIr�.�5�ۓ���������bs�DN�YʪZN�A���J8���PC�9ޛ���K/���q��KJ��0m�7o�֍[�X`��O��Ҟ�nj��[���l�~)������@cq��Y<���4�1i�ma�1�	����5s7i��7n@���۩�:l��g���������M�&�X�-�[˒��)��(�ʡ�q�5�fwͥEZ'5�8[�����z�	�P:��9i�Q��R�(�F�&l_������<�
#x9Y����Ah��lr&���)��Zb��b���:��	�J�쩫tR��c���B��A	�=Վ$���q����p��ڏ�s�}UR��4�P�<�,�J�������{:<�ey�@�=�������" 2�������<nE��F�4�W%Oz�xʷ�x �4	h�JY͇�S��b�Ө���xLNT�	<ς�3ȇ�1�<x������?�~��#�f�b�c�Nvr�ví��/��Z��殲㫅�o}t����Q1�4ڌ�	H9�'(a��cx���q����B��.�HsH�1LNOa�U�		�P/$õ-8�1��cG�d����u�V�c֙����#�iR��{�[�!�Q4��v3�Ekg�f՜a�Jٜ�s����Â� �t��}�\��e|��{����HI#k�-�eiU{�]{��o�6m䒌��7a�K�2�kK�2t�$t�GL%t����^�a�,E�}p���{�#�L̟�?GRԂk�a\�};6�-��	DiB��T��!6uf��i��E��ɺ��-������:^;}��C����4����_��}�W1�~�-}��i��˰�FguL���D�Xe�?�p��XEk�W�����$$��ơ	l#�_꜆���zw����Y�����~������S�(��X�p�����҇k׬��}�[C�*"�7+4�]W���慠�nC{{� 8k�N���w����Zs�,���`�oks��6h�,2��ݕ� 
G�܁��g�~���(��4�{MD�5D�2y���pxm�����H͟����ǎ��ד�?�Re�nm����60�+!�=�����U#\�,�O_z
seږ!m^�@���H"�rh�̝AB���G���2p���O��}�Tr�߄��������Y�15�O���b�#5a�l����j�����~$q�%b0����8q�4lU+k�}s��_y)p�@�_L����!,��YX¾So���Qm4��N=N��V�z_��"�fg�H����bgZ�yj��nRe�-Nߥ{,8w��Wp���h����eTR=#�l�Q{���/>����8q�v��
���sLf�����������R��[���o}/�z#�cx���P��Y�1�EX+	��˴����́3gqn���������qth�͑da!�bf^s��dS���O��m���-�c�����chV��s�iJ�KZpy�B�na�部S����G�� �\��x8�1JL�X�Y;4�u�1����N�����3��ҐN����a8J�&��`��Ԏ��^���O��y���E.���B�����m![�^��i�U11:�*-���HP���Q���oH�����XL�d���?݆!0bS����8h*�����]�,��?8����q5ˠr$���'�����	��_��]%i`�U 긓oy����_��&�/,�� �?5"vĲK;����R*�����y�����^U4JCZHE�Sqdɨ;��w�a����/Q�yj3`���2�M]1���)�r֒�[���j"���l���,u��t0:2�f����ԫ(�+�����9|��@���E���^w�rs蒜�[�)��ee
R)��$$��#?.�d�D�
"�E�.��pNv�pW�.�k_�z�T���Q[5J�~	���` �!�]9a�Ͼ�XP���?�G�牍�5�����#,��?���2CXXn��f)w�YzM�}ғ�eu���?�J��q��ګx��W4���r�,�7�쬁{x�&�ӏ㉧w���%yax���S�h��$p��lG�uʯKt��1���+��d�'5�Q�8Ҥ��g�u:m�=<v_��_s���ɑJ�8e3�QB�a�Y��b�%K�U'�vx�>^V��f�bF�e��g��܉h�'�9Ӎ�%���1��*��R+����8q���8��4Hm�Ip�@�2v��5#���:1Z<cURII"�����;���HX��Ͷ�uś�Ȥ<�/������������f`nm����|���h=�ꡕ�g��_����B���2{Z���7W<ͮ��W+59w��O�{�T�XO"f�u�������+�E|J@��Qi�Q�]�a��x�9�_l�Γ]&��iw�juHm���,�T�m����lj�Zi4=7&Uz�T��{Rb@e�5���V��z���gN
Sb���,�ʽ��!�v�C�9R��F��.�LӬΫ:S�&�����]ȃ�K��u6y�psxߪUS�Ukx��q�=��u�i�?hTl�&�1����!G+C��p�M�`�����b'�vZbC�)�%.���+��T	�,��=�'��B@� D��8�������VOye�>���.�}�M���ۨ�v���B�� &��.<v8���pav߿�8s�$V�߈s'���1h��)��~�p>��0�7���TX��M�I�	ŪTIT�*4�-Z�e���^f-��g������ձ�R�-j���IDLk~��ɱ�4�R�m���%Rs�u�a��x�'�RW�C��/�Z���X��e�6{5��`P���Е��"	d2/+/W,2��X�Z�,v2V?�d����H�4�[ꁶ ��� �v���M:�f��W/�9W&ﲹ2�
�	��}���Vk�
WU��w�_�įb(�S'�JơURFQ��դ��/^s�������޽8�p��'�t R�:%�Xq����2e|�3_��kn@���i%eչ�L��:r��3{_���I��E單;����t.9W�ޱ�m����e5.��e��@���n�E����j����~�����q�{A�����l�o&�t��,�:	>�������i�1ʲYw�<�[�s(�Цhcg������������N�sWX�c�at]��2VI�ү�#�ظ]��.j
Mɗ��C�8����<^���5f早��?�(0R��/)�)SH���$��~�c�e�;`\j�D��4��`����d�V��s~S���������5����u��\$�/���^�ݴ�iU����>���5�R�0"jl���r-i�^"5"w8ځH�}�?����["�$rå�g�D5S$��L�n��F�83�����\�K�N:g��V�B5%���!~��T�u�Z� ���R�3�6ԙR�ަ��0���|]�����J��LCw�:�J�/w���r�,�)�]��g�-�U\�I��41AJ�;�-���j|������L�Y�:n��7�הQ�;IA}/+�G�\52�*;�8��\�5����/���33�X���Ն��\�ջn�r���_�U�^���Y�b��|���PbeZBn8��:���w��3m�Z7�8'vŔ-35�0�Z��׻��GbZ;16Ѧ������Bu��x/W#�'seM:���GW��!`���Uڱl�v���
|�H#�HV[���� �$�Hc^9ӊ����o�8TQ����>r���+/�]R��f@���~`�GX���j���ɩ%9R��s/ՙ���m�AI��#��7L����p��.afZ��E�����t1��"PS!Q%a��r͕�T!ɠ+u�c��w���[U�g߹�<��&�|tIЄR���5�|"��8�7���*l]������hHk�)��5ؼ�HP�`�v�v�!��FU����4�@"#��}9</0�V��N��a���r�dE�h�)��l�V{zL|n.5#��:Q�ρ� M*:Il6�r@uY�Y3�)K*/u/��s,v��n"��z$-�����Nߓ��ĝ_����;���E�m��x�5c�����)�3b\L-����	��3�[?`R���Wu/ra!v��s���gl͒��wh��Z_�2�#��Z܆���*j'�[����lݥN�;!���|p6Zv��H�+���td���B�U��kCW�T6���DbG�F�+8�Y�-�l3&�oR^/p�$��1��34���ȎD�u{�����T_���d}q�ٛ�뀷!g��L�d�Ϭ�������Ie�K�k��z�C��n�\�P�fʺ��&�'V���éx�8�5�g��!�V�x�Y�g�N͞Ǳgp�UoC��a�Ǿd�������'�pv	�#$|x>Y���B�d�*�� ��R��ѦQ?z�4vP?z͖ؔϜ8�m[��Z.I������H��T�9Zg�G��OA�N�׺�Jp<�H5�J�d�}��z
]�L5P��؀h�Ky��r`�9�)g
r�D�S�9��a%�����ZeLĆ;$��\�qǡ�����y�f���m@���x��5�H��xƗ;��g&Jj���r_�Dj�҆�s�,2��%��[K1�e���L�vN�5�ƹG������$��4K�3�\^߇W�^����)�rd]$�+19�\c�|�����~�T���8�����Ý7݂��x-�D±x9����2-B�{y����Y�0���Φ�d'ká9j�=1����|'�+�3鶻��hcT6��7'?�ْ3�8K��k�N�V�䚂�+4�@��o~�(���arh1̲��V��#�j˕�4�5��]�7A�j4$Vz�����Z܉s��r�Q�䩛�;tQEO2��|/��*&:���M�뮼
��%�4,t�f��xdMs�ҁ�X�l�<:�G�
���	�Eu��p��Ɉ��0b_C�p���w]�5���ǝ���6uhM?sF@���WvZE2��V6Z/�'@b��ݯ��]���М_��NB�8V��_cz�FZ'e�6H�$#'!�u[8p�ޘ;;V�S4��aW�?0�v��.�ٳOa��i) #�Ks)�	���f51:�Jȉ���8m�M���4h%1�1e����	��!���e������m"��4��)��5Q2�e�A�����p��VTN��������q��7�r���$Fch�[�Xۮnh�\�"��d�Uf5
~��G��/n�Em�CV�p d�2�V �AP�U��V��2�jx>��%�0�,*j��� ��'"0s���A�rs�&vޏo��qli��A���8�_l�Q��
(�Q�O��1�������!S��56�߈w݀��C�j����'m��\�@��8��Z��[jX��ҧ�6L��`��<���2��ȷ�ۈ���AT�e�:���G�$��l�t�?��,���iHۙ7G�8������q����n�.�`���g��i)�Ȍ�b(	)!i1��:����R�����>hpa�  �@�^�� {Ͻ�}���Z�^ a�;�lí�ߌ�3`���H�O��=L㤅�95�ġv2�x����	�B��g�$����3A�mnǸi��0>>&��t9pZ�U��&����{$�UN�d;�����W*i�@u���Ş��k�n����q�2iQ�ܲ��{IK��f�&eZ#K$���U�BS9��́��	��Z"����v.�H�B�>���?�w$O��h�o-a>�	SJw�K�01�p*�x�� V%�m(�
�=wFy�š���rvJ	�� >�`~a�#�8�� G���a�
�J�����J��dW�2ֱ������X\1�R`�6��`2Bd�/2U��!�\5?���mg]V�i�bR�j���p#����[=��WX��Dm}��q���O����qӺ��hTEs)W4���J�-��9�\ȹQB�ӥE�E�����W�3�eܰ�F�K�- v<b!K�<^z�e�s��ؚ�3�b�����03��DM0��z�Ya��[o�}߇p�U���VĦ�����w�������ïR�"I�����ƍ�ื�bM=�H�}g��R\������'1�v�F�)p��B��G_ڍ?��c�Ǧ��T��3��|�u�B�je&9�ƈ��l�QGؖ������ۉ]�Hd;+و�6���"�{��������Xg�����XgI�%ͅ}$:;0�	�	� �E�y���/}\O��������}<=?�o�/~�؃8ݼ����Z�87�
%z���+%,�p��U$����;p������(�߲�j�g3�;y
���񣗟�9���R�U�Bk�X.�|[��s�eE�'L��.?��XoZLd��H�m5%���^|�j��]�,�4SQ� 'r`] F���R��0��3%�˞da4��Ǔq��I�?wB��+��z,��ک�B������So���Sce[8/S��l"˽�l��}��~o]��b(Z�5���#֭�N�T`N�s�A�m���Bb";�m���ހ�|��XC�u,�\	�*,��^�7��M<s�Et��v�*!��ZWp��p����l���,�#Y>�?12���s>���`��zb�U9���h�;{�{�><���h���̾���z�%�n��?!��q�|�/Z>VH���26Nm" �ϭ����D�u���Mq��1����x��Gq�;�N����u^���jYw�|��e|�fF"����ھk�|�?�������a�s��K�=L����&��U�i�#�ڒA"�E����f���8�J4���Ub��^�k�]�O����HM΢w2�E�X�s���?����s��I�q���Z�b����V���g�6;�	Ɉ����߆����u��²s.�\tI�����7�ґ��(I˩���E�f�&���3�8v��grۚ]1�]����EJ,��a�zx���!@�ş�G�?�CgN`���I�Rp��m֤�� �#�;m9!�S�g�mo,�`��TH+��B_�2]Y�y,�Is�F��K�h�91�5����g99��v�mx3s�
�r�� �8O���.c�F�#�\�̂�CS���KR����,���M�ы�XU�SH�q��A����(�I�g�����B��J����L��.o�l���z靤t}�H���x����{�/�:5��^Y�r������6��ߋ�~�?c��׉��p4��UQ����?ZH,����ԫѓ||.�`�0e������w} 7]�6ڜU�C�-7%��]\ăO>�>�8}�TY�P3��|TJ�	���ԟ�(������0���]�n�Wo�5v���b�!�g5i�=��3x�g���G� 9;;�����r覌�3~��p��D���J����~>��O`��F�ޘ1�h�4������ϟ�+�_C������yمv���Lf��Tߎ���|j�x��/|����wb�!����S�q>p�0������Obfim�7Iٝ
j��L�;��g9�>�vYn�A�(Q�b�:�O|����?����41jbp���>u���װ���m��za#��䀋vw�g+,�[R��Tz+-wq=�S��	�wc��@�\�ZL�:�R��?�{��~V�ʺ��#�A�RÖ�h��X��c�P�V3X"at`�n�V9�����)�L�$�9���8�<�nI�HĹ[)��)�馜Ke;����f9�8�SDͧ)�Q�YL��[Vrb����>LMO��{0����ФqT��ɡv��HL��9���hjŗ93�'��K���k0��\�v�v�a�jFj����TK����ɻ>�/~�����ŕY��S9��᫝�(�����Z�І�����c��V9*ÛHE���ԴmD�3�=�#��O|����1٘�c���r�-����ž��J� g�0�Ͷ�]ږD H-�D��H�.�Vk`��L3Qiu�[ߏ����c���1�r��Q2У9�U�V��0�iM��������A��̣r�$̫���oRk��_Oܾ�z��g~WL�������C^	��ҽ�F��e�z\w��]�N¶��/���2�ݮض�a�
7�.�V���]�7&�[�����I�/�D#5�>�NGsv��&�>�y������n�s��t�
T��"��O%���|��n�@��(�;!VνⱨV�[n��w܎�������S�����}s?�d���.~��1�����	vm�ZJr�q/u�%J��M�=�&'������eq�=�g7�v���\�H�I�p�٬��v����!�u�5�#K�I�i��
�_�K_�u%��Y��깓8����ôd}���V�x:��:�Q�:�����;����W_�@�A�<.�`]\��E�E?P��,� }N�����q/�x�Q"�{�=�I(�Xe�M�@�o΢Ľ������ ��Ѝ��rt]�9��w�>�G��Ϲ��o���`�yJ���J�5R�b��)���&��%	7��"�f;��؆�Uk+�����������N�u@��s˭nNf8�RbƧ�Y~��Ɛt4`\ ��}�;�n���[�@��i;U�?x�g����+N8.���51���@v�5{�����׏Nb���d��Tq���.�\p�Νk�5:2��:��_݃����,�9f1��o .Z��+u|�waz|�����g��SC�)�F��]����L�>�(N�=|�4�q�=��"��,X����Q��"��j�fܴ�ZX���A�\ە3-ݺ}�u7↫����Dly������ql����l��T������Y����d`�X�����C )x����o5�mtx��/�|p�۟/\8�cO���u1�p{�k.�KϮ�����u��m;I�KDJ��jM�1zֻo��0n$HH[�a���$U<qq�ƙ�x�p��mw$]�KZM��y��	6�'P��$�ݸ Mo���qlߵ�o�����]\���{��	�M���u��Q��u �Ҳ�8YhA��%%�M9�&���\STbgI�F%,�m�=R6��6:��ɡ%Ia4���[�d�>�:|�Vu�Hl!���)���~L�f���H��M̳�b,��������R"�:��E�j�C��sW��j�cι6.Pַ��8�~"�R.��.B�$e��pjI3�^����S�^<rⴄ�p�+>s��j<0�Ը�����R���<�MB�j���WY>V��'k0��]��z��4�>�O?��ԕ�����`�Ԥ��k\������R���V7�_�7)��
�s%�� �'G�k(l�8!)Բ�����,�Q�~����Ne=b���D�j��z\6����Lf�HA�D6j��Je'����j]�ŖK{d������l�'�8��%-��VX&��z�2�4���|w�T-�Ҩ���$���k��;�؉�/ϊm�ג�p�"$b������)�Iwf����#{T�9|9(u���$�ɉ1�D��p�&���d��|�ƮK}aç�r�m�lbzʹֽ�cs"�
	�����Q���|	Ov� ���{��z"o�
ڇ
�I�O�h�w�h5ak\���W��bÙè����r����eʾ�yd��: N�|�=-��nȼ�W�N��xLu�'���r�V�u.ZDԭ�� k�	y��M���: 顋yR<�Ν�4�sR,��FT�e�����r>Y��"0X���)����v��c�N����V�ݳ��
�l�X
\��MRa��xp��̋om
�'���7���
\|��^���F;���JŢ�Y���3���c簱Z��E�<G�ns�^oY�a���̋s��t ߟ���d�=.�w��i	\���&�<Ѯ�]3�p�83IN�d!��)�5Q䲛|�]�S�3v.
�S���Tö
9�1Β�c��и�8��L{���MR��}��vP%RH:��zb�"�\�o������X�Q�GU��
�������sg���Ú8jJ��S:R�&�q���uz�dG.�sj�'3[�����eRX:N��j�-
s�,&+)���T܄����Jzh���sܤ�V����L'�"��%���t �."V:Gc[F^�%�~����99��m������]���J�9u�A@��l}W���ƛ߂DR|;�Ox%�_ҕӬ�Cg�����E��ĵ�,5K2K�����J؜Dk&Nq�4��N�v�� 漆4"N�O�uk�?;X$�B۷>�6�,��8���!�+��//��l�+��M�_�c��J��.�P�$ug��L�&��bb�d�&�d����9���q���▬�1s)�$#�`�ã���=����,o>�w������x�ş��s3�j�S8u�HsY]=Q{�F�*^�FX���9��R�+��7Whr����������3���1�/
�������%I�C=jH�e��to��qMNNb�x�ˍ�djq����9�v��F|�����<Ԇ2�ä�?��nL����<�(�?�E��sf���fZ���w�1'^�k���V2�������ɇqvn[�_��<i,�fM�]��9���H��Dy�J췂g^܍�x�@�*�������"� ,R����X�8Nڨeγg�6W�/Wh�	\���-I?��Շ�pb�<�~�%��D�E��OYs��(>-Ey���o?�#l��O�/���;t���)���	gSBH�?v�^���G=(�pƖ�ĥ
N,t���M���=�M��p�*�'����&7�ٞ�*Y ��;33�=o�.�>IDp��D���E{6Ѣ.?z�a\��*]��.���IWg���(?d�3z�=ܤy~�ŧ`j�ד�d\�u9"K֨V�� [ZDB��I���{���~c�'��qN��ʊ+����7�T2��5��]/\�|��ɧ��x?=�
N���D��6��5[��B��*���b].��]�TV�B硁��2^�x���*հ~d5�*5Z,ee��r��Yj�l� W
�`SC�]I���gg.�g��έ���p(^�+u/˜e!e��V��bp�LNU���YS�L�wo�6����#����;���l^P9������݅���{\��υ`7�@*U�Z�����v,��.�4T�E��N�ڒ�q�6�Tpt�4���`��*L��)�2 us��Xw.�vj4�q��cRk@�zt&����y���:����!�Ā�|�i<���RCV*L�Bو�ђ���#d�!U�xk^�,�{�K�,�[0��X�/�>�̱�x���P녘�X;�JTlΒ;�4Gc�s�Ԃ8�G��Ϣj�Z�ͅ8
���Hj��s���5T11<�V=9�?T0KRV��Ӄ���$��S�����:MM����HU5v@��`玫���������� I�6��z��c�Lr�\O+tq�:�\�zm���0��e-�ޗB�%�=�����j|��%�Z�lחet�����A��t�Z��{֢�>���Hz�d��4FWKs���e�z�+|D���`����7Hq�R�&E���?��;�Wޞ�C~s[��TH�	H){}~?>���X�8��-�/P�#�7U
mu1d{�Gg'!��#�a�����זϢLz�U7c�'��J\	O(>�eə�V*l��VR�Vy3���m��p�-׌��/?��HV,��진+�s	|VG��D�tf;;��y�����6�-T�����2��O)V�S�� �qaa��R����2.����g�u�V�}���|�W5u�S��ha&��t�:!1����9�4���q��4��G���/�TgQJCv�*�R�Ff�e9	�J}�ER���s8t�$T�ܼM�`�8qɺSgIݦ���Ha�"��Q9�" .�&r�(ض@]I�H�rFN�߸j֍M�	q��a9K���c���/街|��R��Y8�ܢ 3�B`�-t'��17�?��O�0?>��B_���s��i٪a��}��'�߰����,l��F�s]b6և��z�Y]\�Z��ԾMS��;?�k�]�C�����sI��1�Zl�&�X���my��ɮh\��+�e��w�1�rD���z/f/�g%;ȆH��^��������	7b�-�b@��'�Yڸz�Ԯ]j7i�X6'�=;X�θ�2N�����%�h����%N8W��.�֨�b�f��O� b5����[�.�T�E �W��6���b��jGZs�s�65&��5q��il۾c�c��*�[_�Ɍ��8���q�VLf<�<״��?�{��{��Xc��Mri����O\���K芝���W_S���iMڮ G{�h�'X|-��ۯ��&6`��Ue=iV�����A�6�R�+�d�+�|F�k���9�\�����wg0S��m�:�J0�	���ߓ�;��IOOmR���)�9C�;�.s����	��fw�FX��y��t�t5Xmnv�;��l�6��IlN��C�-���<�_�¯�G��C�>��h]��l;��F�I�gzl
��_Ƶ��E_Ý�����������1E���Q���*���	F��c�g�y�	Vw�<o�f��	$H�Q)�V�-Y�Y��]�^�V��|����ݮ�k�ve�렓%�r:�DRLE0@ I� �30�������W�ׯ�t7�̼������W�WAʹ��{'��=t��[ct	��_;BGO��S�/HۧoYZ���%����]��4Ġ7e��ҿ�~��~K�P�������S���=�e�F��/c�YO�ʢ���~={���2N!�N�xc�*��e�ʽj�q�p�x��裇��^�q�6�%�6���o�L�_��Ν�Z�]��)�?�ܴ���s���l�5ф�d m���J����z�[ށ �X�I/|��>JaG �[*|vo��/?!��iFJ_y��t�����j�] ܰM�����Ѻ5k�ǿ+ �e����{��1p�e��_~F�kQE�+�6����aڰf#�X9�z�}��O��9q߽��F��&�N��媐T6��;�!��^1C��5TA"!�j�<��c҄��Q�~�,y
M�c��3H�3ct�T����\��Ϩ�_;Ɗ��Nb~ݶv���ĉc��JvE_?�cܐ�#Q\��*��_èÓ@��Ěsҫѫ�NсSG�t��}E�4C	9�*L`���jc�&����Թ����L�#	]�'nI%Ӥ
�y~�"]z}�6f�鮍7���!��2r�6���U�i���`]���r�؝9·�ڞ��"���K�y���mH7&�l�n�(�dzg���E��d�!@���\)T�c,k�2�8��;�Q�� {����b�o�},����C�I%�*�q�䔬0��Λ5+�ݷ�[w�A�Wo�G��-,,��m.���?�h���N@,ܑkg�n��ڂ���ۺ^�{J��J�6v�����7�=�)��0 et��:����{���"={�E����-+�%Q�HNz�FVK�|A��K aI�^ɾ�;i��G��0}ca3�t�o����.�2�_!sVN�*�gg������RfȄZ�J��<3O7o�E#�.�[������:��B����PMӔY_��b��Wtt�'>�+��'��b���u�biI�Gm&e˝�D\]��p�#0J��\�����%�u�pMN���Ԭv��
���v����=��D�,;q�J���sD�ĸ�:u�=�{ �T16#�7o���.¼៺�mB����_Q�#�
u��ǔ�vO��zڨ���^x�U=r@�U��X���;NH1�;�+��};}��E��S�_�ox�fjsl�RF���ܼ�>�s�b�S�}��G����7p���ǋ+�e؊A��⪐�W$��i+P�^��c����U�s�N�~�Fʔk4��A� ��[�貹�w/�"�1����uNO�Ӌ#����+�2Uxu�[�Ε��t|}|��*��]6ݩS+�l�яb7�'�����Q/���Y�$vB�B}�^}y�n[��n]������/NQ7��m� `OJ�<{<���4]�6J�g���e)*���<�4~�N^��ya���e�T���ls2#%V�:��9�*'�f�[�_�w[r���N���]�%&HV�h�l�'p���*�:^,���}�{���c�ܱ�?����7�R� �����(�}�]�×_�o=�ki��im\@�4��j���������E���fB�Jl�r�"jK�-7�#?�!���Y����d�<�P*-��c��}��)��O��2
�x�]�j�������Y�E�k��%Uͥ
�Xɲ��VVv�N��>9;Ac�R#��+�802�Y�,�dZ�3)g�g�k/>B�|�Ct��7�٧���חF���0���(�ţ�N�@�2���(�az�;�C������7tiq\&�!�i��S���R�U���+��`w/06	 �?���]����^�&J��ɋctmbR�[��m^�����L����]ȑ쒈��hI~�U�� �x����2�T!J���.�x�=���Q[GA�Ȏ��б�'i�ֽB���2��oP��E"� �lE���KJ9YIm߲���@`����ԗ�d��2��J�zyr5�2]��>@�{+=��F����|+�r���R}�#�Øo��ʍ�P�\>M�~h�����#ߧ�����ik�J�gr�/Ui��w|~\'Z��7�V��U��l�F��5������,�ח<`,
�+�G�<k4F!�ܴ���;V�!����W�
JkB^\ M���F.MXЏa1�����4h!]�Y�Fc�蕉˴�w�Z��6�;y���O�;Q���❺t�&������H/\�+����5YLר�.���9j��#V����X�B<�!+KJ�=9�̺��<�i��!�Z�\8_:�����eԸR�$�i���%H�-<i(!ֈ�b��Bh���P�2���6��D�.cp�M��&v���J-9��N>x�Wm��|����o����2�������~o>��L<j]|�O � ��&ck���n����o/+���b�A�wN�̛cC���b.K��~'|�(=z�����{��I���B.d�.$
م>�g��	w���:~Df9�X&i��Bsa?��w�'����Y�d��f�h6:��Ƈ޶�<�t�q@7��^��$�� �Rހb>MY���~�[�`�����g` d<�&uRd�s"2��GZD�?��@�n3����>V��Y��}�E��jҲ�+��������~�?ӡC/Ӧ�=�X����^��qyZC�-���R�|,����� {
��&���<�����?B����C�/��]��O��5y	����=�&�Z�h�'��װ	
�0���>�VҶ�U4\� /o�ۼ��2 ,����������)�h)ey�e��!�J�1�6[�mC
Ȣ��U��d�޳<�1�(����$]<�H+���5�NZ�(���B���!���4_^�k�t��<]f�[b�[´�	�Y#Ӕ�P�Y��葖�걷�j�->Y��DZ���5#Y{�z�h�Ә�J�wi�JH��TKSȂ^Gf7��[��g���ޠ5�vZQ�>vW�h��|c�<�^�B#%ZD��+�(�f��V�g��#	z�H��u�wd�)h�k9r]7r�U" �#�M��<�F��{�V�@X��(���"��^�J''$-{�}�(I2�][�Bܤ��B��(t�=��!��[h��z�w61�:E�9����(���#�|�f�]����Ƭ�j�,��0պ_߳鮞/��$"jh�������+h� +F�����h��aڽk�^�Q����0�e�Fz������k��Eʭ��'M�=m@�Do� ��dY�L����,��*��ZX�:�Y���|�6n�D����&s�a��h� Ґ���&ׇ�g��V�@�fY�z����K~���������,mX�N��;�?�/��>�W���x�ں
,�R ���1�A~�2g��( �:�����ӧ�������4��ïe�oG�\K�#���L���"���v@�X��4�j�Pc�������w�/��)N�^�eT�o~�7����ҡ�YѲ�,�����,������]��s=Q�� �j�i�J�m��dH"��(c�\(�9e$�vx�~�_���ct��̳��a���LF����� �/-�_}���u�E6��Z�\�^0���PٺЈ�i=Mj�6hCF��\����1�p�=���{0?.秅3"@��d����Ժ�k�)��!��EJ%e���Ы�	ܰ 'Jh/��ܙW��\���,(����RM­����Q�JTÀ8F>|��D��5�1���@��f!��k���	�`V�>��@���hk�{];�����ݟv/K$%�fou7j�<VkoP�,.�	E�i�����a�Y���]r-M$��ߎ#�]��ZZ�c�Q��K��w���c�e7��[��)�ۉ��#Ǉ��3tﭷ����4��Z!�qtatJV�e��K,�$ ]/�G11����$���}�o���_=O�6l�5k�So^��6v����+���0z����Iŭ%!cT!JG[�J��@��k��u�����K�p� ��ha~�^|�yZ��'F^���9���dZ�(,cia��>��"$τ��,K=�6z���hך-��wHbq��p�N6"����Ԩ�;�Y۶z���[��������3�/���d8����F�b북Э�X�g��蠛v�G� #p��$�ob3����׳��@)yZKe�l7P6�c`H+ ���T/U(���Qi���,ý�����'��_����+t��;hu�0e��I	�ذ�Ő��c������ O'�¨�hU�Y��b�m6���y�sę���2�lߺ���c��*2���eg:���L7\�
e�F�.�L�E�<�
�w�q� ����`|N��){��c@�$
�c��,G���L�H<�]oފ�eW}m�p�۸����N�:��ƅÞ&��:+}�̕������T��&#�Z�Q���P��Q<~B&3D:�B(�p����d*m(�/�h��ݨD�X�z�14��&u>{K�&�1hL���-HBѺ�IA�YӸ��NZt����N�^����D��2��7Q���*��o�]����Oѝ�n�w��A�g��2%.0@���������o��mbf�ʌ(�P���D�I�)�Λ��`���k�A�����h'�b� ��_:|X��޸�FF&9ڽe�ڸ��9v�E$\��A:AW��}��s���N�9E�~�Đ�y�o��:�󴆕����$�l1G�RM!���0`1Ӵ�o*�0�*\��*%�d)�Tw:K��s�H?u�OQ��KV���?�^E�W��*��yĠ��im�ݽw??s�*�T2��9F;k�p��1"M�̗c4�U,���g�+�A{n�)�g(�G��/��Ghӆ���jJ'��1~�*R-1G.��Eó2��:�K��c�-��=Vf�Scd�֦gr�������j,�mE�H \X��_�{s��k6�9�5� 	fP9��������f+����+#���
.}�K��������syofg�7�u
���r��"kj�`�I�g5ɬ'r�Im������<���؂擯WC�<�ؠU:�N�D?��h����P�8p0�J��D&WN��ۗ"l_�a�[�dm�$���YAq��o~���_�l퐀�萁������^�/�h�k��oq��֥%Έ�X�
ָ�bh$��j������%���,��6;�V�q&$������!�(�	���;Oԩ��	Q+�5���&?W{���h>y�7�BxSڸ��j[(�����+��s��D�;����غ��2ՠYW����p);�zɤ��M�-K-'#A}z�<mA:u�4-���EVm�۟�MZX���kWI|1yԥ.-.��L�j���^N�_�u��A|�N2����pj�Ɨ�,�^=> ��>I#׮��N���;�����6k(����8]��Fs��\��:AҺ؈Q��g5lt����C�-����U+�(�^/-5�u�v`���!P��!��c$�P�0��$n�T�j�j#��g�Έ�\h��J�cgN�2���6A�C�=�⮻��r(�m�-�`�q���\�s|�����Hs�뚒�L#�%�a�K����+/�W��5��_�5ڲv��C�P�(�#p佼�s��/��"ޙ1`	�h�����R6[���.��w�MF���-��s����xV��;��zo޷I���鰃�h ��F�ȵ��Y	T��%M�����J��Ɉ���
����ʫ~h�y	^g�զ�ֺ*(������f��r�؛>����F����(�	$DZa�$K�D1
�?���"� ��#�&6��3����R0��d�:�@=Ĉ�fv�)0�M�um��H��z�	eQ�P��zR�(��$�aD�⯾sY͵�°@�^���%��%��	����
mcEkS\]!�����d}a�B�')W�%��
ֺ=-��/|���<E?�S�aᾟ��b�j���\���'�Z^$����N92��b�p�`�QفQ%��\���ij��"+zzhhE�`cZ�=�e���u�]��i|fJ( ���%]��ӄ�)z�	��.�_������#��$�~�
��\��JIh9��?��
WZ���B������ZF�?{��=^�L{6�,h�Rf�^�W�-И��I��@��R=hҋ/dW�l�A��Wӕ�Q�!�)[K�`�3�������s���רoeY���&�u$�+��ӁM����k|��(+�%A�H<W���/�BC 1ho��l��� �1@̝e��W����ѯ��ݹq�z.�6�#/���ϟ��Wβ|U5A�@M|�=��n�r�b�D`'
��sdy��y��¤�������� ژ����<�(�%S��`�AjS���'@� R D))�� ��&��m��^�( c�J���Y%�g~�MI��X�d�ܟ��V3�,.I|�B�`V�[Ôm�R��P�$��#&%�����b] A�(Ϛ��+��*M%�Фp�-�F��nW�)��dE�2b�����XK:��0�I�	��I�����ގu*�H��M�&�+Y�e]=��@��
$�o�!��
��|k�P�ӧ�|g�f�%�ܗ�@�{�Yz�����z+#��,��Ԉ�$�h��Mj-�b(�2��m��T|��_�_z��������F.PJ���ʉ7���E���[X�(�g���Kt��el��YH���d�D0}eC��7�~����i��&ʁ׸\�Ӂ#������:M.̈���riAv�3��q�{Zw��$b�X�Ʌ%���������o��K�o����G���/�ң#�%6��������WDߴi�����w���+��Af�as
ɪ)��������_���;��FY�Q_�y��iz���t���[X�NI�*T�8}�>��K�ӓR9"��-�u�*'9S ����왥9	����:6&0��~���O?E���?H7�Zw��{�~p���w_�
][��z�)=�㌐ZU/�,�%�	W�{~��1���.��y��fW^d��G(�F�j�o�3�	!��l�sK"���)�tԚ.�	W_�I[��n�:ix�윊�R ��DFEJ�����նh�$X��J�Pa�z뱒My~L��m	Uن*p
Ĺ�q"���Ծ!=L�D��hw�W�kn�XS�L���Ӣ�I�>bE�1�V7�ҡ�Xٻ�O��h{�uɰeZ��W�J ���^���}'FS�,ЭI1��c))��4�����%��W��ڑI�u��0B���<�YI���>��H���+�];wK��&F�Գjq�Q�?�k<�(@�r��S�<�+Oz���Q��r������~�%t��������d4�?|�Fg����3�Ҍb%EZ��7|�xf~|������Ӵ{�Z3<Lm����f��z���lL�~�x�;t��1qQO]dtk�5��F�Q#�2��u�VF�3��4?IW>A��Wi��m4��P������B���פ�MU�4yJ{W;�.u��K�tef�񂐮��j�BmOF~��i�t<~�<�ޟ�!��{?H�J��~�,}�;�Ѕ�en����߸��k�z�fY	f��$��-ū2+/\ʤa�a�d���\�{�`C�
�r�$DGG�п����`������9:�h��� �U�h�R	9��?'ʛ oϼv�*�'4�b%={�0�1��1�������!��AnZ�O�s�� ��+͘Q��H=F��oZxR{]}I�1B eL����8*\a�PȜ�����:��z�A��Q#�a� 1~Ơ����$"�B��e\@+�3�Z�g���Rt��M�%lDwݒG��,�<������d=<��U�zPg���b�v29%����m�'��Z��Eär��qJ2���aK�h�G��G���XM���#���R	�j��oh�,6�N�2�^Rp�9���*�2A j����:���eP���/<E_?�>7�1��p!%�p/�w0�C~lM$2(-1)���7ɇ��пq��۾��o�B��3�ұc����X�F:b4{�^��c��	v%(��L05�!j��|Q�����)��뫋3t�����Xt�� ��S����3t��I��w���D*�aá�(�þ�h ����c=�'J�~���:�[����ڎ�;A�tS@��_�qKP��`p#+�s�c������~ߪ&H�,J�B4Ӥ�z�����1�Wf'�~�τ����9�}���B�G�W�`*ȀA<M-�R"֔!�B��WjQm�GF�^kJ3�?>�M��GE���W�f|����45���k�9&���%�D���RK��H�|p���8����q:�*�g�i�D�$A�So��x��%%ţk��@�a�5��Q��t3[��&�!����YmX��b�hB�6=��U�����8�i��YL�saA���V�m�2
]����Y*��Ԯ
��"�F�Ёgb�nJ��*�`!o�������%{/@�:9"r����)��!U�~����_���д���DH��VRʹ��ف����J���mM��z�U �C�-�+��b.m�3T�Mq�ޗo���tJ(@�졨�y�쬎y�kL�>�(r�	�Ơ�k�u�xp��� 
A�LS�V�X3�۬�N���3��~���ёQ��S�"��� 4KYv	ˈ�y5-��(�F�l�t�|�:
� 2Pi��[j��(	����4��5@ВV9�JEC�ex�+��(�q\��q��d(IXوҌjY�����#*�)/�j:թ�:�����vIn1�Ԧ3�M�I1�&�0,��w�]�RXVY@���o@C%�<p�K��&��U���]�I��"u-�/Nq��W��$�?�5�Ǉ!F�Au%r&\�F�+)�1r"�&����HM�M�H�Q�F�Fg��뤲��$�⡧�p�L�F��T�"G���X��v��!W��n��V-d��3m
VR,��T�,���[���@X˕l���	�l8��TVcc��U����&��eT獖�� �r�-	%�0qؠitfqk*�߮�[�bk�+�H���=�N���y.��U�3�0��M�n"��%�"7��U�F�E��W��މJr��{��\�7��Մ[[K��(�>|��2Mג�k�U��wa���^\�'?G�a���g]X�"�;d͞y凴��ۨ}���ъ��EO(���؆����#�D�z=��qȀnR�W��d'��I�!3J�j�2�j'^O�:f��R���s�/-o�2���eg�=!���G�S&�(�b�ڈ�$ݓ����e�rz1A�^�h��'lb����0�&]��^�:�Ռ"�/ݎ�<_'���p&R��\�b�=�$�����-1��kʄce*�=Mp�XɎ��y�,8���K<�F"l��h-TdH6Yn߬)^�W����C��ņA�$E<E�شlK�}\µL�.{O.���c�����L'�z�xQ,�xK\�@J��<;YI��6�Q�Z�/2��v���n&ʂ�w��3�+���*�%'��c���(�_h��O(YE�6�+rB�B"T$Ɗ������$[�C�n�����Jކ�FZƋ�Yy���,��>2EB�Ģ�Zi	p�"%��>M���j)��P����_ƴ6����F�G/�\}���'U�Yf٧,�2Ri�1;2��u�`�P�ϗ"��ܜ�C��PF/�L�}�r"C�r)�$��%F|-�.X�B��4"�(���Q@���+%-�^�U�����;rY�PUHr��I�!6n׉@G���g�*�{��ʱ��GX����\.{Q�±w��6�udF��A+5d1��=Hԭ�g�>ԋl���;%�_�jPqk������"��и�S�
L"�)�&@8%�i�gB�z��Z�W ���
<�ÖE���=u��:����B� �\ߞH6��:/����˴��ȭ�*/<�d������0D�	bld
�)�T�.�t����܎Ǜf���!wG�*&ୟ8���_��~�%�b�"_]q�|+�V����b��_[�)rWq�X}
3��%���(F���o�=�)�)�`pq�H���jn-9,$w�_�z���B�&CY�&�߫�-@�������+��"��;���]��/��7*N�$d���"�+��Kn�0�G�P��� {bh����JZ��U�[m����%�W!I+ue#l�D>q�&M��ۂDˍg21)�c��<%���A�3�%-����()�T���i�x�=3�:�ڸ��߁Ied�˭�{����9o���'q�8�a���Y�Ō��k�_�H�}D��(����6bt���g+Hp
������t{~���Ԓ��B^���3��]�d�m�Q�ڌ/�x&_���{�b��b#��_�d�.~`���`��i| a�4�T]�J/�x���)S 
!��B$�ȍ��E$m��'�o�H�t2�YYD�uhmB���� I��u�:b�bU���ǧ�nO�-V�_��x-�rbBvS^qhF$Ҍ��'
SnmI ��tMn�e[�T�����j	��h1�*zRo=�&�D�p�Z�E������[�is�e���	1�{��e�dB΃q0�2}]��.ҥ�#�
=)qHO=�?��!�V9I�(�TFc��w�!ۜV�k
���8C��A�=8
��Je6u9�`i��_&��v�M%B
e��ˏ�!w =��;�n��o�2$��R�ח߉�F�	G����Y
�˻�z�d:�)}	��6�qL\O��HD�BqS�J]rX�����Q��6LF�V'�<�O1�h:�dɧx�S�?<��@o�3�%�z`qۖ�q�!Ҹ�=�&�")��g��x���H�!�mGI�P��r�g?Eq�B���-��e�|]���$��GKW%�j%۴2/�~��p$�n{���uqP��k4c+�l(��t�45��`��V@g&H��p9�-�wd�cI�.�%HC˩���kj2��&��B��bFz�,$e�З#��a���Ы hi�bd7X���1b�_(�cB�Ho�oO� �A�T� 	G��F6�B� jj��
��ݐ�M�(�C]S�ڼkQH���L���b�.qH�֦, i�{F��	S���	E٨��<���͗�),9�FG���W5��kU�UP_�d�T�uC<�p��^��B��l�C	rm*M �$ա�_\[��/�kW��{y�
�.V$��X��0
k��1�օ��gJu���V㺸jZ�匠VT�) 8��D�9��Ql��I,�b����@��	�>*-�ǳϷG0�*<#�)
\�ҲR��<k���4�� π>����۴i#=���T�3�����\>O��4::&
�$����A&�-�?Lv��s��L��,�د�]\׏T(g�&�bT�%4m�4�jJ��	���A��Ny�[^g�d$7)Z>)ŭ��E��:d��4���D�}d�d����\�UP���iG�0ݰm#��Hh�㰉�F�&9�<, ���Z<���r���0����n�����/I�I�Z�d5���gÒ�j�/Fn��ާ�P8��]5�d�'�Hгa������(R����)�� E����x�����:-�����k�Y����p��@��f�ˌ���º����F��b,��=��T
Y�@� ���P2�v"K<������gb0�TB&&�Nk�lR��f��o+�a�_ ͢�{inA�]��b]М��,����^q�{�ef(#�p��C��ZZ\�}�5�c���@�:����M�����kI���}==�+���S}~�6���7� a/L�=q��{���d�q?D�:�5BO���V�D�Ȩ2RW�����0d�2�h6�W�DB��We$N����t$%��r,��Yl1�D,g�N�@B��B�$�5�R.��9H�R���&%��\G�W�I���b�co�J��PG��
*� �0K�KI�_![���@�TA'�uZt����A��bg�� d=��`IϵL��=�l��-�S,�$I���+I���	Z��fP-ѐ5.b�dz�3�,b&!(��6������q["�p����="�N<W��</�d]�pH<"����F@�q?�߱�7)��,AZ	���8t�����\�RF�����qGU,���@�|5C�'�"s�o�g�\�C���JW*2��.�V	��!�R>���⑶��nH�xhG?O2̼�P�P�s����]�C���s)Q�x��M�cA�,��O�޴f�ɕ�D6�Y�7y�fc�����7�Y|+�'\d�M!^AS���_{O�`.��FP'v���� <��-�&<3��L<S�,�"��)N�(Y�fx�.(�LZ��z�1!��:��ǎ���$͌���۱v��/�2��}X��/PGG'���9s�>�����K���Іn�ob��DUdh�B�Ӯ�n�b?;WPOw�����p����h|�d�)E���Ꮾҡ˷�e�ʵb.2(�A)�Z� ��v���fJ�,dkvj��'&eڭ0^��B�R��U��{����
HR�U*Mͫ��=Bb��J���MF�@aW&hU� �D�2�.���+����g�11���)�*�j�<�"��p~A�@���,m_���o�L��2��_�%��WU6$L�([��1(�Q]���N��Eƣ�b�����*�8D�!&5�~�ȋ��ZJ*Y<�Gf�7"�&ɱ cLF{�Hml�����C+�!E[R�2�I1:(#x)u�X00Kb���X��wBƚ��	63I�Ú��&��"F���Pc��75�$V*p���	[1*m�sSwq���R���bl��?h�K�,�ƌ=�����!G(���3j��Ƥ�b�#�u�O��"I>5-&&��x�����Z����M>��A��g�c	��^7�,�I.����D.
�BRH�c/	m�a���:��#�ոjU(��g慭��� �s�Ѿ�]�5�O�Y��g�H�Ќ�dAM��<����&^ՍnJ�IP�(�Υr�֫�V�*>xH�&V��b����~:}�����u�z�re��ML�'>�I����K�T�+J�FK����Ư�fS�)�A��Vez�(�t����%\��J)+����̎MQ��
M◤�!5�`U��U$�j~+��ߗY�
yy���E�tt����X1/N�Re�$ר�%�T��ȃ��2O�y~�V� Gk�so9�x)i�l�`Js477G��%E�?�����"�c�b��B�^W4�����)��Cu����?@�|��\<���	R���V>/r=	��B��r����>�ķ�D�ƿY��"<������J6���ܦv�(K}F��1�7���X��1����B`�#��$����&}ҍ��C��EQ�c�7�\j������2�ڳج(�P��ሃ�r�j{C�هds�<EU9�K�;��
��@ ���e��C�C��qE��G�3�lA>�?/k>�&� ĩ@$�`��)^��jB����4�#��Ȱ>�;A��Wg���Ίp�}���%����D�5mD�œ��I1�k�+�⮸FY�T�9E�.���'C�-����{ ����$�q�{{����QĒ�L���?jnZk�.1��sqrغ5	�ށp\öF�-�l���[�������k:�әcV�X-m�����]�L��-��KwQ�_���ߡ��k�WD[6o��~���蟾�eQ
��V��r�$i9�.D�^�X��EY���E���ezff�*��Jv�lY���r�oS����<!�X��J�*!$�wvvN�]�tii)���a�ĕD����0�8VH�Jt�Wm�焑���h�4�ըT*I�H\<S�!%�T���[���^g�� �J�*a�Ύv�z�F/_���q\M��=R�⢑ɑc�����@��~��������3JFϳ�]/ުȉJ���&�4kf�\[sY���ڷ�������42;�����Б�2��=�P+����̕�tf�U��d��a�E�c7���-�`{>R��e�Bw;�4�E�~v;����jx�F��/��z�}(��� I4 E��N$!���d�?L�W��Y>��Μ�
_�7=��Mӂ4R6[Ak6*���e����ƛ��ωK�ib~FZ�$3*�֖B��<��w�^�m�d���q�-���%�~�ʫ��#���j*�2"��p{��z:�%>
4�8���0�g�Ev�1Y �[M�4wakZ���W�|/��a�9�
,l�(�MS'������"g��H��:=3M�JՊ�o��ņ6��l��x��D'm��|=�����w�]�|���|�M�&���*+���%�[�kb\9a�O�Z�Ξ�H�������@H�1�s��J��/�=���2ţ�U);���������HY��ZI���@bnjj����E��%~�1܆�i���b]�I�w�W%�2���E|S�HdF�5����FN.�[�}�R2�	4�㴃��dM+��t�"	L�%u���g��u���_�liH�s�<F��n�	�H���Z�H�bt��=��ۄ�9�"˾"����\�̷�~��.a����de�^�t�:�:�?7�u{���b��U��.;F��劬	�tVft��e*e�d��0� �H��a��\�O?�����#g�ҧ��9F�#�]Ń�I��@�]~������b�.���+�t֧��<=t�����CG^�G{�����=�aF0W苏|�Ν8B�6D{��!*�)1��)j�5e�������йK��{�1z�����a��P�U��$UL4�nPU{=���m���YȲ��o<��\�,n\��x8!tH� 	��
j���}�P��j�Y]��E���gh��dٵ�iaz�Z�iOh�2l|
mi�lU3T/{i�*��1���y�@B�!�)�V��Uih��1,��E:
�(!f�n���k�T:WRbp���,�$c���FM%�n��9O�Mܑ$���K�;;izq�EB����)���5���}�+ը6�0�5e����"�=Ny�x�V��ff�$�X�,��_��g���U��,��@���U��U:���F�./�C�A���X[V���LP��;P�J�\Vb�a2!�k�	%k��К/�,T���o K�l|	 hj�;I���6�"^+K��	\���#'6�� w�d{�gE2��7�S����I$��tk������Y~�2���!�$��:�h�������:N�����+aydz�M�����~���gP�d�4��j���&��r�����d#S���q��z�I�=�3W(@ɣ��mʜ�d��߲g�2b=76B�s��q�B����=[wЍ�����s�U��gw��F�;�Hj;�պg�>���}�����/��wʎ/3�i��jZѿ��m-NNS_����RT���?<E�
-U�Ȧ����Ѫ�����#@�\��mٸ�~�c���?�iz��aa�A����ϚH',�)��D�؞�������~��9���~�]�<x�9�z�*MMNҮ=;���z7=w�E��S��jP}�Њ����
-����ۤw�Zo
L���d�
�Lm��!�u�����`�+�[
���o�!��+Ֆ�I6���A����T4g�F��]�5�d�_.����Ң��2iZA<&��{5�*_�\����B,s5F@�Tú'h6m}��lJ���0q2�8�bZc��4Q���P��RBT�@I���vF:e�ReQ�QZ�ť��<�/�-�C�P��	�� @��:�MUH�3�HO��q*�\A�{p({�s�����@�������K2�)eP�/H�t{0H�Z�LLt�I��?�%�R.v�T.\Ʌ��QٰPIU������wwuu�g��o(��U�\�<��\'��O�/ƾ��Q�%F�9MC@P=T��� ֳZ-K�fݚ5R���y��!��]7w	�.b�?���kPp�#z_�)��[��M~�P��'�Uy7��WB-��{���8v��I� Ƒ3P�@�ϳ�
��@˨pp��u�\!
薍�����tvf�����HP�Ms�4]>��Ku�g�nZ�f��w-5�����E:>rF�N��
��v��E�z������AJ�b����,�yjϵ���G�5�^$#n�@�əI�D�,,#\�p����:f!��`:���&�Z�]<s�N��:�;:���(-�g���Z
kډ˷�i�4��׎���s2,�]�i���q/M�NK�pEo�$c�l�)(�+�=N�����C�b�g���fJ3�8r�K�75����A���I�H��(��������q�P����`E�=�b��S�L
���KM-z���4j��d��#>*��p�M)BXh�9/F�/��!J�ح[KzN���8�iO֋�$�(3�Ak%�Tm��.筕k� jAUX��J���P�l���u������]�Ps (���E���W�T>�=����$
W*k��%V�5�H1r��죫���kXI��>{��p4���h6n�Hݘ� %b�<��� �������3�����h��(a|M;�!E�6=��厭����S�x*W����]b� � C׮�g@��$���g2�Z�]�UeA9gBv���g����硣��Z�ҹ���ᗏ�kGߠ��yi��cxN��,K�����!�~zh���-� �t��HN���Y�{Yk�O�J6���3ZA`����~�'�����Ut#Eа4��P����w�TB(�4+,Lx�
b߳-U��AZݳR,��9V��_�����������H���?��ʌX�*+WLA}��O����Y*�����ҵ��TY��; ��y^����G��.�/��Ct����gT�AM�}��[A��}t��U�r�
��!y����h++.&������$_�A{n�Q�~�{���s�3�A�8dT�)�K�A�`5
�*�q`%���@�@m��B� �MS����׊�3�@���3�qW)qRQ��0��H=�L��CU,lP�$����K9�
F)�B˵�i>Z�Fs�*R[�XZdE1��ˈ���j-j��	U��`�Y�3��L�1�yi�,tRg['�g�*�E5>�9�X`ĺ�(dIP�*m$�2���lM+A���t�e��.��r�>`k���P�9	)tS��.XX�p�
$�KK%�g�����EA��|J���(���tG�,{��n�̗
��]��:��$ˆeÆu����;J˺X�֬^KWǮѣ�>�����i�3H���l)(a2H`�`��T$�r:0@�}ǃ�}�.*�A�de���|zv��響D�?�(I�Wm�i�(��M�տ�fˈ���s8��Kw�~mڼ��Bz1�����jz��'����VĘ�V���Gh��z��%�T�Z @b�/��J�U��;
�a�0��iO� ��, @?qL�9��C��q���"�tw�ʕ+���st��ـ���3��J"������,=z���
����"����`���S�W�䌯�]H�!6QF�$����}qךvD�|��'���1b,��i����j��iF���=\�*�Y�����������-�Ⱥ/�*��K閛n�m�����_��G�V*�{_�D�ͬ'٪J�7n튕���a�[����'>l�8ܽ��v����^)���E�IR$�l����[��M����\��k7��{���������䨄e���]��#�F[7naŗ�J�{︓nݳG�BŎn������/�+�����f>4?x�j0�;>Q���3��Y� �<��R�d⥯9,� ����|'��l�!b��W٣(t%���EQ̤�i�4'D��ٖ��~�и��ĹC���Vx��aQ�ˊ������-�R�=���z����5r�*/I#>/��T�#i!�5-) �a$xq�Ps8�p�P:�ʽ����:�ge��9F0H�Ayud���e�����99�Fh�F�-,I�Fdrq�=��N���<躹|�|�@�b6O+zih��Μ9E'��u�6�:V��lN�P��ף�
�(枻���ZR]B��l,S��F,Ӧ趱}���* �!,��o���MFfWzA��)��pmtY��$ה�)�z�?3�G�t�,]�2B��>ڵ{/ߋ�[�C�4��>3jR�p���>��(��Gmʹ-�3�E{������3��HL}x�zj+,���R�m�aD�L8��N�#۶m�[o��C�/�֍8o��mķ����	h#�_m�+�8a�%sv�&���+�%�GS_�r�2Ȧ�ti	��dLqZܸ������yC�k(�揘����j�2v����c4��Rb��7�8U���'��X�ɩ@C���]�@���/�Co}��s�.�*��@�s�~�zZ�q�%�R.�o=��w���t���t��yAyvIR�2Q \������v��DL�����Cb}�r��z�^�e���Ї�i*�"Aa�'Sa�/)_`e'
+%ɊJ�L���vVJM�W�xh���kSVz�u��{��B]n\��A̲!B��;ug�i����}�v�A=�bY���a)�G�qٮ�N9��ᬏ^�+Z���[Cjv�Z	��sB�~�6(Z��,+�T����M붳��*���k�� eQ0��+� �|�ϓ�{��g������օ��?&ٛ,4(X ـ10u��]=Td��I�U66��::�exn�u�cř��[hα��d������'0yee)ڔ6Oı�:��ћ�G�.�C{��Ì��ep$���y�#��HIg[�,�m��������5\�c4Ti��Ƣ��cŊ4Z+�+WӾ[����/���F��h�T�B�è��Z�E݅���3�Kp��4�P�[�n��6JXb۶͔����cc�)Έ�������xi�8E�(��K1)��+0F����B��	�:�h�?����N�9'���u�ʡڸe3�|�(F5"��n-��	=��G��d�����n�nȩ�	ѭp���ɚ�%��;GN�&��/$������~��ʭD�C����E&ʓ�й������T�3��G2FU|�u}4ؾ�s�t��}����!,p�x�v߰K6;ǖbz�.]�H�@g�d�:��}w�6v�^c����y��0ɇ,�ʠH���ܸG�U��η����zz{e���w1�M�s�^�V΍k�Q�X���Iz�����ht�Ʈ�JI�葬B�K0:z����������s����H�S5����r��-�vӽ��U����+W���E5z��hߦhM�0sE�!Fna�,�����Q!��M��|��5����+�`�$:�4��d��|�r��|��D�j��eiYp �B����C�L_��*���"Ji*BآY��V�����n�ca�1��W�Y��k�7�o$8�]��;��gŝ��ncd�{��40����(�^���iAM��<���1f�tSb���dI`�5Y�$�TW����ƶ�=��7�B�cT�MgΝ���I��J� �n��K�\0Z�Sz�A�ꍡ���E6�i����)0K�i�\ 	=����w�x���c�c��܋�D��h�P[�!�0��=�c�6�T��G��\�H4�A��5\�n#=�wЩ'ip�0�^G����C^���2*��c�A�W*����:4�k��v:[���{�n�e���_{��]����wӉ�ߠ��9�,�)p�2�'c���$c��:P/�����lg������?Hӓ�ȧ�l������ec
H��Q^\�E�$�ڡF;���^����ƹ*� ed�k����һ�K
T�j��5�8�����z���֙�B!���-F�L�$ϼB��Z1����-7���W����I�b��ʚ�az�;�F{7n�Lu���3�@m��ڴc�L�2C��M7��vH����Aн�.��w�U�ȵ+t�}�R/#/��t��4�ɂ�g��M�L��|���M"(�Y*슭^1(�pt�*}�K_����Z���J:m�ő�ͺ�dNC�>�u�H���Y���b�P�Ic�^&�S�����_����ZO���&V��]��=��ĉ��q� ���oY�f�FJ�h�Ua���@������;�@�|
��і&�������7NPOw/��u*JS@M�����Y]�x��o�@w�yy/��3KҜ�%ܧ�1�D�[��,{���C7�t;]�0&q?d�ڂ�G�C��@Ə[,q`$M�
�Tg�B�4����܄O��!i�^�r��}/˨���Y�hx�J���9MƦ��l�5.�������9v1Y�c��Q@�~��"�x&j��}G�	Q����K�#�QF��.]��a_\���qV�Z+��:�Zo��N&�z��0�H�%9��}�粒�y:w��`��u���V�g��\�jM}�pAs�P��+����G'O����+�y�� �����{��6&��^��R9Fd��֑��gH^ˡk�5������I%eZ��._�̊�j�Y�{ۭԱb� V$8����h��8<LT�ke�~��lB������&LC�ջ!��ODB�s�#U���tkً�+p�%�O�Z��%�ب��%�B��!e�"�a!])���ѣ��y&�NeVNSS����� ���|N�b:���=��'��%�D���2z�z:{Ey��8�Px�rh��ؿ�^;v�k^�yxh�XSl�4������G���w��.���s��.H����u��� ���?�퀘����-[���+ƔTMDWr�C�f�umf\�Y������V����vq�I\�����+"�87�q�qj �^����Ȳ�PH�~����>�aA#X-Ui��mt���h`� mۺ��\�L3�3�Mj����!�}��A���i��@���	���J��-͠8����}w2�������%jgc�Ni)��⒒�kR�.m[!Gs�����۰�d3�Ș�1gK+0�y��jʱ�ݰ~�^����e��JVBu�u�PJ��_����N�?>?C�|J2�PySId��qW��HdK�|Q�{��%��0��U���}��4�T�2t��3i%�A�G�Ѣ9�G���EO�W�,�K���}���Q�&B2>5K+�n������H|\4����Z.씇�X�G��gX�_��(�� ����[��9M�I�/Fy:�Ht����YvM�rN���Xy<P�����0�D\���+�G�Ǵ�k�ͤ����[���S�$$��^뺵���ٳ��$>�`|�Q�Ȁ^�4�z�ҡԥ�~��kE��T�3�����U��~�0�I%����T��~Zk�,��u�a������QĈ���'_��l�R�4�ZK���ibb��z�IFx��{�b�}��oѓ�>EC����q7�_���\�FϿ|�Ό���ӣtv�mZG���C{w�(�1�l����w�;��Ni9պψ��N-Z7�ڼi3�ټI�	mZ��Q��t�[�@�]Fn�B������q��)�]S�D�q���dU��6��$V07o���x�=�d�:u�5��F�z��I�ڋ.�I�q3�#e�' 锶dH�,�1nu�ٶy'�H:�:�K��j_�LM
�Y(ω�g{�b��v�1ft8�0/��☞Yl� iGI�ĳ�t��oc�� <�({Tbc#�T�h�l�����+�SJ�a߾�S��Ǥd���*��w��b��W���iFSq��F��\���P��G�-�����S�"�3��6BpS����J�q8J�	�*��m����]�x)��x�����פ.8F@�
�r����J#��ZI�6G�ixZ�������<F�7s����]���ZiG@�,�Jv��gi��I8�@��
�������''�^��#��G�x�e�-���M3���n�iF���qn���Mi���Ƒ���_�EF�#�Fs��]clH^?y��g #��ޗ�{@π?��{$>o��V+�(��N�eJӶ��hɕv%T��,��ŗx(�t��� �;3~�^��]�5�6� |]:��-��WʡR~��̚��*4�h����@�I��u�#I��z���G�����볇��޹}m߼����U�XN�%}��y���ct��qF>s�u#+��n�tYF�e��骺&YV^���m�[��������x�}t��	~}=n��=����OI��.v�ׯ[/��ݗ�җ����o����z�L#�77��?�Q.���mUlWA�|��
�G�5uH�/O��%~���r���1��������h��*g�r,�Y��6l��n����I�Z9D��t����2i�z��ieq���S��**��Ŷ)��LX"#wnɥŕ�ǃ}��&��������������
uw�y+#���������MC�F�����"�/��~.�@�{��&������2}m�:���/ʤU)�j���%Y?�R�&]LQ��o^��؋,{H�6M�&���Xc��!��t�	YF�$�C�gF'�P!�8w��F�׺��?'��@�3�p��6�[ʷ�_/�XյDL]����D�!�����R8��C��@z`�M7���)R�t���< ����kTp�_�#�(vժU�|%Z�n�(���I�<�%�y���g�1�3#�G�<�RGq����<$={���A�)t����r&�Ktu]c�T�T&�z��B��Z��uww�ɖ-���uh��n4-�d�@��}���8$@-��&�~�9^;+�x^�=.Q�7��	�� Z�CuYŝ��2$Yv�}r,H��.j��zعe�q�)�B�V���(F�Sݾa#����i��Z���i��(��wi�[�M�j�{�H����t��X)����d�+=u�$�6�Y/�����=���+� ��s����6��0b�%7���ei!$���ZY6$-:cu��6/ Ȏ�ڡ��~�z%��-=s�J֭[�®�K�Xp�!>�N��gea���e�JWT��⺶8]5Yb�XCt %�HF�K��V���/-B��PUif�-<�������yM����!�����Aj�i���u��	�)�f�i^�-�:���y���3P�-7�Ȯ�4��^��+r"��{έ֮��P��p��qC���$�P�����f����U+��\�F(�fV��T�9�ٓ�k��"���:*�+R�	�X���Q�3[�)����7��<����.�Š(^��D�_Gg�V�����pq�r@�� er��F1kj?q?0�7 �<��:�����`��#%��!.�7�kB�a�w3QK./X)Q�%��*�l�l���b��c�ע�ó�2U;%+�2�H;�7f��`m���h�e��`4���R�z����	�:&kh�$l��L�e���C�F)>'NY.Ӗ��r��<�K���}���_V�T�[/�/�%5��\?�V�^�T��dk�xd��#Dq0�:+�|�S;����������#i�S������s��-ed�s������� �D�������g�+S��&|�7[�� �̧�����+_����ӎ��Y��%v�+�լx׭Y'(���z����t}I'�*��v�D���+�x��>�P�1"3�Y W�YC���>��\cŔ�τb�b�Z��~���r�سtߝ�Rg��p"�n���k��w��|�߿?�aik�q�6u�z���l�+s�4�8#n�� �@:�Z��K��h�d�6�/�j��1�
��ꤳ�O�!Y�r4,d����GYW+�S��h`�z��g��[�GD��WK�B�	֌�R0%�;�������uvt�K�!"!����VR�~X�� 0:��A���*�Zdr
4���(��A.���݌SgG�	1�ڇ�~���"P��|T`/�-Sr7�ċY�--��:��;�)��vV�m�LaP�@��P���L�NQ�3M�֮c�pR�8D@�0`�gg�]+�,�,\Qڏ�o$	��_��x�C�y7��Ƙ�Pgg���ڠ�  �.�׃��5�O�to�J�w��If5ߌ�J�(h2����鬆�7�4�b��gQE�J?���R�A�Hs�k�c'�o��m� ��\A�qo!^g��ڵqA�)/#M*Pl~]kۨ��sr=!�A�5�&����B
��i)Mj�]�'%�ӳ3ˋ�+Y�'���bႋ�S(��)]:H�s]��ѩ�atӖ�3+Ѡ�E?}�h��m�T������_|��آwv�k���`O?}�g?B[7n�����÷�N���4�(Q�5h��镨������a��[��`S�y�)������w짅�����~s�t��̭��FjLafSZ*�ĝ�5f\4�T*Ǯ=8S��7�7�Ͽ�yz��giú���~V���}#��8=;�m��	e������jIbPh�DA������Ff&�?���B#S�dIvA�6l��U�I�i��^/�љ�g�T[���k�rr�Va@H�� �)�𚍬 �i��#�Q�G_�&fY��0��F;�|���䙓43;I�C(&�u;]�L�.]��=�h� �q��t{�C{��Ez�T�U�4�s��Al���]�����v��6X֐/��^H�hR����ԡբbJ5�6j1���h?�(Hŭ�u�P��%*���W��% ���1�E����e�,9�,���ϕ�U�| @�h���j�H���������k�V��&vC���x.g���`� �@��k����_f�s� ��X��W��|�5�{.Rw@Y��	�����ͤrٽ0�F�prQ�0gkB.`@�n'��P����u
������=�,�g�zap��'���6V+����R��}ȩd.���k��:��3
n$��4L0f��`:��6�Ă}�s����Ŕ��c�?C�c�����f��yp.5��v��4���GC}��m���sg�F��}���xvq�(���)ٲ���e/a�xa����{%���AiN�+�������&�>�B�8]��u�`�Q�� �?���#��(Q��>�i��?��jT����?ȝ�;־9�K������Zf읝u����/�k?��D��E==����~��4'�!�X�rO�������i�/�+W�o��r�i�^���r{���Z[�'�Y��'&e����F��o���t4*x��g�>�yn������*�~F>��g���~zaNN;.�x����K���?�y�vv��/�X�z�)9�����ǎ������{�-���������X�܄����˼�fcJ�3��o� 3�!� `��(�z����e]bOí]y��/䱓ʚ:5D��+qMJW�]V�pN?�%>�����ݸw[n��k�l�n����PK+�md�2��d'��śo�?��}����2�A{���i���LO͒]1��-I}l��16d��cW`���;j�FNJhԃԞ5�Ib}}[^}�u��(8$�-���s����Y�[r��-�4�pu��'����iG�=�]݈[{ۜ�}_:fhGM^+� �%��(Vy�(��U�קgʪN���8��^[��=�PÐ=�:�bt���Ť(ɥ�C4��Ύa���� ��Ľ��G>�x����n߲I/ޢ�9�Ǭk�����1 �m�|����<s@)��}�/�:����t�D�;>S�7f��\��D]�`NN��N����5R$Ō<#�� �7��f�3:\4��2�nNXg���ly�Iihf����#�yo�Es�0qkFt�5k ȭS�;0qO�K@�4�f#~�y(v%<H���Ɔ,*)_^0>��mUO�~^-�cP���|��iT�[����7��_~�k��w_�9}�O<��|�����(��9�4{��e���U���J<� �������q��/|Y���/P�K�|�I9��������eW���Ԍ���0Z<�Hx��kD��D#�6�핋��o��yt���G:DNjZ���>��ћ7nȷ���|_C^z�ġ���/e��Q9s�Lkڳp���t��{z��;w���?��ɟ��,/�p_�{�~ ~�q�X�(VQ,�y=w��A�x��]��)�0��,An�[�#ib�&���ɩ~�p`�"�E�"�;qR�:���dXY��u[�O^~I.jd���AcJҨ���exf.mc��f_��A9�xB���V�g	��A���1&��9#��l˝����ޖtG}��2��!�@��i U���_|E~���D�>Z����ut����9wJ���i�%�Ԫ��yjB0=����z�*���9������U+� q)|R}p1Gj�{����2,"Mf�����m��iۀ1�qDf���{�ZcD^Ү����M�9ůn�וØ���#����r51*���ܑ�*���uody���-|�!s%���g�߃F���f�n��bF90ˈ˖�,4>��	,���x����fA�o�b6���m���L!Ѝ�M�����\>��Ž-0:o���b�69	��j��+�����W!#�.�jČ���n޾�8��ޖ���w��������y������H�j�����=yᕟ��kD��wߔx���k-�z̖��+�����/���8tL uA�vlr�KH�}�#�G�?J������4��M�����2;13)�n]�����dS���ξ���(,�2����KG#�4��-'N�/�֗dcc�3�`���>�i�0xKs�����_��Ώ��w.\�?�������E��tt[#�_E��ޖ�����	��4;3-�����Lit���>%o\�1Дpɂ:�Vݦ�ư�{x�m5�w������3�� �a�51�����FG{�;������~7��//^�W/�.��[���;/L@s�~Q�dA�J,�C�����������������rg8�Y7��~� �ÈD��Zo��.W7o�Sڗ�~�Z
�G�� l���ʢF�C�w$����^�S��ж7��O~B�Ј�;G�� �����c
e^tom���>���h����m�X"��zN7��1"�E�%*�"
3N�=�����+8�[Y�U`t��\�U�KZՕ� ���L��E�:�0@��k6|���X��1 :)�?��<4X�kF:��XmUTFF�11NE���,�Q[V��o�?(o����Ƶ�G{��T�?q,�� A�� �>�i���ڃ�z�8�Mא��/o<�]E�%�o������p^�ܠ?)^Ʌ�����ޕ�W�it��B���%9�FX&FnC���Ʀ���{���'�]������L��x�3r�0��xP#�����+?}��?��<t�,�N,-��<��Ú
�jzPCڃ��_�җ�QN�ɱ���[�{^6ww� zWފ��#�ֹ}�tzMu�eiaQ����4�M������`d1	uqeY^��\��.��[�4�%j� e��򅟽$���w%�h�A;����'[���@3a
]o�m�L��)4���quL�����j## ��h�+�}��:TfzES�7oʇ�?)s����>�����<��	������r�����*���h�����\Y׃�јA`eoؖ[������|����h��Ʈu�hd�xt��X�]����X�ْ-��!���Qe�o�)�[p����=��kwoSUϽ��e�`��cl�)w�3�u�Miv~��uj�v@3B!$����;����!zB�9$&����nU��eB��!j�Yc�>������ ��)#�`d���
��Q0���(��7������+b�2�nm�
M�j5<���`<��Vª��pRo����&~��Il㰫U��5�����"��s¹���9����bi��<�e�q��LR�߽B,%u+��m	�v���?�}�l�hm�?��%�@��:���`��D�E
f_7���Y���&yᵟɛ�ޒ��C�S`G�9�F ����D�k���?��<��g�-M1��O��ܽ�/ȭ{7�|�srr��)�B�aQ�B[JT��~�׾񷲹��)b<`� ��歛��W^�/~�T�M4Wш���^mo�4ܑ��Y�h���An<�:�H�'/���>P���D;����Jf&��X.K-1��wo��?�>����Q:��Fd;VDql�E����i���kt�E$�����;rR#�SjȆr񝷸�65E�v��eM�w8�g�ז��8ڣV�K���z�I��RΖT`�}=��n[��|�|wKN����4�[����F]F6��<�@��Ձ�afQ8u�<C_�h�s�i�v�/�z��62���Nա/�-�-s��1K�"�;벩N�n����N	ƀ��g�#s(y�<��`d��`h��ĝQ�<���RH�?'�4��kl|��%B�Vx����Jڎ�n�P>�mں�v���]�b��I0@{���iԇ���(5v
ƺsj�v5��>�D����o1�{�k��ќ���0:d���,M5������?����c�:��Nj��|q�y��+#+�_��\���1
?�_�
�)Ӈ
�&�	ĥpϡf�0�7	C��a�R��P�r��saf�8*($��������7���+r��-n���=�`m5�L�"��pzn�]�QA ���@c̿�˿�_��U��vW�ݣ=0�������/_�f�����SS��H����bA����o�!��祗vY����`p|{�Q�GG��|�k��P䛝R֨��x�L/����;lnh�1ISC�N�/�\�D�������\�{���P���p/���l�[
Gs
����[a޹Ή����6�ۤ�!���]�f}*�G��i_�����r��M��k@����u�#�mȶF�=u�<5�Xp���CDc1y1�XI.m���4�;�i}��1����h��� J��3x���,%�4�֨/v�K�Ѓx�+��7�g� ��J���^e x�����;�(�/�	��ԫę�V��E�b�fG١��u��i������Ch��v��4�-5��S�@?�v�:;���a0.�(V�7k%����+,u%0��"��X%T߀�nll�����{������
F�zb�`�0�Y
Xx�p7;?����v�K#��nĴ��Y$?��s��^�K@��܍�A��P�y
�i��N,�.]��~&+"�P3���%�=�B��x��ь����e�It8����yZb�H���!	��_��o�U]Xo^�@�<�Tu��n\#�3�+��-y�Ƨ�C��h-np�>2�(�AD�=C179-��{���_"}o���Q�>�ۧ��`�G�I���S�~�]����^����XT�^���Q����Ct�bA8+[[m��˨��oٰ94gd9!��.�-5 {zN8�Cg�����2��F�~6���C]����8����F��S�O���۱	y���d��G�n�
^���H��Y���Gy�d��"5�]�ޒW~���w�2�<�b�$*�8x򦳐�x�Ʀ�g�"(d\e���������e~a�Ɯ@[A��� �-�d��ikQ�Ь���	�=W�tHU�ڍ9\�U����L/ȑ�#�`5�>~�FqscS����\B����HM(��#�H��)7��@�WNR�R�yv�2B8���Q-Dc?_�����f�k``�R�U��q�GgTu@R�z�znݺ#u:��&�ԬS:��&}q�ڵ�\��;G�
La��,8�áUE� �������dFg��2���}�)뀔C�W5z��z��
N����ZBfF�k��hϝ���ڈ��h�^��ӫP��1�͚��M>3���#�f|q�V >6��]c�45lЧ�����1LT2��h���q�B:N���Ԛ
�n��QĞ�:��RnTp%)(��A��A��Ц洊�.4gu5�F@����Q9�	�,=�t��c�7�`q�S舸)�gL@������� uW'_Z�Uss�O��}Cjw�����*�z��������d;lxzO?��<���!��?6'Z&��_V$�e4�
CI����MXڟ��/�@��{:�e=6
����XwO�����3�xn�|�ETSc�.6!0=�ZQ� ukӵT�(���=���¨Pr/���88�}�8���� Ml2-��&x�0bh��ϔΛi��~�/�z��P&��/8�z�?�ey�g/{/��}�ӻ����k�U�����&��aM������M�[7k�J����"qa�J�9Z��n8�Țdp���E��m�0��
�l0s	]d���Kr��r����� ~8$��l��{T����#�e��2[�fK!;0�����nL3/��خ<AN4��'�S��ȑ��r�}�A���Ꭲ�'�V_����?M��W�+�l�SCk8�zq!
Sl�P>�Brad[zfS�	���'Lk�3�i�R{���9:�k$2Do]b�Nyh���:�+�01qȽ�1O}�r��q R�BF�	gDM�	%K�I�� �4�f:���ޔU�$�+�3��b��~^��
��v����։A��7�?�L�����!Ҿ &'���D�Mr��f��`t�+3���n9?ߔy�ϛ�=4W�87��(��S�B�Ѕ�9Y�]��lL����yu�j��]Xa�Pj-���Y�
�P�I5��rlqQ��%y@��ނ����c���ܙ���"�kX#�[a�h��V�|�y��0&+KGx�����	���d� ߈�X��v��ի6�;�bWج�NIY�:��i �3Z�����Mg�3(np �G4&Rd�mm�tj9;���K�_�0�U�I��1L��b'D�A����<��2��A�?�g7�����Ufi�����֊��!à"�^2�� {Ma\'"ϕ��)p��~��s��F9� �����1h��%֔�I'z�y��']�R��qt�m�c��l����F/�Qbûm=�y��Eݞ�/8P)UƨM0V/aؖ6u����3=���t��J$�E�n0� (R����W�\�"������%+��KR�]F�R��CRcda*����y����J7�,��~�43P=�>x��anS۔�����^D��㨦>ar*S���3
�gi�e�q*h8���n-���r�9q�8.�y�g���w�D�*}���^�U��
"x�F>�� v�Ԭ�o:�ዑ��������K0>�}J�3�v�����q3�)��cæ��d��0���i�ϲ��5�jj���2�i7���7��c!�2<KF}x.����>�Q\�E�g�O��xr=F-�}�c�,*���{���B~nqA�=���om2s��4)W�2EE����XQޓbE%�ƑC�� �7Ի��c�NZ�X׸�q��=�bc&	
:���оXL�̟F�S�3�_keA &v9Γ���\���V�����o�k��)�V|�116�b�*���w��N5c$�}�1�$�#�=v\�Jd15+d�.щ���([��wS�/5RtONZ�E��,0WZ`�����=���f��O>!��?�F<W:��I:�'�.���s8�-1ּ,VER��_���.d R�Y�_)��rU��d�^�2�=p�V� �]�&�2�o��'��o�Lk�xV��б�Ad���91�χ��(Ja�	ɈR��a!`�����gs����7�+)9���DE,Ǫ�maa����B:���(/),��[�/�{Û��ϲ3�CO<I	�W_yE._���ˁzq,V.v�)u5�)b#�6ı�����$q�iXX�np QE7K١���2�h���Jr6��A���$|i:��P���A!%�M'�s�+2��s�,8T�9�����@ �W�I�6ǐ1XG"+�e
]�kdjz�)6�Al��^DK8&��iq|=8n����z�1�@���EQ*D��^�x(�ܾs[:�:M�Z�qHk���/���"���&�BB1(]G?y�dQ³���y�h�8���~g���8\7�k�9,�{��ﭮ�������Y��h�?h��W��0CKvl�a-�ߞ���3�w���g ����P`øw8����,�(�>Ϝk�ȡ)|�Oq��N������轳1=�Ԇ`L/1q�	~��h���\�zK�٥�b�@G��"[�g��_�l-.	��Ǵ�X��f����WT��P, �($ȥ�-0�P7���W)��5�I�2��͝�����t�I�u���E��P�YZ��zt��y ����1UJ���K���R�wd_d����^��.��<\&a�ԅW�yU�$�W:�@��V`�s�b���F����{�«\t�(�kpZ7L�����9>ex �I�Y0�5�%X��+K_��%s�b��+���G���=	F��{��"kKkBk��a���Q�&��8�=��Q���;����&D���-��9�iT�.Efӧs��[���F�����γR�9<@?AGT�`�K,*�dsy����+�����X�"!�`�?k��_��p(E���!�=T�= �(9<�]���,�q䟙��&@si��fdG�a�5����5F��F�z���<���2<û���<��-3����S���5u�8p��a�6�(j���� 5�@�b)����Pg@�B��]�
6�v�>� ��� ���wYL!�3�ya_U#�~X�[ח�>��-�> ���Q�}߀\*�����߱�h�ۨ��:�V�2S�
��h�M`���p臇���Q���Az�B6V��i�{N�u-�O�"��`cw����V� �P�P2�f��qj�ׄ�HX���P$;2,l��:��~�7����s�L[A���������
7bE�'ǌ/���E��q�Y��F�Z�r�xq�U"��:�@y��!��8{��>>�Rh%T��ޅ_�f��KpV��8���� ]���/~.i0�I�=�>�1�ynh=�#�.��l�` P�P��իϩ����6�]o�K��D��>�#���������](и��|�I�P�"�ic�����F9����Q �ila�bMΊ-�)������׭l8d��eri1u#r�K}�Rl��k���;�K����Ш�nL�(! ������]#]GA��S������u���/֯/�qp�(�q�/�Ϊ�&4�Af$}�"(��|��[a��n��۔YQ|��?/e4k]��,w�SV��fF4�F���?J�@C��HOV��Do�q�ho��U���~@��P����`�Gji���i���*xFXlY�Z�YP��h��c�\@>� ����b*<(��G@eA4w�y^;��BQ�vg�_`�v�c��P���Ƈn��%��Kadb74Z	����Z���a��*X#�n���XЎ�k��NUXd�a�݇�@)��7u@����fg}H�9Unh0ĉF�+ʃ�0�����0�l������g~�+�jl8�\
0{�`>ҩ�����"-�W
�!���>V���#8|#�/��8~��Wׯ��+�SdMA�$K8����H*8��?���]����;��̘�(W�����yU.�\������C���5�Q���DG!�y��,-(L��{=C�R���y�e����2&D�-���٤�����U)��e��!F�`� �����K�6���+�X�%Y�kF�A#T�:L�[���,"�Zg(�Ǘ�=�99}���u�+��{��|����ѹer�Ձ���E4|Ǧ����#�v�x��^Vyx�J,�Y�O����8��c��5�/f�����ǚ[]Y �" u�v��g��>������C�N?�oPɃ��a��&c���1s����qQ�w�})�G�a��_E�WŔ>�Ž���V#�<	Wj!��QT �v�JJOu�e�1e�B������wE�rAD��±�J�z�����zE�Пn�]y�,;<�ᐅ�|f��Ի`�;E�L�3�F�{�\�F/�����k��R0�"�+���{�_��Wx/���M�����~�^Hˣ�7
G"�*,R�)qQ��֗ ��s��eG���N��G�f��5Fiώ�Ʀ� ��u��Ʌ���7`>!���MTM���Ź��������}�:t��HV7�DV��~���3���MK���h�+�iM>������O���j�Fi1��{[����_�l�aY�kZ�G�$�ȧ��Ġ��Q���/c�C���)��NL_]l�J��U�ٗ���Aϊ;�Xq�Ām<g���(G=KumH3p��.,x�|��5ٸ ;�S�x�<}�Ԉ���ۓ���s�N�3-K�����
�m�(�`�����<�.�`i�O0�"�޿�������y��"b�����c�����I�Y
%����}1�y�u�+*�Ai�}N� #�.׹T��ǈ���#�/����?h��U ��4� c� ����9�p�p=v������>�u��7�x���?��+���Q�'Q^w8����_cg#R��j{l�~a����5��Z������`��"7��ퟔ�-=B�4�٠�8b�V㠞����Ϯ�H���C��'܎ʽ(x����Y`\�]ǌ�5�G.�l��e.��+�Dk�k��/^���Y�mY�<���30#Yc��=�^�����cm(�ٌ� *ai�X7+~?����>��c�_�}�mL���˭�-y�ŗ�n�61�?�!����2+���A�Q 6*Ԩ,#�E��KYH�PA�t���.�:�!���7�Zbk~G�^gό��<#��'5��.èXQ�uV}�Ԡ�8��R�
��|��&����n���K�tL��Fr~^(�DN=C���v�&4'ȡ�ң�pm��e�܉�{�ؔ�p?�uƫ���~���%v�ZTГ�a�C�3�x�ϫ�v��x�V<�F�__�Y�S;�z�wf����G��u%���͋�8;�"h1��ᕆ�za,*�zA�����*"��Ǖ��7�.C�f����\�ቑy�-�(>����XDn��(�z16��}���d���B�W�rýF�%Q茲�<��B��H��`l��fՔP�2��>)�E�1fc	�$5ÚJطISE~�a�� �uWش����e'N��^C�6W;X�ׅ?O�Dk��I۝m�|�=�C5:��ȁ��S0. �ד&���'Ɯ��[bQ9�D?���9ε��~���}��Ҍ�����j{mG��\��iY�]��=�Q��ռ=De��XP��ַd����~��t��?D�
6���Ɔ���+b�C�������oiT
(HE�#Da�G����4rSu�v���-&�ʆ����]e =s�T�kSb�>
�[>�D*QZ��[��(�mA�e���JfxVX�_.WRRҒ�q�oߢlaĝefг�������L�.>���;"��b�v+���rhRv]�uR��=Ø3ܫ�T��}ܣA_�Q�:� Q�g�N+؆��d��43/Gg�ّ�s�eV�gJ�(���ܠ�
%A���=#���!�`�b\���+D��2h�e�`ȷ����$�88����Oa37�Q�|x�Bfъʄ���%��GΣs���b����f�k��Cv����0Q+h�]B7#���G膀#�
c���	aB��Z�BC�fC�&�k�L�`'�F&��۟�P�q�$0'��b�v��ϊC0�Q��n+�,DO��bL3q�n�*��=AЦ0����|�mzH��3ͼG�Sy���{Ɇ�!E!�C�|�6/�c?���!�L�SKX��ɋ?����r����:��VWWess��$C��7ސ�'1�o�}�-��/���7����^KǕJZq��<����7%�"�Q�2��Hģ�������Y�d%�	�lH{�k�V��O�E��)3��I�0nF("O�a�����p�8|ߋ9�Y��|��x�x�)�H�f�e)$���oݾM�0��0׭�V`�����E�7�ua���\�1J,�a�&�"�6����klۅӡa�I�7	�_�!�
W�`�[�y1���4��݂u3&Q�h���>�-6��� ��!�ϩ��Թ�s/���.��ch�	�zT�E��y��ƚS�� �R��b3�pn�g,��C���(�N@�Qd��'-0���c����>�a4g{�`���˽�-�X���MY'ր㈍1xp�l�l��6���V*^����w6edĊ�#�I�����
q-����޲'в̕��t�]+	Ye�"�׽n�S\��f�W���t3� ��P���ۘ3����'���zë�y�	��Ȼ�r
�r����k�Z��,@+$T��Ŷ���������{T���F�@"�W�pL&�^�|�pպ��wl<D�0ܯ�����:M��0&t�=z��i4s�!��i݆�~��	���c�����3�2�FDBt�i��&�e�_�z���'�4̋<�|���"�3cj�f�&e�_O}���{�Ř�~�ǹe��˧N��̜\�r���K'����������ʓO����U��7Ǭ1F*?M����h��::}ꔬ��q������/_}�z^�gayY�t��ؐ:t����{�R|p�p�(8�>���ѣ�l�����f3���.��/ǧƍ��� l��vf~��f_���އ��D���(�-��ܪ�� ��Y`Mmjo�)�z=8� ��g!�y�U�d�nJfC���.�ދ1�p���e�����H����_�/pW������1�7�$Χ�BH�xo��]�?�qO�>-Sz�߸Ό2n�E��0�(;(]l�=��gն��q����G���6\{id�$�9�&^�C���z�������1"15���x��`�7r'��h��e5��0�l�SD޹ukJ�Z�'V��"v�"k�Eu:�>�ɧr�9లx)c��ӏ<.��?���>z�7���#�j���y�v�F�ZP��Ȏ�O��E���h��Ѣ�E�7pumU����˽�w���1�͂�t�:"�+�� Z%��с���E�	��[N�l5� ���A�!�8�L5'd02�cE�+V6D���n������%��e0��Ji��p�@T�(�}��Rl�/�V����ԛ��3�kM��Y�K�&��e���۷�G,���o���5F�h��\�T#��/��w�~�Ϣ��Ae*��s�-��x<������pc����;�dwkWV��x	�w�dws�	9�ܫ��� y䚫z=��^o�Rڀ�O�4L5��j ��ta1+Nn��pi�-���@�6u� Fg"�� ��c�|\ڕ�e�����}����C����y#�O�U7M��<���D��;�Z������ys�Vl���N����.�[��~
�f@h�ث���S��!�-��:.p_�������4�C��[4��k�5���K݆&FK�8"��?�h�X
ʧu�R�F\#;!��E[��έ���,+tw��YBC�Sf�>� 	��)9A�юOP
F�~�[��桺MA�����1գѨ1�^���dlrB&������v[>}���{B>�̳�y�x�P��%�H�b�4k�⫤��̋��"���M�f�K$��i�ڌ����bFPj)jU���60��~�/� 0	k�WJ�T���\D-
� th�jiŞ�o[-^vU^.��m/]����Òu.��!�U݀ [��Z�'q�~��Iy�̃��O^�FL'��܋T�s6c�i� G
�2�Xe�G�Ko���u��ZD#��ܙ��ǔ\8N��w��e[6$�~f�
k!��;��׶FM���b�țY�VW�k&L ㋬ѬFs+A�֨�)DC+��(��Z��-΁]xA`�שa�9I���%�^�ӈ����x.l��x`Q`�q촰��0`h��b�`X��a-��o�܋x0�Y(�lvK�i��.h�ah�a���ʵ�*|���(�bPU��Ygɠ<O;��u=u���4~X-����o8��y���N���9��PH��Eu�Q��"|���·���=�C�$���Q	���HL<a�0B�8W>��A{o�dL����P�f��l��~?�K�/�Ï<"��K���Y�Ih<Ѱp����w���\x�$AF/PB�(,��}�xE.����{���t{�_��7orq C�&�9��)p�A�@㢯P����e��ך�MS��8�1�b���e�1,y�5s����]�I��Pڋ�a�J%@?��O38v�!�?�z
��C���x����Ao��S]e�H�%��WF���Z{d���P��uDqnD���U�^inϡ歙��(z��þoD�T�%����:��m��[I�.��A�46�h������	[�5�d���Ho3j��2I?o�f1�#�q����4N�����TW�]U)�Š�Q�R<���giɇ.��,;���x���Wp�YFq|�e�l���70Y�r�ǜ{i�B�ru���X�YD0j�#M]H��J�9�[`�Q�Q-/拱����zd���P ,T�l��<���ז���D�����`0��1�a�Dds�v�jX�"6M���`x���f/-�lmL�f��ڽ#��o���/�cKg��1�H�a�����K���^�[�-���^oW��i�j�-BOx��7�f�H��()��fR��o��?~A�����ߩD�� ёD�nH�������Cou0)d�2h�s���FHӚ
ﰝ�"㩦:pa�k^��7���U1�a	���*+�G����L�>^�G�#�_o8�I
�1�����B�4:��l��a�}b$ys|�p)�"$R�a�FgA)AM'[����ҭf=+6�\_?�y���dA�����L���c���Ş~`{��]���� O��"56����o�?\ލ �)�[�F�16���s�-*�z�e����B�,
 U�T0f������)`��e�G�.7�j�C�bL���ҧ��&q\�ɡ5�М���+�H�*�]���[�p�⚤����5��q�(8�ܘ'��;MK��K�[A?Dڑ_w)�Y��AA(��I�%\vZ�����A�ದ�
�lh�	I��0��{�C�c�O0�����*{�g6�J<[����3�<V�V1�y�:㬦���\�qC>��G���	���&7��Ȼ����ͻ�O&rewU����L�'ec�+���QWDy�C�6�P  ܬܼ8+��1��y�=5�=�3����|)[amS�>l��6�*������p��H:�233ł�ED��DŐ�8iT�~���U��)*�%��"�4@qA��R�C�l���0����>Ҋ4��z})���V!���zmI�'��ѣ25>.W.]fJ̑71���ᆞYT7}dY>����K/�Lu�:�A�i��࠭�uV�[5��Pu�����	����3��v���~>����O����Sg��V���C9�ѱi��\��Lѳ��埙�t�	��m���m��4�4��F�Z��!���� 8��Bd���r�[�FQ��a5(��4�t�+K��H��*T�ȇu�����s&8<^`~8888A��ݓ���sA�+z�Ñ�B-+u�D@-6-e�Q��&��(@���$9��=v���빍y�o����7
qƝI@l��}ג���V�Ė�lݰ���8���P5�<����Y�~���ٰ��S r�~N9�)�٩i�.�����3�_�찠���{'X/�PJ �{K33>8<T��:���9^�*��ؐ(�l���(�c����ު�}��d2mH�?��U?��0Q�^�gt����e�7*��ڐ����Hƣ�<���dzb�}�wnޑK��� ��{��
*���B��ߣ���#��C�=�4�4#b@����-5.*+�a�AXƵ
��>��� 1gj(9��Ϣ�u_�zȖ�c�m��e3d2���2B�o�=�H�c���xSOa�3�ei�\0�H�4��;�C/��6�
U�`d��b�2�L�ei�.[8 �4dj #r��;�r���r�ز�9V�^g_9?F%�Y#� � ��,@d{�zcj�Zs3r|qV���l�b�j�Tr�S (�����{��)�U����*���������bv�u&h�{�뢱`GN,�ʉ��6��H`������$r.n.ͱX�.L���=5�=�ޱ�fa��Swވ����Y��`#�F\9~�F�Q�,���LOس���rL�-uZo��6��`hC����skg[?�_h�بg1ը��sgd~qA�76%廙M�@�l���>����_�/�L޻rK�Ő������EiL*��u�}D������G�= �� #�I  ��IDAT���%�"��B�FQ߇}D���țo�%k�9��(d�F����k���=�:�Wa\[�+Y��t�8&���ڢ'?�Q�}z��%�i[A	�mVL�{��Ls�·��؋�š>3����LW�����敦�#��w�nh��CF��U
Wř��JGj�>�`nfN~~�5y��u��h=�a کL�B�,�r@9NzR���/����D����_����^�4
���B~LDX����F�ߪw8)x�86y�~>�g�3 
6fM������%�XƈX?�toM&��_�d�e�}�������o�Qs�G��C�gt����6��~�{�_Ӹ�f��Ӫ���e��.�唨���)j��˱���ı����s
l�"�HM�
P}�����g���v���2;=���q��Yw�^�:Ad,���[��ͳ��(Cܰ$f] �F��%�f���L�ƚ�T��e�(��t ��P�&؝ǖ�j0<r|vZ��	o BE���C}�ǪiJ�ר#��'��FfvCwe��=Bg5_�v�^����(b�G�	�lh�./-ɑ#G( .�����iζu/ܾq����ӣ���*�����88�-�!��TmR��q9�JKs�{f��[C��ӝ�P�037-��:*o���+;`�����k�b�,�1u��r��t�WgY��U���Ϧ��Έ3�~�7gp��u=���ey�S��՛����m�*�rR�ܧy��[��f9ǖda�!�����J�5�(͘N=�5��M�u��?���&�^�,ۛ[h�!���GG9L�bp(;P����k�n�䡓GȄ����{���%�5�$�,��295BK��dZ����^�}u����}�Ɖ�P��.�3�+�_��239�tN�}�{`��}�>��@�%�X7��E��-��9z�(�T���!橱HH�>s�q.��0ؖ|���䡇���}iL@�y��\W=��+��Ν{��w9�**�B�m��Z�|Q�ƍ�w
w�#����_����Đx�E��x��]�.+|'�M��T�&V�!-e����Q(\���y!�h��w={Fn\�)]n��"?���+y��eSK�6�O�@�!�>��s;.�) ���bS��z��y�p�BQ�~��#��{�ޓ��o�Q@�Ɲ�����g\�8�3_�T�1���}�K5�1u�ȣ;���UBr��z����xuL���h#"�{ro}S�{�#ˣ~�Јp�0�̒	F�>��VS�ᬗ��4����%��4j�=/�%��ll��zS�?a��48 �N|��<d����F^�F��/X�D0��Y�:!����֥�i�����3�,��!m�3���O����EDWo�(��f���k��f4��3}�:�!(��9��u����j�c����7o�K/��]v֡������<�c�@�z'��&���kڕz��yE^P�����=�hS3�]��Q�Ew%{�A�
���u���M�f���PF==F���]uL��<����5�i��l�_���/a����0ͷT߭Y�"�<�a�ך2ۚ��Cӆ���9�Z�����R#N�d$�0�p�MYt���DLc�$��褣����=���}���ʹ����vL��N;&�oݥz<n�B~c�G١�3�%, t�\޸lM,��b y`ͅ*i(*�����&���Y�Ţ.Y�B@���VcLS�9N�������k���j�ސ&)5rg������Ѓ`���<��ic���t����!l�\��E\0���tO5�kB�y������a��*�/��'�x�B�H���F9��.������QF�i�����=�����[thx�1B�Yb͖On��+KOfZ��C��QO�6r����F��A�b
����(�~W���s`ٚ��5�����ƴ0/Is�S�}��m��J����e�p�&ge���uȂ�戵q]߈\�aQ���99�YD�],MsϜ;'ׯ]�{�cF��w��e�<�0�x�����Q�F�w��������P�Vtqit��/:�&&�����4�`]�A�D��U����y�3�di!���R(Gլ��C���u�.��0-�m0�5g��u�lFj���a���)bJ��˺m��qR��mM���/���t�X�:��M��9]�xrDڊ[7�ӆ *n4�-X�7�/���<u��6�OyK��M-	�0��௔:,
>?�=�P����tmA-�z �N���Ԑ��̀�p����K �� ���}%���b�����.< ��'�ڕ��Ʉ�����=9y������	�u1O:.�i� p��@��+��2�(��O#0 �A�Aɸ����
:W���jCD��:�;���FC�m��295C	 ��.aD���I�C
�4u�޺w�&�r��I��, �dw"FA�FSBd�Q# ��gN��c� ���ʣ�M��H�o���qF�x��֚7/D$��ax�൱�NgI�WbE	�p�0�0H5F�����T�E�	��x� ���Ў����c44|PD���%��5j��=�@�g��{@/P{&?4cԎ{�V��>F�oN��{�i �FĹw�@F�rB35�r'�'Yb����F�*��&������UF>�I�*w�v��F�B���RυED0`L�61 �|`ȅ��c���H9On��D`z�{�Yx!��u����'��"+�az� N#�0`U#硏�OÒbz�Q�w@���=���b���!��*���������[��+j��{����.S���7��{`�3�����k~�O���)�K�O �<5��s�mT��|D����U=�6	���=��W��O���Ď�E�7	���g`{Ph���+��HBĖ�6e:C�$�Ʀ dq�
���Xb�����F֚F4�yMo5�hAq �,�%:,L�02n�����K�v�'�υ�<l]�m��q�ZI1���O��,%�B!!p��σ�T�'E�U�e��"&<ԇ��N��)�!��Jq��Y� ���
l��п/L�0C��6a�5�s����C�ˆr��)9u����ϫ��+{��qj]�S�j}��f|��/�&.�A�`f��nVc����b���T�h4���
��̬*�.�J���;�i���n�	!M?hw̱��KR>&�F.�n���]9D1���������ݓ��;�ա�ӌg`�(
�4SZDW���م��@5Tt ĒM�(�K�*�N�M�
p����ל��ZᲯQ|���6{�z�y�y5ײ:�h,P�Rj�}Kű��j��HZ1o��iǢ���O���tk�h�������Ѵ{ ��7��Uc��'��]�������˂>IS�Z����KN�vdY�J���	�H���z��&��U������cǿS2"�0Q�ŀ!4b�k�:Xp��Q?�)\�F�Ŀl�g�E�Cvb��@wF��]�!�0�z�"�^��%}㔮�]]�-Ȗ���Z�l�&�(~��}@P�����N���F6xW�����Ұ}���р=Ù߸(�K!ҫI1�3qSl�FlST�#
@D�.b`V�iϮ,a��m�qa�����[.�ڏ�m��*���Z<n�\�� sUS�P�d�0��~ї�����V��I����,-,r#!����Ѩ��á�wc�kV8;;G<:�x�O&�`��殆�g[�[u��v�mع��?���u^���<�D.&�$��Z����,�*�=`o���]?�}Ӹ������SI�k�E>��~�Zz�M�����w߽d��ܪ�0����%�<�zdi^&Z����!��S�0���ۦG��Y؀�Rgw��=�b��ҍs����ݦ���e�ÇL�O�>Ǝ�4�B��=�Uy�4 ���ȼ)�2��3(�$���]��i�I�ac����52��zЀ�Հ,�ΘQ	���T�\ �(����g��\B���M�k��I�f�9���w5�3M=��X���
î����[po}f�zn�����e��E�g�{`@F�ZL�׈�Sdc���&T ��|�[�z�З���-���7"@5E�CQ���u㙁U��bg<g���|0������܉���hxn�e¦����	%°�yF=�JL3ӸNcu�wej�!��9�\��&Pb�o�>���A�I�n��7��!-��T#Y��XD� ����H��h*ךWk^�aoS_��\��*-:4�R�����\�ߋMueS]�ء�#'��Ŧ�Ɯ~���'#RsО�`?9@F,��󀛋E����U���&�@�<T��a󌫱�ӨF��D�x�8sK��bp�GA�=�{{���Ý��b��jb�|�ZZ�c�v�	��0��"�
:��m®�Tȋ[Q�tA!L<��qb"p|Ĩ�~��m��@��23'�~�#r��i}��4��"0�o���)V>15+����r�=��F��B ;)�N����="�����j���d'�MP��^&؃]JJ[fs�!`�0� /�����?�sޡ�8�m�r\	��cq~F>��O����c
p�Q�pM0D����b�2���G�% ���������Ʒ��/H\oz���y�Ѱw���9yꩧ��<#�������76�b蚬xa���!kkz�����LF��l�P��%e���⬜>sB��Ii`�4#T�L�h�
s�Rd�N�Wp���{ǵ3a�8�3�ƽ�o��O>N�� �G�5�3�=��H��
j$V�΁���&�3_{�u��_v�n��2�df	�}�3O��ţG��qR�:��h��w�H�+N
h�3�QP��_������lc�u�k���:�2(���'��m�~�Nܤs#�Rh�ٴ�^zYv�>�n��f!�t�ph2�)���VG�K���+�7rt�֛�Q7����>��;*
1�W]�QLᘻ;�p�8o�>�:�%�V�ȇ����ո͍{F��#O���{w��{�L%HO�{��>{pݰ�{�#�A..1���Az/�Ȯή��-&,�AJ9s�w�E��BI��R�xk��\��������r�|�v��; ��hh4��hnL�ʄF�c]rﰈ{�:�T���<w�� $��Fl�pAgC�I7RWF�[�D:e�kE�bX����g�N�ܡ4F	?}���ӟ�<K�����r!���4<��)�����$Æ�Z�X���[k776�w��҇z|F#��'��������A,vȴ��%�g��(V���ܾy[N;��7&��_�yg^�,H㑵l���N�u.6Sy�ѳ���
�,�Ùe0���s��� �BU޾u[޻tE�������c�6�0l&`�1x����krd,�c�3)@b�>�&��6��%���B7�i(`m_�yGb���!���p��<=)��ȞX��3�>"c���:��e�&oȉo��~]c��ؤ�D�>K��x'����J�a��ԔL��}��Y8yZFQ"a���qo��P2"��ӎv����zF�wF ��:5)<�"�X�I�3��\��������pW�ʻ�xh��gl�0��=͂߶���-F��!͑D���@�����ў<��'d��	�c6xե��o����m�����o]��WnrM˧��ה �YYt��^X(ha�@��_�����Ze�n��0�'2̌�=Mr����7�O��7�8�cJ�]�{Kv�aYʈ��[v9�d���" �!{_��gư}Z��S����l��w��� t��t�6V[��8lhM�bt·MH)�����ִn��uss/"=�4,m��{�/V3v�=�����o��ʙD\c���ښ��2F�A�'�����#lR�b0f�	t$nL�p�6��D�9�>� ��禩����ӌ�б�h��5�P�YH��4U�{g�ꬦŐ�˝��,b��J���8~C��H��t&'�NP�b(&1塍���c��a�n|����ʽ�W&(Z��5a�Ȋi���Q`���f4�H������(�2�lm��;S���������Z��������+�uy1����?vd�n>f�(a� � ��=�r�f N}E#Edk�;�@�L�Z�^��"%�>�A��@�ڨ5׿�/+��u����(ݦp=�0���i0}�A:*v=��uP%�dftT}Vӻ��"
M�r

%���
�1����>u�yر�Z�r]�w@z��
1����6��Nh�u��*�<N��?��>���Ƚ5���m"�&v�M-�9A�%EG�S���߱�ג���ˊs��[�g0����7ؽ�=)�l�'��5q�R��]Q/��O}J�g��k�\�������Q�u+��5Wԏym�X����牔�OUh,(�T����'�0�V�A��*愦�����D�y��Iz�7/�eE���*�/*U�1�C��bҔ]ě;�\p�N�`w5u���jr����´�fEԧ���d�5%��]�1]����f$�4��#MF���:���eh;<`�"�cU*j�J�X495MQ��uF�alH8�BxƝ��!����ѕ:�����o�3~Z�?���F7�3s�l�q���oȥ�WdZ����IC�cջ��� !*Bt�������UvjnFϷ�Q�OH�ea���Z6����`��k���4M���7���� Tc#�S1��Aa*���P�<�!����Ա2W�Q�mbr� ����"k[���youU64R	'���l-o������8�X/�DI���4����F#tbM�5X1`
��s��Ű��_탎ܻ�&Oԟ�Ze�M���]�FcRY$��E���:ʚFh0o����#)ܲ�w�
W���!��i���ٹY];e��\Cͨ}hj�0Z��M���6{?(�O�{@ѣ��B��7�ns9�8)���tF��(�yA,Q��l��kl'@,B�%��L�Lsey�N,��A�A�#o��kvcs˜2+@�<��`�TT���ؗ���FV��șs�{_��zac�v�ίd��e!}̒=<��v��dd��>բy`�>��:���Om�6��H�:K(FDl5�<�V�����Z���H�OK�&�\��
ć^���U_�!�ĭ7���=M�m"&.�������2���;ۨk�<��&��1�c�ֈ��Ҕ�9���n�."wЊRfl7��ؓ� Ռ�����+Kl�#���5=5����zB�n�#q��0��7��M�|�n�6�^�*�Μ���dv~�������hF���W^a�4���#�eB;3�(hh���9��r��-�����/p�A��j��S7��qW�;.���M��K/�ѥ��_C��3f?(�7>~��,,�xL��n��A�$�0E�U�N��:���MY^9B��͛���S`l�N����r�@�ͷ5�;z�9v���j�lC��S@R(�yք&���I&D�h���{l��=L=�R�m}��r9��j��1b��a����Ufl�q�Ե3�yKΞ{P��o����
�}$M�W��2ʙX�,9"�+�Fms4Xm����f}��\��5�N�z��}G������֦MN��B���0�L߳���,=��s�N��(fR���ޑ&�y�x��Ӡ���ҥ���^t625>f�X3��D����&���$�:`ò�,���bQ��ך��^�[�o�=��gߟU^@Q��e\N�ȳ(����襞l�b��F?��[Q%w��g�0�4-8�y�X� ���0�����8>�"��`�y�PX���k
iv�&��ٝ�����!zV�ů��j�e|Q�P9�:ⴈ~ǋ��M���`�ڹ6��>ǻ,�Q�a�� ?�9�rdR��B,3�9GfDqJ}�T��p�b���K�@l(���@�8�h�T�F1|�^vDs։�DBl��7u	:	z�衟�M353-�48rdY�n��A��$M���{�	V��Ð�H�7>+t̕m�v_�~�YZY�������Hx]F�$qn�G�R��?-5i���
\�����E�����5��22Ko9����-ȇ���� ��ds��؝�5m0k���7`���j���8a�p$��F�OQ�8���C�2M��"�5��j��3�)~�3�'ģ��`�V/D��4�?�����ɚ��QQ��ŉ�5��w恇��y��$7��Z\	�c�d��iu�G?�Fvz��L�<��=�$q^�
��-6������У祦N*s�e��|�dA���Č+���s��Y��_�'	�?�*�'����^X\������sQN��:������#*�w�9��?���/+R@#lx���<BT�k4;��,#؉�9���?%";�g���W���sR��{�.��{1'r����gW��̻��]k�H]w��B^ᕢJ�GȽ�F'��p�m���6��j눤����Cz�1>�ɲL��4*��8��i(�K9@0@a:#N����
!dYɐ(�>�=O�լ��H})�$b��ޟ��	��"�|=e�˂F�+SMiECN��ؔ��C�����̠A[�\���c� 0�Tk�@�!y�� ����Ss.�a���0?/���,f��6�����3�oF�z��:�z����gӔ���@��7�W�P7�@��p�+���5V<�1z���N+�3v[H"�N�	�Ig��I�⦌͌�SO?-�K�r��>���2 ���K1��T�j�;���(b)V�ѳ��6I��Zc�X��2۱;���k���c�>+��){Ќ%9~T�PjA���C�5�x�32������6TҢ�xLHL�� (:��h.k�H#��Sp)��0�����29=�9V��f��5j��5�2�+�=#��4
���}A�IꙐ-��_أ����cP�|�a�^X�~4cCVX���CƃbR��a�P��-i�0�����Z�
oX/2֏}�9�_�{��]�.^C3!m,rZ��I�8�9�m���q�JGn�챛�����N�/��Oc/h����"&e�UR'M�5 -%�Ҁ&��~</qQe���9̼A����ml��c	aLB/�*&��n��HÔZ�9�{�S{��I��f�2��4^;��� BL�f!����ɖ~MQ�`08MP�
^1T�����D"-�>�2�E�����?�����
5prk��5N#K����$�=��SO���E?@	hO��`��@�5"���Q�(�Ǣ£�&���&� HE�����2m[G�?��ٮ�:�ȣ�J/�ߟ�������gϙ 
��M�+�ML|�1&K�G��ŷN�ƹh�Т*VIe!�;y��Μ9�.`�`4��!����Э��Cm ,&���l��z@�>��G�Enװ��Qa�e�6�:{��7(6��>�q9u��;y�"O�>� �����t���(�g2BQ\�4�iq%j ��c���v�zˆ�E�G=>8U��|��T��V��u���{��f]���CA���&�~���B=�w'f�O��P)�@"/��H��dܠ(!Df��P�]�x�w%�������c(��(!� �e���Gl�۷uc�R�p ���:-���t��hlr��3�
�Yݬ-[U\-����Q.2�Ff�D)'���M�l�Sԣa�L�%�5�@��tqn�]���؝IDF����hݳ:\��+�Lh�/�,�݆�vml7pA�	W����t{o��y(X.[��6x���*���D
TnD{F!�2c6��݊��vx��5�,~,,)�4�LCgof��f䅌�bY0�����b���cHi�x��M�B����D
,�0��Xd�cb�H�'4�j!���R���a]�����.w�z2匀�F¶��G0PF��(q�����4Vg8CL�rXk��g�`��xD�3�����7�K���}��-
}�;&X`Da�]@�\o�w��0�jS�2e(L�#e��P#q���s{�Oo�#Պ/!Vm���������Zz��}�g�r�	�D[ި"Aʎ��d-����k��ʥk��tC��0�S������q��2��m�`�H�,�Y�7.\�'&��A�2��غ���=��}�w��ߡhK(�F�[%��1:d���Ǯ���)ؔ���c6Wk�]�M�� M<�V�-`�cjxO�>��i]vz]b�W.�P�CD����/R�r��o߹K�D�Ԍ�L�@��1H_jdW�C;AȨ<�?�N��#=�����k���$D|@��!�D��✆�֭U�9�8��Xw��6������C�	�s����?��lln��Ԅ��KJGVC�B�0\z��Alꠣ���9���r獪�,��:��h/�s������7��,;���޷�˽����^��Hds)Q�42F�-[��?�/Ðaa~�o?����m����20�P�,Q�EQ�&q�^Y]�]ݵ�/�v�����8���/��5���Y��򽻜'N,_|tei�]���o��l��l',�!n���s_�����;�>~�BJ<,eɢ�)�h�g
S���ӽɴEI��N�ef.���?#�{�srg�.#�A�oŻ��E���7 ��d1�<�Z�=$_h�����7U1s#Ѹ������Di-*�}����QIa8�n\Ӌ�ܐe(��=��
u �{۲��}Y]®8�aa=�@�Bf&Ԉ��dY$��8����O��u�$����
p���F>˖����4~뛃2�׮��n6&P���;�������$�h��-U�Qi-���EeK�Q����x���IL��Z���^�?����;��21ɚq�,�m֝�
�\�ɘl�]H��@N`x0fB�u�z�=�=W��<X�a����(_������|��y��*�:��Y��F��3�����(�+v��	㺠kinX3��y�����	V���*���iݚKu��BWi�����݅��s�����,�����7#��ѻ����
��o~췤��G�߱Z�!�6C<nH�%�Μ�0��������zO�t��ԫr%&*u��<X�?��w~����s	�{��!���aƇK7�0���]�D�w܍���u�mΡ�omn�����P����s�Aơ'�N�[h�r�*EG	��4�	��a�gY9��%wb� <x��ľ��u�����Y�\�$��e�<��޶zv�E��+��H�cz0�9���rM�߸Ao�f�� �P������n��>�;2�J��I��| ���t���.&]�׾�1aV�L�ʗ�l�������|�_��7G�_y���r@ڹ��i�B�I���}�1��U�r16�"v�`x���;�TKb�tetr�:�����Ԙ�/��ӗ��e�{��

��jW�}�\�ԕ��� ����F�d�B��9zη�鶔���Aܔ�	�I�PQ3f�2�#'T�p}�\f�G*�ݭnbyP0,��C	20,т��� �b��m[�vgjQ��"#�:���k�ep�L�����@XX,�b�4����{Ř��F�i���b��LIH �5�4�T1�Q�5qzpx Up�Qb�sX",�0X�ŋ6?���̲�V�GW�hվB�*�X�p�d�֎K�b�X�9W�yz�'��2�yj��yP�QQY�nK���;2"�s*��4R!��Z{@e15�,�a-(ģ�н�s���Yϫ��6JD��pר�Z���ץ�>��ؐ]�js��Ƒ��1�U�R����xQ��J6&����˲�n�Ge��ᅚKB�j�������Ђ�"������W.��m�5=ds�JK
�0���D9k�3YZ�3�ͪ�Pa�O�#�'��$\0��bi�d`����>������vH0�]���Q��1��������z�����D}`L	s��i�%�+A�ݾW�ᄮ��x���O�me�1q�H��J�w�o�f�,-����i��7��ʑ��E���_��rO�viQ������$K�{��M���{&1�N��1�7�-�u!!�V0a85:�,(����hqG��L)���a�@@�9Z�L�����1^�f8����qAX�Y��g'�Lqʕ�W5S��=�I�nP�(4 t�/	���O�Kj0·��m�ZYT%���Wς�W�W���Ȭf�J��uy�u�(���ݲ��A�nX_�!cΥ0���1���WN�J�J/c�Q��j\Oǹe� ���y`"S��L���Rʑ!�%6��+��^{���&UYd6�̃T���T�Xh
m��Ks�y�9vck����,��1_-��3c#�9�N��{=�3�JSͰ��p������0��	�`��K	�ۜ$�ӣ������:�N�� D֚�PX��Ʋ�i�/��D��%�6ވ�\u1j���2:���.�n%�� �J5GE�0#�,yHɣP�2��4ƕ�̑��{G\˵� ��=L:���|m�n. `�9�q;-�j��u���&�@�-!���әU�T�j�ͩ-�0U�#�K2��΄��ܓ��Ϝb�C��*�U����P�U�mN��~T���`�P�u�і���JY ��P-pb sZ��&��W�%��ș|0ё+�+�l����e�鶀��"��N��*�i�獒R��5�<�%���4�2��GQk.�ϼ(�,��[�RE�X���s��A-mE�=���%�bĦ6��L�U�����-��X��D	��'k�D)���<7��녭+�1Ĺ��"$�֦��m*5 ��(�h#\���p���E��r����o��wH�_'�`[�k�'��|k?0V���x>MXNb��K$W6���J1^%W��f1�n�cM�f�� `i���s�o�/�k\�(�#˞D1ST�
�S]��25�{�jh�t�\ Aق��x���+���o-�?���d��"�6��/��Wr{;�,y������C�}D~�w˫7n�_~S[�`�6�
�yyE�]�*:��vW�"�p�m�a�!���瞓��m��׿��B��5Z��<��
��G������_��_�}��C��Abd*���2��hfU9
�޵4�u�����ˇ���g^���D��Z�BGe�G+@X�����n�,��.tAJ���A!cb�� 錾j�ah��.v��9�m��[-.�d���
��I����[0�Z�R�4X��E����pLd�J��}e%�X[I%c|����6Z5n��%ҩ�5-�wT���i[c@|f��&�-S���I�.��v?�bw��/t!����E������ʺ�2In������s�ׅ�R��u#g��H�m�Y��qJ�:\�"
+���������4֭��.R+�,#�WM�	'~A�s�f��];��^�a&Y�I���u鯳e�S4��S�ض���*e2���D�%ɍJ�(sb�[�7V��*�,S/�LX}/�aa8�H�<�nD�Ly!��/�X��g�U�n2xV@)��Ceۈy$ā�yRV� �p$���$����ߔ��E�w�) s���y�#o���������`��������{ī���1\�fA�e���N�ÂJ��?���0���,-C�b�	J�?��.\� �x�;H�r�}��kjk���K��b)��db�)�r�4�yyQ������'������`�GkĐ	�B��IX�S�c���X��j�&�c�&�d���w�").��c��eB����C0�Z���&�������e8q��#M!
�pr̒�b)�~׉%�V�s���4[L��UqU�ݤ�:�	8�~Z���0K�J�v���O��Iba�R�����{�'�t�y{�h �g�(��7*$/KW(~����� GD���'V��j$���1�أH�Ba]2&(�5+Ϋ-}=E��.�}꾧��~�=p��j�1IV*z�����C+nᦡ��3 �ia���t��|$S�w���8A��hY#7�Z�i��s�V��	�*c�au�Q'��͛M7�T�*k�ÐX�*+a�\c�w[V��c����$CX@�Ϝ����^/����=�&L�G���ޚ,���ſ���3מ��K_�{�m9���yG�]�l,���]�At4��z
���o|��YX$��3�+�pkֻ]z���������?�q����R�&�u����7&�r�Bd���@[�r-/䉍Ey�徬/N�����,ϔ����T�y-�w�94�c��`����:�� �N�rZF�>�Uf���/�ͤץв��[Z��T��%� �
2�Q�9�
7���ѐHcWÎ��iK��]>���4c�S�6{��В(�x�bsM ��rjC�VcRCL�~��ͣ���2�G�P�T�ҺkxQ3װ���W/Z{莆b��Þ՟�l��fS��Mx6Z߫�ekk���Ҍ
�s���CF�R�k�������ʸf�7𫢲ml"S/rv̪x�y�I�ޔ�C	y�U�7���f>DH��\�=C��}�N�:��a=>�[��+�V}�PP�J�]�r��
q����ƅ�\�oa;��*�JCP3��Kt��d�3c�D�voph�ĒUr�,�����zV~�~V��{LTd,�mqn,�j������;����[��?�grX��G�;�t8%�zcAj9��F�M� ��na��}���5-��Q2,�T�di5��8	���4UdXo�=��}v�T�§��˙�\(���>�yk���ڔ3!}S:t-�����U���n4�����aƢ�S��B.���3^&%��I1iQN��v�E4�Cy#H×�d�]�������+��6�T�Z������HߖY�͕�Xkׯ�-�����9﹘�8c�B��v;f�]����Yh�<��lT�ub��=�a�!3��hiU�����5gC���[��Sll��̮`T������^�v�
/��T96���mEl�T��G7�P��V�S��(D��3�k;U/Þц;�yv�3M�/|~+37�;[̄9j���xb �#�G2�T�湷���窎��z���T�t���M�˂��b;���W��l��0>`�C������3���'H�t䑍K2���ڢZR�ԅ6�C[���e��c��)�L���@��Ĉ�*T2���:� �|�&WZ:�Ӊ��@u'j�3t�\\��h����AAg�=��
qdAa x(�����N�dR�,�e�y�5�J����rxۓ����3L�u;
�F����zŖ�TF?�%?7.�2ם_�%��I����C���J���ʭ���Ú�L����3����y�t@�<��3�\j��' �QE�$á��),�)�h�*���%���lZz1kԽ�F�ٖR�HHlլ���"L\ө+���kr�J���h��k=��n��w��m��&���~l����I�Lb����o ����0O�����+�ZI4�2�E�:NH8�����ys�Y?�*�ט��&�O�|^�.���|�Jk��&�f�Um�f�Z^R˽~�����p���H�h�OÑ�["�Z���0��<K��>c}m������O���/Q	رJB|��; y�{Dug��_M�Z������wX[(E�ʫC�$G�J �Bhi֜�f�KD�!T"�~��@���kqqaI�Ptp({���w��	*S>��&�Jpz"�!v�N��2��7M4�:P���֬a��m]������i,�aQWo��������\
vu!c;��=�r&�
#���:B�%WJD�d�6#ffe�"Z�bTDi�����j%�~o�N��I�6�\E��R��(f�%���� �5f����3�Ǆ��Of�궙iwH��$�J�޵�k���4,�y�/U��R�g���j����M�|q'��ΙZ0\8em�E�˕�.��⵼r��vK�@p�q���EKʭ̸�%���*��'��?���t�S)���u�Z��1*C�f曏��ˢur(g�4�s��U�RoP��J%^�<Gz�Nt-�������y�y>�sc�"�s�u��B1�o�\+��t՘���Qf�"�OK�W�R�+�J��L&��{1�%=��g�R�gz8Up��f-t�l�$��=����m9�i�<�}X��w�8 �a���	�zj��R�#c%�@�&�W�8���G��Ɲ[r��k��?�eǅI��2����t�ƥ�JS���`K�(
�	���7A���;�b,���kK��7x�h��q�16���4�IK?�C�2cU�U�ni6^�ڵT'�c��.�@y{r��ōe���� 3��	Q�G���z{Ke&�~�T̩�µ���b<,��i�����OZ\�߼����sb����(�-j��6O��bi����*y��d�>��RE2s톅x���K-W*�,��Ô�ð�Y�㯔�(X�m�Xժ?��G��|�yן�.��B]q5���R�sg�����ֻ�����zU8򼾞��4� �Ϫ��^�}$�2B�`���)�w�/���g���ٟ�� (]w�2�9V$�΍h��y��P$6�W��ū�ȕk��֖�t���,�vP+�V���������?�#��؏�2�G���e��;���1�@Zg2W�P �K�M<b7��N���L��\ΟY&)���ڞ[��(�)wΖ�e�]��~�6��+��0�Œf��G����a;���������w��w`Mq�2�F�cE�:���Φ�,�!�R+?W�GcaGQ%��q;���9�%��?��<�G�i<ầ����/�.G�jL��kVy/o�H�	��cy�qT��nl�9o*oG0�'�H����r�k��x�)�(ܲ�f��潻qR��-�Q��� ��B/©>E%�~�hҶ7�gP��lN��5b����B���p"jP*	.�fM��y��.�^���_�����G~Z^�sW��������*�1��V���-,˕�ҿ�ݗ��.;�3X6wY�����%���$XN/�s�
�C�R������d:��`M����bG�,�
��9�2U���O��%��5���,mA�%��p��jTO��[�����YV	��I�'��y],0I
?\�c�����(6���J	Fƅn��*���	�hTa��5�⦧]�3�ACA��5��qVQ�~���VɦV�I�8��l֪L�=Hv����`�C:V�UJ��l޳��|��t;.4p�gq�$����5�p�Q9�(sd@2�b�4�:�7�>R��Ǒ��H�Q��X;p��9,z�j{�x��`nO��/V���4�1ږa�7%{�w۠�-���f�UV�^i�/�	$[ʖ,w�kO�J�/�_���u�'�Rltt;�z������.-`u]����,����v�.U��MiֲH�����HM�L'.-�k�_�+�?�օ�sA��Z�`Ӻʘw����}���,�����!	Ƈ�<Z��
��/&����T�Z���*U�1���} M"�:��۲V�:\��a�z����D�ж��OOWZژV��Kl�[D:��s���]k�U4��mn'�kZ�^�iQ7�?ދYOe5��gB,o��<i|�c�qo�WS)��:7��xos]�^�q�<�=�s��h�^��4�q�����a��n2�y� Hְ��B�<T�YU`+i�%j���;_�X����	
�U�D�ApݡKY�g	����H���vQ.TPڵ�]Cَ� AU�M'2[����y�����_h��a�\:��vH`�b�J�Cou������QEw���ϛ�c�xΈ9窰ѝ`!(Õ�%;%oA�{d�s��")�RVa3%���$L%�*:#뙘u��!��V�aP��4E���R�K���)�{�c��@����	�h��S��aۓnG�UY���3cˊ#N�<���1=����8k��6ϚK�4�1�n=��<9ΝM���4�����fV�<��
�^�A��~?�gO��yG����t�fx9:N��t�������O=6E�Ԇ�VĢ���@�{|)�"i��4e�-mnG} �,��hJn�̺)�"[F=T8�v�+�]�I"ΈY�e.��4XHY��A��?043��Tr��;{F>��?ο������!n�����w�~0��2���a�Y7�8��9���GW/�:�ؓ�^.�]iw��3BY�(;;�%�#2���W��%U��Py��,V-uÀU�6Å���|5��Hp�*�9ʄ�䂞eD`P)��De*Zj{ ���v
�L�����tOg��F��XϽ�����f�l�h�xR�y�y�7�H�N38o7cǧ��8.��|���q�ޒ5��9���i�H�ooUɽU�z������M1f�O<2o|2�J>�>f7�*z�X�X��&�g��F�����W���K�r����ۯ���{D��縐E醯NP~�K�pDF���aM6.�;?���%��[��������ӊ|�?�џ�~�I�-/���oˋ��$/~�y�X9���J]�`m=��c�K��Kr���ݏ�^P�/�aP�k���󹷳I�]��˲����l<���#�,��Gw%�E�6��>zCaBK�g�HSt RSd���t�O�~B!6��*����h��#�pK�dXş���Z
���Ĉ�˕�>w��7��(C�CV�TG�/�9�o�I
k�$Vfcd�{�3ǽ>���]Of�3���L�ϴt/W9�(=�}8�2;�~�F�|6�8;t�AVSc��+"+T�K���=��߸/�*��q����ļ��ѣ�qy�$��� �GZ4�`%o�Oj/��CmURH���rm���{�
?����2�o*(�sK������kg���=���������,,���}�Ȉ�|��6����X���d�ޅ|�_��O~=(����{~L~��o��p��Y�	,r�-���I+����d��ַ�)����X�zKt���#ݰ�,�x������/�;,vsy���#�~Pɰ*�SkwwPCeNP-���!&"%^0ዎ"65����z_¦��O��P�6
.8Σ�񈜂d���^hUFT�����,�J�Ӌ�E]���.+rm���@��=�����J��m�b��T&C�6��>� ¹W��d�`�ܬ`NC㒼D���-� <,�j���)���M-���u�:�*<2/qq4_Y��|?�j�%W����ɣ��-+�f�[�5��ϫe��f�F~*�x�e�9 �>RW׹Sa[��7��f��ϫR�{q5�%5�]	RT�t7�.Gp�Q���S��2��WtyI(/Z��*�˽�/ٵ��V��QX�E��<Q]Ű�R/��V���A��M�G�#�i���H��i���!b�	��խ�ըp,u�eQ�g���HKu�znU�1,�ܸ��V�w��/VߙX��b;�i���Ow��~��>ؑ/}����j�Pp���v��+?�?�>��?|�Ѡ`W�@���w����,����>b�n��Zd�^����v�x���=ebo�c�G
h��������GnPO?���z�%Y�ud�2�6j,K�)��B2������fd7���5�<]Y��A	A���),ݮ�^!d�����,X�`2D�1��G[c�wH������}f�2K,"�R�Zy}F&�D�	<^���J�L�-��o(߭T�Qe�������Iy��P���i�����J���l��}�-�lƞ�E��ڽ2k�+�s+.=�/�h�e3dD|V��ޓ����T֕C�K�ĉp�Z�����q�1n'h͠�P��ԕ��'b=�m��f=h;��쳶=�-���5W�Oe���!#'0J�'oQe��4sr�ʴ��7�d��������}^h*�A}�ӿ��q�C3��ENi�U�P�:NX�����vR��*�ɪkJ
1��{��9�����ݻ'߼u�qC�Oɫ�n���-YZ\�
��H�p��=�����GzX[=Yj���z���3?Df�o}���헾/ۇ���������|��o�G>�a9��n�TkT�|�mO��?!7_�5���M����Κ�5�mn��Qɦ�eu��ޕ��`�DMY���.fĘ��c���l�uYY=�T���D!�.�_U���	����j��N^ZW�	J�Z��^{�,��[����|n	z�R�BP
؉������=l0;�N�>����:�=��t�Osޙ{��.W0��;�}F���JfH%�x�sUiJ�������&�\�0����j�Lٸ(���lD3���Y�U��2Zh���lϫ���e!��kwCf�)@+U��Įו�>�d�����Qh�D�V`���=���o,��M��:�
i��q�ied��8�HCg�����%ڹ@�����jw�:���r��ⰌPs����7��R|a*����K������ܾ�����˲��&�g���׃b��g��Y��t�-Yo-�c?F���p,����o��?�A5dC��pݫ�.Hk�M�8�]!�`ŞR�E���/��^�~�5����}OV���_��6�I/�eh1�t�z��M߫��Ņ��]�=�Sa��`��ʺ�Ν����?,��-�^��[ߓi؄�[h���i�3��TGt-����B���d�^�ƁUc>r��Ę\fᎲ��d3���0� �hY�,��`���銘׬\���y�BE�B �&�%Q�{}Fس�1���qN�k�y�ްi��=Z�U�A�xǲ���qoy�����]���KK��w��3�Jn��γ�n��lS�L��B�{+"?9��4�T�%�5�~�ҫ�o�Kԍ1���YX�`�e=�@�/����8�ʹ3g�eK�ܙyT
}���C/Ԛ=����*��DU%�����xeL�نe����0�ڵ�*�7���'�jxpl7'�x�I�ᛡƓ\�d�7l�sA���.�k�ز-�$8Yt�̧Y�I ���ݻ��4�)'�����IyxnqUV�K�{��$����d.-Y�ɣo{L�;)(���@�n��N�]`Yml���l�=��b@0v44e�
�c��ܺs'��-��v7X�o�	�V5U�*Y>sFv�ñ��;lP�
�<;9KI��*P�u�i�ve�E�л�M���YT�x������/?��R�v�3�-P�;�ϵt
t��m�%�H��R����A�W�p.��s���(��b��?�dZ�i39�u x	�[
"
��p_.�^-5�{��mfXSA�7�o�hZ.1A���H� r�~eqIά�� ��ġVWW����i1��t�!��Pz�S(>(+*��<���u|fm����6�%�׽p�|<����	��v�����I�к��4���[9���	���cj}}�y�G�ԟ]�(�	�*L��Bi�˙�|�H�E�����Pń���pƆ*0A��l���餈u歌���֬�,G'{�5��;���LH�Gj$5�ѕ��d�MX�|�K,�O)y��#�/�\�{a#�t�A��j�8���aw��y_�\�,+�y��G�?���]���.���{���~Tίm�h���6`�>`�JАl�?��r/(����۴r��ec#��V��A��ل��);��E��E������|���&h��ܗ����/i�ڰ��*��;�c��3��$q�Hd���>�JX��I�0*�o�Ko�'��`�`��K>����o,�h"�Y�k�ͤb����z�P�%4���j6O��3�Z����%�T�2P���D��J�7T��4�������R�3��kY͜Wr����'���ül�l�U��:�`�Q_�s?WU�z��h��J��V9�兿C�Mv��Sļ{���5BI@���l�T�l��Ս�I3`����� (�Q�|ѯ�ܹ���}�1���Ӹp�!�z�*(6��A�A��k:k�pM��[]]���M��%����m�a?�΁��`W����;��r(�%��ϰ�>������K�,B'G�R҂�T�|�z���#�<��������{�4���lp�g����p��PA�����!�s|$�*u<�����s}Ấ��f� �aϵ�)a,Cm:[+ٖ�"N��L4���>+�?��|��~ޑ'yT����R�)��8
J�ۯ�����Vʌ�e�A8(��ٯ|����{��{�%�� �@﫰c����vtħ�%�
��N�!7�wi%�
X�/˅�W��[7�`o�q��7d)(���_�q0���>0p���v����C%E�\+-Q����+a���a5X��
��+;����H����~�n�N�*N(ЉB�@c8��T��0#	tƤȴ�����*��\��	��m�_*xB�*���~{s�e��M�k��P�^HPS�u�B,.��<k!u�Ra��O[R�
��3�Ѥő�Hf���g��%�<q��;gjkYl�X�9^��_���$�hQo��
�k�L..�	��``��y	9��S���l�T!���g�X*�{p�hx�6���n���!7��T8�a9�k��daa��&�*&���s*���gΝ��`�noo2FL勿�F�r�����R�J)/g�&2�_��^Zҵ���o�v_�Xp���J����iI�d�=ǅ��;�<�{��^&��M�Ϥ6��lY�?C�ʁ��`��5�]���_+��b$��ܟʸ+���r]@�Ͱv�6)�P����n]��n�V���8��-������M�G������B�Z�L};L޲,�WH���`tpH� �/ �;�y���bF�y$[[j@�^~�t�@���i��d��헲�;���y ��
�#[;a�'��n=f�ٹ!��=�}��ҷ>��|t(��V��'���tZ���T�"�)d�Q	�0.+V�e�3��#'�Q���w73���g_
���(����g���i��q�\t��:ޙ�0��	�9��I�<�������דD��s�0�Ow��� +�����wXQ���m�t7aIQ�Ֆ��i)�"���]��z�zx���W�}�����i�qp8
��x�	�ġ-g�DE����"1��Z�t�SkHK�rV9n4-�C��z���\� ����`e�σ1'��Zj�0���"n�k����V��"	����!�-g����!/�e�S����f��0�pĂǃ����BG�(	�w�cqԐ��d�L-EH�Š�!�r�l�=�.�E2$��-<���0y��P��3$��=���'�.^[`�f?��+��+Z�y�#ctje.&��c�`(�V�֩� �p�X!v���-�s�MZ���=� ��c�p�*L$������*吂�D�p��|�wL�g�=~�䠴��`�I�e�1w|�,l֕�éܾ��N���V��أ2*�as����C'�)]�)���CHc0BuU�l*dZba�8[BUU�c�Kziz�⮕* ��dzI� ��x��Gؖ�����lD��.�0X{
0�x���;N@�=��y�b�ܒYȟ]�����ŏ+w���5�,��=U�h�[�D!Bx?��K��������@=e/��/kq��^p}�j�p�#�ͬ���w�2��g�!�ω+�����a����

+�Q4D���-�t��@GFŤV��X\bY5���`� l��®��R�*I�jwx�"����6"hF#��\��.���-`�Ļ�����A�˖�!YW[�=	| u^ Kd1A)46��1�0�7cDϩcLo�!>Á��	QdvO���&������~`	�q�d1qAe��o�e,�q>��lHk���#��׾,?�ӏ<!e�����@���?%ۣ);��_�([�Z]�e�1?�a��Vd��(5c���]���[�����D9L�SCon�UE�[2�J��߭.O,��z�il��,R�Ą亐*�}�����ڭ;���q����l�X�N'�m�Ga����qp�$��l>�T�����o��QZf�JVy�D "�9sgMh�T�t%[+�Y��0�2h�������z*nēz�h�?�b��!N�T"�J�����q����f�.)�G"o��n�Y�AW�(z���w����n�ڀu��Q�pEO��^X�ck�o�2��1��J�У������?0���r>��<���lW�,s��C�f�����pĞTd��B����TVn:t�N�|�3kW�����G�L�i=O��@ܙ�o�&�$`�"$E��W�ʍXӘ�`4l���zP�������*�_�#�B�,Z�f�s&k���*������l%�<�e��D��μ[���9���^�_�X��2cQQ�Hշ0<�&�!���#�ٰ���]Y���c�;Kc�AX��ߔ��w~K�aⰠo�ߖrA�,�����My�On��4ࡺ­�NFm�2)��Xǐ*[��fe�b�+��c��n����f�f[�t$<��X�Jj��s��8�����7g�1�7V�4�~b���6��ww�ܪ�bw*]�=�hv�pC!���p�Iɸ��
Qk��l.Z��J�|���I(QEov���vl\�c�y���C�@>t�����6��l���[j�Cz�t���Gw%�1�K�4ߛ���r4�#�I�)��iſ�XYnNh�,�"��H�@V�Q#f�>s�#��P�Ӥ� >��\�b8��Q�wp`�23�h�ZY�أ�F�f�n��sG��ܿ|�]9䦠�n�>־�ͮ=���5���4��
��P�]�F� :aM�Ah��"�m�U�P1i\��4��J*W�6݊B�xW$ƺՐ��A���]�S��s-'����.G�C�����))nZ��8	�6y��Uf�+zT%Jv�f�Е��M������R%�XM	�Zʴ~��&�C?�Ay����[�n˯��?e#E_�i�ۭ�y��m���w�K._�,/��23��hϟ?/7nܰ�E�����W3Í���O?��|��_���1όPR���^���0����T��M�lw,���9�PRT���Kf�+�J�F�ʨ`ǀm��E�[�`Y�U)����r� (�,��[��K�j��ƞ%�� :ă�=����ʲY~���2�uc���\�1k�x����H�+�ܿ�`��
�cȚ�h�"�]�XдN`9�^\��dDˎ���,V��Qj_5O��E�����*����X�VG�1q��/�6���HKigw?X�CC�0@�g�^u���9q����N[{ϳ�f6<�޿�w1l0:��:I7W�[W*~-|���Ӫ������q�r UB-Z)Z	
�V��VZ|W+���<I}�ei��JP��wp���@1�{`�+Q�i���}����Ɨ׹� ��4���M�s8s�\R���a6��B��Ƀ5�A�jT��$%[u��s��w�O�������²$_�ꗂ��"��\�����̢]��m#9�8,�_��_�_��_�;����Q���C ~�4)���s����5ށ�i�#ޯG�x���pooN��v��JƝ�ŘZEw`jn>,�Ѹ�P1��h�����_l��b,�8l�$J��|<�j=�$KH�!�k���� �`��\���q?=żd�<ři6x��G��Cs,�����ռ�t������Xxa8P�m0:����
߿�)��P�z�8h����e����!\nXwi�N�)391�@ˠ�Jp���F��*ٙ1���� _,�I!]�ͬ�I�����B_�a�����Q�إe��L�[:w��R|��x-�k��4|�f=nT��ou-����u����|<��tF��Kʞ|�B���F�x���ɓ-�V���v%�	�c#d,�M���W�F�b�W����c�L��֖G._��<�.�z�!y(|]8sI��%Zc�!��Lޠ`�牦t�b�X9Qy1��t�|���'䩧���^z��ôs�-k<�״�|�����.-�M3�~��1��bM�2��_+k"�Q�I7��}�;�bY���t�U|,,X�� fh�)�¤T�Xĝ�U20����*�J{�FK��ʯlsv������ ����d�k��~�]V�Lc���t��MoZ%��|�9�nM���:��Pj�\��Lk�ݷ���5룗[�<�B��hfx(g���� �T@��VnV���L�\ ��kW�K(K}r��wP�]��,��������?#���ѭw��������[ȇ�`�8��#���������2ќ[A�U^�v�w����)X�����㜗�ƙ'�\>�����I^T3w�/�õk�:q�>��ƹSK��̼'Cdd�B햖䇞}2i	Fr0�հ�.�_���.ʓW��ӏ=!��/�B��DU9e�2�W��bi��AZ�c&E�R*�"a5\��0�N,
R���E�'n������VCj��w,$����R7�cDZ�UP����9�B|}7l�3�eTO�Ω<���+���"���Ś//�9�8bp�U��]�5��3���&�E��xg�؀��}�Z
�CB4DF�%�xVn�<u9a~�$,�*��,��%s�Eќ�y�J��7�>�PFKK}y����q{�dmss_۸O+rv,���l���6�RoB��J�4P�bΞ�ށ+��e��y����.d��Z�|�,������-�KBE�:���k�KShT>c��oP�~2ͅ���O$�GB28э<@x���[�1�.^?��$��eU���8���%$dlh
���F�>_|�T֜�H���&	M�����U�����^��+�5��~lʘބίrJh�p�������D�d�6���X�q�q�v�`�^$�V�j���0*(�Bv嵻��;/}O>��/�0��������Y� s,S8�2��(��}�G�'�'��_�r�=!>%��~�|�va¤x<̭`��
Ïۚ�b�t�@���XBz��6�=*v����ƁB\zm�]q
�)u�++,`��UqAɢ�S kvjU]T��v�
�g��g�ĊM��V
3o��R���A��6J@�PͲ@<�J*W�21*8s���ɬSG3��5CD~��߻wO.^�@Br���^
��]���`$��I�7f�;�5�yGv�$K��tO`&���r%+AZ\Zd9)x|#���۲�!�XT��={6|��90�^Cd��uk_��I;Xc
�k��#�F��-�����j�c��mz�����<�X�b�5WZ홐Eꍸ��]���-{�S1��ȩ��|m�&��'Vq4�雇[��a#u�YqÎ�v'%-��0A�ܱ��J� f��Շ��3�<%o{��Zɢ4v)����G��+r�������k���{�p[vF���#/�z]^_7�ܒ�;�eX��&���o��q�w��w���Y�цm�Q�2�믽.�΂\�p����>�� hZ;��`�\ۉ_y�
� mµ�f(}Ě0w��`Y�a
v&aQ���2 �ms�SY�l�	��d6``.2eZ�
�7����,C��pY�K.I�Y�ʍI1��I��$T�y�(Ɣ��_7�9�3yn��BM�Pl0�)N�L�k��z�R�MH�%�~2�>�x)QṀU��8,�e+P�T��P���b�H����&.��=7�pv�,2Sn^YE�t)��oq3���ev����0���w��ߍ���.��A�Y�4�[g�gTj���Z�Ab���c܀��c��;��2�,�%���\-2,;��������UJ]�h�zuO \�'�b��H�ׇ\o*&'1�"�M�Ţ�"G
=���t�h�*���$Z��)��h���?H�4����u~��W�߉��hx�O{�7 �A��������]��l�Y
�r��JNٵ�U��y��Y����O��|�Ƌro�+��9�J��	o��j�嘨���<ovP(��V_V�EiMs%�	�R�O����?�gV��3�<t������T���kD�B�v$�]*�5h��p�	�[��\�]�t�}tS���a�H�2�_T�,�z��H��X�F��5�W+����v`j3��̀M3s�iy��Ű~i�+�D+�J�ݢ�>�^1�������M�����U��S�	���9:�T��uθ�5ʬ���΋���H���52/�T�"�]�v�j��3����DzE)wʘ�����gu*��.�w$��VZ_4��mt%?7�R̩tŠ�-V9�޴�xzC|8.����&�;�٪�Qn��8E)o����"�sP���
�w��t,v����\���E�(�@b��p.�<��-��U9����RU�iw���i��Y�|��ӡ�]��9O���[lP�G�wKNܹ�M,9za�	�����f@0�LT�ܺ��nc��^]�Z���f�f";M��"�!ZGTD�`-L�  qwx��X���>��s6:�:�m��@�W��7�[�_N_�ޥ+	x5�`�>� 啵dz��u)v���ױP��2�W��&f�d� �.��W��i9�C::�����������HE�+x����쁭]ZÅ��ekg�ma0 �@�qg�;Lϲ���4�ts�"gQ��3�q�|�0z�a����U0|��m��+�0c)e)
ֶj���R2����_��R ��-���J'�%Q���!����Ƹ�a�̳ͨ��DE禵TU�ѿ�c]��(����)��2���,��c盈�S�3K�!(U>�ވx�S��-��	����~�w����*��6�er��ʺ���&�[��pd�{o��Z�u�U@*xoU�_�e9n��Wɦ�6��iKK�)�>��v�z�NL6X|8���G�e�O�kK�"������h���*��(�P+K/}��0C�7��V�z���ܚ5E\X�='UeGCQq�Y���^C;�Օ5��_�B�]����ݔ��+��3������G>$o���W^�oܐ�v]nݹ%;��`�2���q�+7.���m)��'AQ�"
$YZy]���lY���o4��t+(��&ZY����ߎ����9��
���6H��<����KOIe�@΁�`����'�tJSB��@�~��0��\A{ʭ�݅Yq�(ٹ�����=7O�s�ǿ������X��ud����{�fު��DE�b�{��x�4��Hn�-����ӤL�ZVb/+Ov%�˚�'W��ƿ�E��=��Y��[-^����C��w	A"F�(��zC3M��fm�vaۢ���5��1�*��*4�F�!Zx�|�Z�@I�d�i��N�\G�BE�`�c�=�h��P�{C�Ly��ټ#����j(�2dyY��{3�.��]����3��ū��ÏɵKW�wF;�.-?"�]}��to�<������|��+���=)�G����/^p��=Zm������r�M�:�8�]���ɑ
�7\DŨdR�+�[P����4Bn| ��������	3G�B#�C`}c�����T��V7�#�W����W�d0�+�����Rr3n�&�M��{r1c��~&c����Rڧ9�s���#��SYD��轨Ǧ
�J4�[��9V�^	���Js��N=��j+1�3�g�]
�f���Z��_�?f�ݕM� E�����>�	=�C�hn���Q���Xi4K=[��F��CB�yU�Z۪���>���dv&�@��h�Yk���WWV䩷=)�n���C#02ZJ ��h��H�^nJ�\>'~���;�k ���ii9�J�Nn������ͦ�/+�M�Rɵ��
��>Ϲ����a������[/W.�mȳW�k��+�ɕ��i�.������G���O|��?�����eܪ���V.xY��Dh� UP*Y�����!*���*V2�2;�`���P	+:-��\}��p�ҔL!E8n�ﱹx��7�S8�Z��..���B�$!U� ��t7�,��9d&�!�("�'y�.u�R��$���3Ou��j��q����J�qn����;�q�I�o,*K+N[#3
��U��lç Eʭ�_����p�jy�t��BE`�ȁ[���J�e܋�$���qeL�
Y��V��U�0߅ ���q�Xj��r�2��~U�?��G�	�wz�ْw���nY�kc�d0yG���r���4,�t>�9�_�����u�An����&�RB~\	��H�I�P�߇�_���$YK�1�;�(|���X�j����c�]6�"���,ׯ_��^W|�߇��[jɫ���/ߔ'.=,�^{Z�x�Q�v�a�z�rP�$E��k��ޗC�;b��7_��AM*rpp(�%.�l7�$+�q��I-b��Y0��V�C���;,fp ������F����H��uT6��E��Ru���A���a]N�+�exg��ݺ6�O+���yF�B��b��vZ�4b����c^Ib�[�IG����|�'�;�P��s�����������ٹs�Y
�u$xP�iʙ3k��1��Cr����/+�a�^���5�%w����.D�������xO��u��G&�.m�(�۱�@ �o]#�F	��?���k8/>�E�1$ׁ���]Cd `i���r���T8V��W�i-�5������Y�U��#��ϗ��I;�Vb�`a)q��:B������ X6�٘��#�̻�i�f8�6 1Gz
Q�VG����Ē�)/��ޕ�_}�V�Pb �-0�N?�ax�w�^��߼!��O�����>��g�-O<�6R��%�)�FXsv�uak\LB��֕CGx�u������j��,���X���3���SI�(�2�;���4G&�J��cUk�����"�Tz�q-��3�lɞL�7Uca�r����ъ�{��R�y1>��6��p���	0DꝾ���8��[��I��
�y^\�sN�6�1!}���bO[[_a|�
���ȽɘP�%��	�mog����9�tᢼ����?���~h���~�F�d����衄��
�t����2�Ne���x#��+���`��m��:0��������g<g����?;	ϼ�w������.���Z�2�dJc���r�cB�E�6�X��he����&��/Yw��|b�$L0���ݲDW�F�.�:� �F]��_��R�:)��hzL�Vc6�C��DhE,���Oj[��*�;�]�
c��o}K>�?�$��$�Fd(��a8�1� ��v2��^���_�o���r�ӟ���=)?�C�=X��R���T����I���_��I���^9��N���-�p�G0�W@�hXW��T�������5��$V,���+j��ϛ��j�<���m}�� Z<�fD�>*:��J��k?����hbؚkָG��ٌՕ��3;v�,���?�O�3��'>!������{))�2����Jb��f8�qi�y��{os�=����ﵸ���XP:�ڂu71X�R���0\�
tkK�����|�*�M(� #��X����#�P�p~'u����C��q'��T��ՠ�Ϭ��haD�4Z��2��[��O�Mpzl(�}�t$�;���=����+c�C�� z�^X9 D㮞�T�7��2�)�ˋ�>f+�%K+c9w�7!��Uƛʍb3��r)�8%Ή� �.�w�ѸbXgj��t�3��YH���L��%O�t]kDe^iEqyt{��0��r�s�*Y�oY3�eV����������/'T�\Ho�x-���l2��|eA�n!���Ʒ� ��f@[b3}a�A- S��O��q�1]��fև�ws{K�� {U��Z&p� dkK+r|�lY1�C��%.;ᡷ�N�e�q.:$p ʘN��L���UN&�S�ՖH���*ʋItܖ*l�FYl	�.�A;S������L�EI��{=��b��Y�%��Y%S�NOh�v�n��S2����0�^�L��C����׋��/��م�@�Kb�����zH�m�s��S����b؄�R���!W1H��x��
�Q`Q♈���$X< ʣ>�jɝ�������X�y��a�R���r��ue����9E�I�m�� J��LI���d4V���|n��m^���@R�L�z2�9�ٽa��"/,
�%�n�Pzx��`}���\�ª�W\)\	����-@ƠY0bvwv)�Y+#w3�{euQ��w����z�l.s\G��z9eg��B�����9����E��Cb�o��2(�'��������I^�L�QU�ogBkR�`��~Z�V��Ɍp%[�e��
� ���5�%ğ�]����ݭ��ϔN/3Z�����i'͛�U�0p=�:��H��Wa��!�C/!�����C��.B�0Zݺ�J1N^�(����@�rUa!�.����+w7��L:�A-)����)�\aWLMk-�
�������,�E��nj�;���f�­��lކZ���VF��P�6��EYu{��Cf��s=yn��'?��O�'?��Xf����Ą*d'�]�bp�)�f��ߨ�c�~��Rh8)(#��Ye�x�C����b�-��Y ���XA�ńD�%�q;?�����ëT1A��&6vYT���l��;;h�	%�E�;[�Q�ăB�ƕ�Qf-�,**�P�^%\���W����a;�r���Ƅ-���j�n�m�+���b�9v!�dsk'���9	����2�2ܲ�-�z����4���%�aNz���ey��k�P+�ƪ5٧�GR�q�N���ܽY����Ol�9G��%���<9sk63����t�Q��Ls�4���]��b��	X�cV����?�S�C+fѵoM}\�L�`�O+�L"|�u.2�쩾w�l-k�1���J
v�n�a'T`�u�ۖƢB������
�n�	Cf�'��56�
w��˕:�+���JStDH4��1v���T����T� 0-
�L��Ը���b�f��ػ�ޯ�X��1�$;|���P���w�V��BXcSk�o��i�'��u�8:��'#��v�z`�s�-[l|�n���V��I�	�*V}y,�����܃qNX�޺�N�(:C{���kXӀҭ��͵O��b�J�0��kH0DXِi��5C�p	\�Ä/��[��b͂��V<ƴQ ���y��O�(�`����<Kb�h�уrx���W����"�k8
�-��=U�lk���Q��ߥ�¹�R�5�;z�u��z\�������|,��d��~��NR���7��b:j�U������$ǫ*~���Eך8��0P� $._�\�}���	Pl����~��\�3g7��g����f��ww��k�Y|�qF���`�jr����#c�I�C� ��n�& t�l�d#;ny�@X.J�Ůt{K,�TNKb"i�	�;���5���4�$2R�e��C1;���� |q�Il
�9��=���|����0�F�Y�%Ű`A�����mU�ȥe1e�/�P����;��+���@�+X'#v��\��06;�(��9�t�O��a���'�����l~����;ŏ�`H�I�>���A����0 Bk���/W*�N�įI����k���������r^5ƴ�Ѿe��B��a/��C����5��jWj ͳX�a���d�x-���f�Y봬a;Ӛ������)���/�X*Yf	��5��B�ep����n��Fw����'S
/����Nk��S��v	m��p�ֺ!��`îp��9w�ܺuS�|�*䀤����<;A��{ϿH�	4�sAI�G�i|�SxX;p'�hgS@Of&�3�l�n+k�a�[B�\5.����f��+�.[2	��h��
[�1>s��u:r$k:6�\�_���xC���sc����&;�i �M�<����L����Sq2�b�'���\8�LoA��iY�(��8�C�$�NX![[[,�jo/(�ñzv=Ƭ�*�/�yp
��@S/
�U��%�����Cna��'oqLj���`�$C�c������K�3r�*&|5$J�vi���F|cu��7�6)jf*��*#i<�1,=$��g�3�B�	�Z$��7�1����YE#ʁ��o�ǦR>v���?��4l�2�|'��h��e�'���Ә)��_L��P�ϸÚD�:��H�K}B�SKߪ�<�DY��c"���� �;�N�I6/�d]�x��?�7~F.]�,���� 3���-7���T��o�.��]Z�P�]yH���rFI�8Ϣ��v�K�� �]��L��p�v��"%�Qa� ^�;�z��tîbhE�L{��[Q�"�&�����*�sG�v�����ʂ��U6#�f
�u��L�խ�PS�aӒh
m�r8I�S��s���P3�����p�aс:Yv�{�,�V{��v�t�1'���hI����t3̭.��
���&9t����0����ܜ@�}h
�m�`�����I����(-F �X���L�NŻX�]��j�u ���X���y����qR��a��ՠ�,�\X'���}�;T�*�YIc�%V�S�ՆV�
�&y}1���glz�f\�j�'���dSK=#�拿;S]�?@~O���yE@jhX'��b}3\x,��fˏ��������ꐁ��ͯ�!�H�~'�ra�[�X��#A9b����^�}f&�����pv�^xO���vA0�ݘ"�		W@#�ɽ�F���るcV,?0�t<�3�3*&�l�v��0R�$-���j	�<��T��+/�����mkL���~o��Mc~G�+�-u����
�P�oP�))���,��..�>o,�H��H��B�x0�e�;�0&Iv� �W_���Gl���A6�z��*�
>�o�nDx2


<�Zh��"V�7 6Pm���#�]Ӿtpq.`l�,�|���NG���󲼲CS�dއ�Y�n^H���[�i�j�I7q��ސ�&P]�yG��LG(xq]·2&����"zj%;��l:��x��` ��,���M*;鸥��[�Ǧ��o����2���2�O�L��gq5�a>/&��^�tG��������3p7S�^QZ+tI��*���ԓ��La�����J���s��ϑq�_���=wF��u�>cq8P9(�Rp��tH,�h�y;�I�2UY��F�{��:�R���L?�q�N�GK�w	�(���[�ι8G,T:M��889~�&�*{�킓Z6j������ȩpE?=z4��y�i�q�g
os�m��a�k���t�RZ��v<���.������VPri_�iyz2�����51���ޓ���\�|�	)xؔ����e��ش��Т�6HǑ����T����\�^Z��\0:�d1^P�ix����id�%�)���Ƃs�a���4���F�� �B,u�b&C)u�UWό�������|/`c#���>|�i����c|R�����ϞZ�5�ϔ�=C~y����媤F�b9*vǩrAŝ�L�V���I��T?�t�Zh�L�\�Ow����n]d|fE�ұ5�T�;r�������lPΜ� �09��"�Lbm�C{mY\^�'��w��n�;N6pf7I~�_A܋�+xv��KMn8X=���\�����
% H�%�[:%�`I�KQnL�7�A���DVh(�6�!5� ���Ea)��}n�EU=��FX��⏅a[Y�����VVVo2�y ՜M�AI������s�,
5Jb�D<��|�C*7C��J��h3�eOb=[+��X�\c`�|O�,[blW��.7�,Y����7U:Ax�, ]H$�V����UB�XD1��*~w�2K�c�N�%o��	�UQX|_rB���������ږ�7v��\�Cq35����EX7Cz��`�9�-жA��?�;C���lNcd���<�v�y4����;C�[�������jl�)�e^��"�W�}�1�}U���k@�^)��*��Ojum�b�Y0������&1�L�J�����UA�������PȠ(��8�?_�
63��V���X��7�&{����U�>6��Ͻ_n���Lv6�.-��W��/L��{�?��o�?�x��@-�.h�J#�q72$�IP\U֦XC$����C��V�^X��g�!&7�X��k�GBg�����_������Cr�n`c�D����{���AkG�&�xp�LA�x��F,	����Bw؟ӞEטr�B��(G�K�l���RNT�ݎ�m=/�;�;Y�OxwOq`�a]�?����<R��P�hK�9���_H."L������@t��_���9Tf��РUU����Aq��������������6���.�.Y2$lAA��5Wt�W�͋{�ak���FЦ��܈�&� �^Pz���bx�=Vk���C��q2�����2�3�c\c��AXGg6dyi������><�%!��]#|���Ly�>D[w��h8�x�v�3�β�L�f�H�P^������YT���n~�.��*�ѓ�l^����i*�̔}�q�j1�-�c��ib�]/��Z\Z��n0�����b��7ӣ���6���a�u$%FA峼�"�a���	_»��(O?�v�ȇ�r��u��W�$[��2��bi�`ڣ��/+�g���ЃvFڑ�-�Sb�H�R�/�����Nh�r�.�i�&Zx��I2)d��{=v:(EXNUP �����Ek�>�+!�� N�msHx1��xO�-��{�,IG<�U��F"Hy�W��s��}�e�'(�y�œ~n��I~ܢ�4�Y�A��꼿��X�0>��T�K�b�x�V�ɥ��"��o�����;D@3��B\Y]��5�
qT��{ �	����/�s����dc��Y�a�Ѱ	�xl�i�ܹ�ſ�o��5�(���
ʏ]<�b�N'������V��{J�����^�n�'q�>-b2�]DI����5��鹠 ���>-��^�l�=6�yBynw��ɳ%�J,�a��]�BmʗǊ=<���(�9�jʝ�[J�t�1/��&���Vr�G�?�dzdr�u8��B�L��,�������j����e9wv)�A������<�����+/ˍ�/ʍ7�X�6�|��<�N��;��!�'��]���X:�1~僘9�CY��n,����dh��b
���ۊX�tD˧��k�������{��*�EuR(�+~���4j��A���O�i�GI7�����0�M+�NKf��q������	,$z"�y��KF�o�K��ʡR��7���ͭ�1ܲ�.�����@z�A�E�ʝ�w#'���4��rsk�a���'�P�3���E��$��L���o�p�O��Os�"q��Ylk(����}Y�تg�Q21��rj�D�L)ںn&���i6�V�=�7x��"N91�m��,vk�c�Ҝ$MTK:6�%�������H�-<S�7���vO�-ߚ��A0�0���GN��ͦJi���$P�H2�b�ߒ��>$�<yY޸w]>�����/v�ʥ��?��Is������l\�_�o���7_ ��E��V��B��
iƔ2�Ϻ���7��SY�r�=~��	p��-�[��_P/��ʹ6��Js��D-��&�4vV���5����a���𫳐�X�R�J��+ȦU�ϔ��V7�yJv�{HǈC�&�V�R���f�4A�Y\nN�G�mZ��"�G�޿�ʲ4�]z�'o$&��BGY/��\�(����S򶅚��9�T>�p|�a�xx������Js�x4Amՙ�ϫ�"�ȓ2]�����Բ��la��?�r%���։9���w�j!`��]�3'�ǜ��BO(��Z'����Γ��ԴX�m\������� �<�ɏ��L�!���1��N�"3䄩�2���<W�`�m��y�'�*Sn��΃EVi�M��"������]y���r������}��_|]V���g������͛7Í�g�b2&4:��zI�z��f���ҒGw��I�d��#�
�7�>���@|���B+���QqTBI�?R��L��q<tp���i�h��ͦ[����՜{��#7�V��,�0�/�4�
R���
ͅ�������ĽY�-�u&�v�s�;OUu�d���5���m�5tKh�6�!�6Z�6��`���n��n�Ԓ��'QT��*�V՝��3�^�v�8�d�{I���9�s"v��{�oM�Z$u��56r��9U�d���[�mZ�U6d�A[)$݂���w^����� ���)�{�����w�=�LUe��JS��d�����5��\����)}���z^p�{S��3�WF�����k���d_�u+��,[S1�ZR-�^*SekXf��2��?�&�Z�����e��7�J����m��H�s:�Z�[�:��nȹ�����IvA	N�KD�����h����B�̚���N�^~��t�u��Dѣ�!=:8��nP��#��w�g�����}��U�a�;lN] �R�,5o&Q�[-X&��������_`S�-@�f��4�Ř	%�A j�<3C
��F�b|�&\S�G��&u��^����Җ�S��i��D0��`Q�<}��7k���,����5�rwT�c�����z�ϕ��*��!/y���"2����ֽ�����!����}�^�9�T@�}���J���,
&�
�h�c��J�W.>�tm��W(�ʅz­�5���}��vo���'�\*��s�����6������d�yn���J��'|��c����_�ʁ� �ˠ�f�FH�*Z+�t��+�_ݦY���GÉv�E>ݓ�o!GF���h贺�e�UL�N��2��y�Q���Q��HI�ߴ�QQw>�ˠW��I�����3����5���.<C>s�<:��V�篧�'�)Ҝ��ާ���,��-=MZ�D�B�jg�y-;��D��hȅ���2>�j~S.wq��F�Q3��}�n������ocLqX��#�|��W�2�B��v�e��?���l��.S0˭�E!����a��%����)��G^�HȎ홁���'-k�ڮ�=PC��~=�QjY$΁$�[�hZPou�z+�4a�ü>9����I��R�O *ټ����)fv��ј~�*nmoH@���;��ͱ�i 	�:̙gAUu����J���#���)Y
���������E�����4![ĠW\$濭��!��e_8�{5KQ�d���?ov������"�ya<?������ZzjEu��E.D;���W�Ậ����8U��K�I}><�,s�j�I�Ug�z��&Ī�d��a񓋙�oJcZ�(�6��yI�"~�N�T���4+��^-��*��I�)���R��[r4�e��'{����y�uG�Y�	I��2��t_�͛;3%&r+^ʆ���4�����޼DYع̭T�6��H�*e�y#��UZ��)�H7��_ ��Ј��b�R~�^g�Z|�n���I˟�7a�&$��ᄆ�������ȁE�[�Z�/�U� 9C��_��t�|��7nН;whZE�	���.�ή��$ז��e�C)�t�ҵ�����M����֨WyMGȵ̵#���Uf��7�F���EP��)��rt̟��H[9 ҝ�����M�4 3����*q��x�+l!;�=��B�R�?�I�9����TwRV��q�s���bf���s�J$n�r�5W���k�w'=����/�_7�߷�C�����?�h�f�?�μu�#+�����ҊW#l��q��E�߲8" n.O�}֘��D�7��1�#E����''h���5���+���LxA�U��"[�\��BV���_���F��J�V5��gW����L	�p��,�LUT���`˸��?T��N�}���ZH�x����&����^���{�Z2���{wh�����1"n,�Y��<GU"�UK �7��W��ɑ���~�~�������>~D9ꫧ��
�h�,��Y<�c��SmH5�N㈫�^���8<�f�!��e!sˡ�-���J���P��!AD��ҥ��2ꦬ��T6һ����7�R�UGL���fYҴL~͂=GͶH�4'�o8
���ԿY��\�C@XK���Yf�VՅX��-R��<��(V	z�,��#�Nj�C�}�	��r��(��g��B�Ru���r*��G��e�O#��[�9�C�y�K*���o������@������:>�hv>���):P�+�JxU��Erb��0���:��l+�
�fP�c k�|���SoI��E���#o���;�n�{�ta.|-���=�H�<�SCz���_H��`��<9H/��P�G�A�\�I�CWmݼ��)��a�K�7���t��V�*cάo�g������g�������8<!��GjZ�b�#��b=e�5�f�}�MqVzNp�S?�yyo���t���}Y�x�fr��?/�|�7�~Ջ+҂���n�L��PJ�/YES��Sv$^��\�2�<��B�"�:���|uq�R_(�+���>Q�5��Ul}%O#����˾�>��3�Ȥ�I���Qt[a�b3��A�l��������畀��XN���I~n+�Ԅ��67V�3��Yz����_}��܈��>��M[�r�vc�O��E�Qr���x�My��_�"=|�@L�t�dG��,���H�dDO����)��]1�f*��Hh�N,���R�~���/)cd���w豼^��ӟ�)�)���	�nz�{���5�o�\�$��c2w�>R��(��(6o�%�A}�-#�mHQĜۅ[/5��y����7[�6���B�����4K�Έ��?�4A��z���L��B(�]�}���es�*�ӌ���j�m�D��{��I����x̍�r����V��JtzOiJWw�A䘽1PY#Ҥ�*��=~a\wumM*�m E/q�䳢���;N\��h�T�k�C��>��� teʒ�2Ч�����M�nG��bZg��A�S{�ɥ#8'��VV������EYg��ރ`�X.u�A�
�d"�Uq�DɞN���42Mq��c�za�A��.���2G覄|V��?�;����\�-+c�<LA�A�.l�G���t�h�*_���7U���������l���
,�s�U����Ԓ��B-=6���Jl�[YզvT������Z���2���Rhw� ����t���h���J)D���,yn~H�q��0��-�����aQ`l��_LF����e�5t����40A�����yRT`M�;/�AUy^�#������[S�7��ʬ[J�m���`XZ����5��ݭe��^���I�:n̬�Ƌ
�n�pŮ��/I�|O�=�je��y�u��h����F<�j��~��{��[o�����{��$@���aH6�2�``�9,��Pj��/})��b_�D`��q�@q��*�r%m���cb&3�|[hjU���f��%�2�A�/9��R�\�s�e$�^j���9��R+���ᦦͥv���D����\PH��=}f�>��v�B���`�0ۤEo�cK�����s7NH�+��쮫�摑�qa�M�a������ʬ�~=��4�̔ ��4�I_�g]��e��@m!��N�Ő�BVck�<�0��T��K�ɣ�DgI��H�;��L�k�V	T:bU�'qQ����IĿJvn�)���L��Vh|K�7�]��X!���<���:Y���:�ŴВO���)~����>�Sc�O#�NXc���5i(=���\;��-h4���`��m�T3A{|��"?~�&p�p�h�W9zY2,3_sc�Re�d���p+K�8q�܏���:��~�#�^���G�b"�g�v)([v�i���H)���Re/㔲W��̑";Z �_;��ôp#-Un�:�l����o��D:.~���E�I���˅t�$�-޴Y���/4"A��P��������w=��{��	�����Q���r+��jYE�?SO��E(�*B��K)�4HY���*׈��6�QȻ IP�Հk��}��V⊜y��\H;:��6<�&Bv!�OZ� `�L��&�.�AI�h6�w]��ř
B`�"Y�gr�0�r!� �	b��:���Բ�"�.u�$��w�j�F�t(6N��O��/s�OHn��<�C��t����Z?�N[W/���ЭU�D�m���`P͂v"��k�zR���LKi��� "�/X�^=M�@d���;���e��y��\D�C5>�<Mк+j���T��9�AG _������}�0�C�	Q��L=�@Z�[-���̇9����j�rE�7e:*�:�&�\I ��]J�,�/A��kDSiJ�<m�.h��s����ο�'呼aP]Nk�At�����)D�E��s�7���G�թgn�ʟMkiuFS�cW�{�`�*< �"�2��<�6_��)	f��:)a�k�v�BZV�*H1�A �v�mm_o�?�h�%�|�� �cf�>YpSH�!¼�w���>By����լ��z@�L��+�ye�*1�+I,����]Ⱥ���	����-�v�,k�'p�����۴k� ��t�@�O\�x눭�C��J���������>m���SMx��I��:�$&�����
���^�K�v��,Wd5����ڦFd\j�k��R}!�Ю�d�L�s�]�Q�̸s�|�a�(5*�H4����(���-��9��`xs�>q��@H3=�	9M�~S�mw��,��8ܛQ1R�/�w����{T��1��A"�3%F�X�J���NA�u���E2��pp�v;}�J��+mxx����)H�Vd�ϑU?(���$��̐	{KPc��L�Y9��dJ~j����D��S�N��rвJ$-'�醠�|2��G�Tn�Z�y#߻��A�[�ﰬc!"�J��f"��q����hvf��2�gs����z�|��(��	b�����ڣ��(!&&5�s�<W��j&�D@������ ,}4%�ã��������ѢrƖ��D��h�$�=�����@>aǪY	Zݴ�7��J!�������̈́@@[�h��n�%��V�����y�Ii�Z[�d��y��-�s���Ĺ	vw �wA�*H�����������v��:X��h{A��M[�H�Ԯ�&K��B8�]��Y��/F[aO�f����~<�@/Ka6��֐�,X/^��G^}�>��K,d{���/�;����/~�o�%D��ژX�|-����~��������X8w!lLkIw ��\6�^~7���p�/<��_�������g�l�E�b�,0[�6�;U�s^�i�9�u>��~�~��>)���W��
&��g��y�t�ʕ���o~[��p4օ��������k�&d�����ݤ�;,,�B�s��-id"`5�`�d���н��A'���wx�%��?>LNm'�h��l��h}�<]�~�>z��y"��q� O��!2!�&{�&<:����&",&���u��İA:���M��������O��u��ɔ�)���5�_cu�╖���=��_bs�X�l�0���l���� ݵ�Y�̞��)�V"㝉�Q���
����.'~^��NƔ1�т�1�,Z�x�L;�h�~.��c�U���E���P�JZ�&�c�.����Q�m���8h�h�9��y�6i�z�J,�8'�P�3X����R��Kq�蜗ń�O���@*�kk!���A�y������k�֚�h��<�#���3���F��ٞ�g:�Ӣ���i)�:�� y�`3u{���^���7���4�����'?~��рNX0ܺ��~t�=9�;�]
�vh�� y^ӽ�v�����I7��(��M�g��3'���d��.��Ȅ776�h��F���,�6c�	����EX���&�d��h��/ɂ����]z��o*Bc����A7�� �������1�o��o�������:�k��"geD+>���Z���J5��l��/]�D��뿡���_�roFJE(D7�!�A���� ?�Ҧ����K����O�o~���PZ��^�%�xΝ��/�ǃ�d����d@����}�o��5׀-PzP�jZ���h��_�}�g~��<�`+������R������	��*��
�v�Ok+�����O�����E�	��F���~��3��s?�s���}N:4r��VH�Li̤�E�h������'�����ʡ�n|��T�l�aHJ˭���
�w���Ѕk�������p�Hr�.?��Y%���p@?|��������D����A�,�5�ϋ���?�Z[�	X]E�����?[�bi��V{��|g�������+O(#Tn,w�2��Q�����������_�,�x�G�؆U,ܸƑ�u����xD?|��E�$�)g��T��L�t"Bd"dɐ\X?�Q�9u�� �����M[~tz=ZC0���'��t4�6:�=O���>���;��[����}2���t�'��F7_���"h��L����D!����bǄOQ��_<'��g^�I�L�'��XI���G�sh�t)�A(��j�������!]�|�ַ7e��R���0JW��M'��$�t
mA�������B���`Zj�L���.lӕ�)c�&��w�̑H �H�%/rCÅq2��ҟUh�B��甅���F�^{�%j]��(ঠ�:�����'��F�v+��=���?�՗�+�u�\����G��4Ĕ�/���]ߦ���M�����l�&�����n�%��MUSAy��c�<}���"����L��1�>�	���/����Ư�c�,Y���ĳ y�����sTM&������M_�җ������k=��<��_@���ӟ�(����j��I��`�l�iT^!G�PY�������������ߕ'nY���aW"��Ȣ������?��u������oUzJ�W";��o�B_������ޓ�����&q�H��R,����/]����/h���5F��pD7�4S�ш����У���ѓl���p�������ǵ��CĞ���0O����Kk�{m�k��2ʷ�ָ`�9���G����mM$���`O܁8�����jm�t����]�񢠎�� ,��)]8��qӱ�)Oo
u��?H��u�0��ms� O�-L�0~k��7�6簙Qb�T��\��ʡ�)#G�t���Ç�.����>]�z�ֶ��'���N��(`B������6����"ؔ�:>�7(5�x����ӓ��^꯭Q1'Y�!�h3���t��+����߼�.���rnAhQ�Yu&�0�y�n}�>��i�Y�};��<-R�Q�V4eU�":�B�Ί �}F��^�Q�
[xiY���_k���#VP���/�kluuV�1�Q���ҹ�lKǌ�4>�8�	��'����֭��A��˺E�����<�=�ş����Gh�f�	+�J��h3��enQV�'s䤯�U2��2��Nf�U���@ pt|H������E:8:�����ȫ.�X�P�8�V[����`��fS�bp�3f�H�: ��2>�'�n3��P�'����tN�b6��O��"��|��wS9+�T+7w��4�(ϋh[�W����<���}�xn�Хxb��đŠ�b4{(1�u�O���
�O�q� ���R$ks�Ε�s��%eC)sTLA��aӀ5n�EQ��X	2M����N��e�_=�J�Y�v�6y�y�vxһ+krS�ߣ{��Z�%�$��i�R4���ޖ���G}-� |<1��nSӞ�@1��H�Sm|iNh��>�,�:�q(���7��w݊#EҾY�� �JD�O�� �?��G�_�A?�����f���6�i	�=J��?���z���
#�c�7 ˌ"*�rgV1����n��O�����|�g�j��X��f��ق=T�)�F�� 4!|��w�����A�kt
6�2(�+F����;����_�%�t�0�ͤ��D���!-��\�h����D���_�=�͉(��T�阀���*5# ]Y鱀�g��6���q'��pKȽdh�O$A+E<�H��yrȟj�%f��9Z��bHڶH���(��t�����+���v���Y���B׷.&APr<�6��}����DR(F�Ri���С����w���i��~����ٻ�:��jP�����'��f����/�J ���w��mo�"�y��HA�n�>_�Y��gFĮ�8S�,=i{c���?'
�p0�.��AЭ��X�s}����ʸ�T����%���,���&�-�xn��ʾ����!��\0�{��t��Rd2pY|��sey�pM�|�o-<k��A��o���18�:��2���g>E���Ͽ�����mu酗�Є��Ν�Z��u�q���k��Q��!7/�m%I��xP'`�u���Lx�KJ�j����1��-X�q��ε,oR�Z0�K��J�������U����,��sm{c�n߹E���DY=z�X^��Q0�N������FO��͗^���Tq���<��,h��e�'��uE���;{���1�$��lndT����Z�P���)����W?Jo��]:�s�ϑŒE����(�U�z����2�n#d�ɍh8��|���|\���f?�0<�O}�t��ޘ��3��%�ֹ�ri����;��ߢ�������ӘZ�ϱt.m����X2lڭU�����ؒ��[b��>���Y)�qFv���w幠Yc.-�3u�ZA�9�fE&~�i0.X�}���k���7���yW*-��a(^�v�/�Pܾ�sYJz������bd|��Mlt��76��u��S4z��Ѕ ���_�{|H�>���M���w����_Y�ѐ�1*� ry�5�!m���o����w�|���?|Y�����^���sA�w0����ۥ�	�hF�G'"�s�c}*�ѕK����ߠ���7�����%��;�м�5��9e3Mi��Ǥ�	��um�je�T03�Bz�æ�^<�����f���%ɡ��/|����o�΋a��p��Y�uh{k�'g(�RJUkJ�8��+�ڙ�:"��Y&����bm��<UΚ�~���"�U�W�l�h,^��2�נ2���b�V� s٢�I����ի�3?�	���ܷH_��vӌZ�����H� $���X�ۄ�O����dwW��.o���2eB�j
��wJ�)G������+�Օ6�~�(T�r=��n��Y2?��р��Xk#b�XX17�����C�J[zȢ)o,d^ �P�,�Ӗ[s�|ª�*a�l:���_Y�����FҰ0�{�I��D�4	C��i�㚈���Yy����t��ҭn��V�Ǡm"�����"%��-�6)؂0ș1�� SH]b! =L��\;�{��{@VDY�H�[�J�HWK׶�Y��W�C2���Jm��ۮ�bUb�a��|<�c��;!����-[C	Zͪ,���ed8�J'@,_��X�4�B���X�ZQ���]�����o�s��
~\�OAP�QJN(�y����O�,=~�K_�����+����m��1�&�M�k�Z�8���A������׀{@8y�N���������1з�z�'e�p|���
��zr��Pv����b��k�[���I�;"���$v�j���oŢ����7�7P-�7=�EK�P$�]$��U��x����.�������5XR�({`BBM�U"��J#�S��2X��F� ��@�9ҋ��K%�y$���K/Q��%7��Ps�A��tʦZ�]�Uz�wHm�*<�Z���F��E�6T��"���cj�Whuc[ƙ��B�)�*��}fY@�NX����֝{ԻpY{9寖��+��i�G!�M��=g,�;����#���Őe�[
V[�q���-Bw���+�2�2D���s,5�V}� B&c��3$�-3N�@����ڡ���H��� ��-�D�4 J���{1ӎ��u#}x����Ǌ3��Heૌ�Q]H�u�B�:+lq�G�؀�A3s�W�5�>�JJȦ4�>��_ni���H��۽
힌wL�e#Za@&�e�dR�FZl!"P!c ����;�'�˻8�&�|/�<h�����k����*�
��S�"ISʰ~�*��w��?�^g�Y恼�8�b�F
���&K��3(ۏ&�'� r�T�"Q��S�2��O�6�b�UZ�#-�+�5b����?��M��jO�j�U�����Q��$AA�R�iے{��E�˦�+'6("����Xe�2Y4Sk���
�`j���*,d���ltE��ܐ�UcqŸa��Y6e3Zl���/�D��e*xm�i��Ql�F������D����8�;�����x���O�_K��E��;�"��|�X���)O�$A����eSuumCHɇ�P�FT�e=zr4��{[0�O.�oZ�DR���4U�S��,��$����z� �Ye<�p�r��v�p]�8OEw��~�6u���:��嗨�D�%!�,C�s6jT}$�uV���E�� .P&ʽ',�Ɉ�A�u���I뗯��`Fw��	����$Y8	�����$H�6�*���ZBŚ�	����<p��.UN��n�	?�ۏ��:'2l�Y6��P�U"�Kك�����rk��� t#��Ǌ.��n�ʩ����u6����!e������Q��B\#(J��uk�(�E�[_g̲T`�V���t���kvek�>x��wL���ڶ�p�����q����*+g%Xd:�4L����6V������+/й�����G����,W3���+i4K��z0k��ɘW0��b�Qۿ(t������6ꥫ��j�	ڐ�kV�d�81���J���:mk�,)+�TTa���8��+_���G�t�5�O���V,����Ā �޾����בW���j�bŜ+4�GnIα������$�-����y{6'd=��-���#�&Gӵ���T{�E@Mƞ��_��Fm�*���X�i����=,|������}muE������Ts ��h������pNl,�M47^x���У�c�mY���>�OvĪ���z豙�Qv
a���N��	Bx����J�%�2H�K/� ��%b�
�~�?x�=A��!��f��08@?Y5�M���`��h,����,�7��ᱴ�G�j��}p��e���4(�8�<>���[U�X�e���z��+A�=��-�	F�2����c����y��HL,�_(s�Z��0CKI|�d�f<�CF��i�7a�`A��$�����9�������'�Ǟ�3 jK�j�.\��{�X�D�����pw���y��r�~K�a�ć+>gMND�J��퓇<����K���T�S�H�Y�Ӄ�C�9Č�"��tK�����8�,AO�2Ӽ]χ�ۧ��σʟ�ʥ
��m1rfpƿ���V`-t{�l����)Dqa��mx�	&;�|VZ�3+����P�m�Lk�cmX��_v�"]�L،@=�uʎKA�S�hn§4v��M��׿Q0�~�#��W4���!���k��<x ���7��ӓ�]Ax����E��G�N�FN=)Z�c��S�l��ߤ��<����a��I�����V��*���
"S�ZlG��Yi�)���d��9ߕ���(<�?��?�|T�$�!"܊B�#@q1K*���-�v㺤;� ��r���#��"y�_��Wt�3E?]�yy��_�_�N$��`<��I� t�;g��TY������ث�I~/�ğ4���W>J��ݧ�?��oO2$x˰e�����^�{��w����3���drlU��e���Wip�ϊ�#�|~}m�}h�+j�y�p��ؐW�p� $����`��,�l�R��E�.�q���K�DIa���E޾}GKrlda��1�VZ��kC^p%�G3q��\z�9a�by���trG�n����[<�~����	�_���{Dּ��y^�`��{؁�CbU�Y�����ߏ����&M�}��jք�E�/`��0 �X�C�G0�e��������:�(�FP��ҕ��B�"RmAx��>ޡ'_���+`qa-b���mYd�d8��ۓl'�_��������H�lt���R!��n����%�b[]3}���<7UL�R�HE@�t�"V8 ���� �k�.ȷ�v(�8�:�wx�[����8eUP(KSG��L�[vMXYMZ\=M����i�w�
����w-P$0qd���R�-e�.�ԲX5�������ohb�RL��lT�?�&9A@q:�� J�[Zu�Wz�R��4�<O��{��V�����WDp��y�����Ţ����3�����x�#���e���`Y�F��#xV��_`��	+�cT�LGR	�����?��?/(���H�Y���-�_e�_��LZ�W���Wv/��P������m:���o7�ȼ��C��Ch��H4��M�ω�H�	^�:5�B$D�_n AlSz�c�{��޿u[KC�9c;����R�S����5{�HK��4	�,��|V&@έ��:4"�vN�X ݹ�H���?ٓ=�|V(ʕnO����2��i�����k��)mT��:*Z��Vum��_�L���mQڒ���)�O����~�L���M�8�㩸W���m,[����6Eɠ��Ռ�=u�����}V^*P��B^v:-��UW����PY��/���Y�������U�����	�S�S�q�cM=�m� lK>�F^�\1q0w��Ӳ�G�WO��٣<A/�fajj���Ap�T�����-7d<Uͅ*yr J�ŋ�,�Y�$_��gW�Sm�L��ɹT�UT��tA��)�.���P!FSe(�3���	��k` �iS�;Ll��}F�[�k��h큲l_:�J;Еѱ��%����yԪ��(Ţ�7V)(���HQ����Vn;����ʠE�}�k�p��>��,r[a�WXHwx�O'#e]���^wYxN�������]gA�����My��`4�1(GishQn
!.f: �"  �*
bfc�fV� �"A
�WP�%$(B��VB	s�נ���_V�6��\������ofUr�g��N5~�y��oHm<<��6�	A9��DQ�7\<�����)�k����\}Y.A�kj�51�i�@�Nr��rN(�iA��B<Ȟ��yLb��Ab,KL���tG%��x� R	�C�	3�?���H�;@�_�q�\��tW\� ��ϋg)q#�S�D�3^W����������L]�Y���y�^�-G�Y����!�Dn�~)�z���p�fe��΅U�b�� ��D�����~��x@��c�8��4�S���Tt�J`m���j��k����J�Cq�g��3�Ct�.=�_(����9��!ޘy��T[DT�����sZ8���KP���3��WyN�кBt�s�+��P"���:�'�C!��l�I��H~�g��O]["���aL(��s�v[�¨m��Rk��V��L� g$��RFP�jv��@ݥ�G�51<s�6�	�%��6�ws�O�����tn��x�K�Nix�
 �@���\$� �㣁����l�����%/.)7�����3���M�Z�����P��j�&�#��0��a���p,e�EeI�梯2�]et	T� �:�.ȟ�3b��l��X܃�4�>�}�vF�U����$��O0��ZSi�2B�4�|�)P!hs�4�^�[��o����6�g��k~;i�^�j6�tM�T��n'
��x y�UҠO�Z��⚳�zQ\#��N�
 �󣓳�C�u=K���v���j�zE�89ָQ�ov��q/P*u�,�qPJwd.��b��)��%r��
&�2J�\I0"�SQ(��o�!��B��h
��d�4>>�"�6���t���*�zh�{�LS����-©�	^b����И��o�����9� ��l,����/}��]���F����I���J�6Y�@�n0�[g�h�R�*�|emC\�̝p�E��ߗT�A��πo����w�zH����V�a���u����� 2�
\�V��FzH<�ED�?-�������:d"�=��js��]Y3@��+����+}��7"�LU�\�_+��PS�z���;dA7F(���9�;��la)R��y�=����Mˍ?��{ěAr�"��KĞ7-h�H���?>�<V:��,�#$mL,6��q�P�d����˫�'�^&$�"ؑ�@"�R���R�N��L+��<��ĵ��+�B���h0�٘A
��r<U�5wG�H�t��F�Z3)�!��ϙ�۵I�%g�f�=z�(��$�6fT~(�* �	�T�|���"i����(�$厪zh+tX8�q1��ᱵ�M��x�-l	��G(�A>�x�]�!�C%s�J��B0P49MZ��"����-�P�>'�/A��	J7v����r���ښ �><A^�I�A.�	i̮�vu�6���C����2H8�E��{�PU�(:����bJy~�hv���8�tyS6�����φ�ە�.���%)Ǭ�S�,O��ݾT�=�q��V�\5�l�~�DQ�@���_���TB	����	\Y�9�Y�77����-t��v�⁏�w�?D���h2�M� ��ޮ�R����Bg
G�`���w�+s
�+H��r��Zg��������05�%�u�� NX������m��@���wh��(�}PN�,��+���@4������u�4�	����<~H����� ��u�?0R�2�n�A4����q?���z|�#~\���
�o��%�T��}�|���%�=O �̊��[e�G��uY����GOb B���t����w��=���\.��m	�[A�۵x���AP��J��Ahu�����vP|�\�oݲ��X�Y�X�<|�B.��
��s�[b���SH.�ڤ7��Rڴn+�k4�5���#Q�P@��9�f7����	�/�A���n��WQ�$�"�W�ց�3��\��3���Db7Z�����i&�r���C(@a}a
	A[K�u6����YK�|&������@p�t�����D�p[����J���HZb�T�X��h�jZ{h-���ҙ�K����gCy�fpW
Vm��]>���6Y�\�|UM<x��U��YG,Pwy�`����7������t�����o���G`� ��#ͽ�0��L���L\�v��Z|Y�����"�Q����|�E&���������j�l���\���.Tn�_"��o���ݧ�	䕚шvO���� �%��s��~+��Čg������tt2�T.�-����M�n�fo���@j�+���%�6�i��2	Tj9��ގf��(��
c�@��y�HkC
�L/�@@�l1������@�},k8�Es4I�f�mk�$����fZI(����`p,� 9�=�#��� �����1+	)Bԯh�7���ɋ��>�Ϭ�AMiGx @�C������Ni
V�6]�pA�4�,��	�[�Zrn���QP�u���\��=-WRv�ca��& Y�e%[$z��e!G�w���oD�w�э��94EE����t��Q���;�ԝ������$Z�JxOϤ"S������^���=)?����N|��%��<�5YC��{(���:9�K��<PU��@��!C���]���/���m��� (��L�}\�`�
z8f�����p�.2���\���m�`�Hp�EhI%��f��T�#��(����f�8�5��h����1w�TAP���l��������4W�na�'km}Et>7��#Nm���H�'�/4�^����@O���k�'q9����f��%"�H ����WJ�#��S@��B�Q9%]5ە�����N�R����K��r
	 u����U�\�H��y��j��ح�9�N�qws��T�K�e��N����	hBLC���)��A�5�π�!��2FQ�D|�� ![iR|$��*�.ˌO��x����*KUau�x7ȗ���	���iG�R%"�}r|b�!QL8dm�u�֖��m��:��|�ے���ն���	�H�e��'�dwOy�-h����hY�AK��g�$<�P� �F���h_,>"M�t����)���W����r�p� %>^��w]Da_?���?��[��
��p^��\�ueOIg�c��߽wO�-q�+�Ha\�i*��O�g��$�_�|��2�F&K�L���Vd�� �'���9��6܃�1`p'��o���&�BZ��wp(�������5���r1$�Gi�$y��ۼ�T|��-���3����,���"=���(�C�H��Dh��dM?.�R�"~�L��  ٽ0�Ͱ��*�
FLz��+�.�qB���y����<�U^�[ۛR�{ tf��d���U3	��,4*P�!��<�Vw{���o3w$��YQR��l�k=�ў=���/]�IHǝCa߇i�wr�P�Yb,�^}VB*܃0Amlm�� ����
!
���!$��]�6�"��*������ں���?A�@	�
���+�� xSTb� �aj:l�����d���8'��&��@Vt�k��� d�P��\e�o�����@�ީ���u��0˃5������ �7�y��O���3���vߡI�%�8���B�T;�\��#����)Eg��H��s�$[�-����YaETщ \k1�� CU�p�"�~<�ʳ�>��M�XQ�Ӯ��[� _JЙ����^��at�4��X� :���l���({g+��ɚ��*��՗n�}F��+�2�Y'�5�D1����%�f�rGw����*�J�\Xc��A�[ݤ�˗�� ���L��bр��;W�v����r�:�f��9㥬 Y��������<��խT�3M3A0����Ƴa��M�gV��n�X�c�;�<���h�J��Hqб6�s���{��X�f�{��ز
	hf�l���X���,`���s���!x�&r�Ȼlb��2ϗ	�扅�6��Hh�X[A��.C�y��{�Cr���"�B5��g���K/��w2A�Ǔ���\-p�#�C�MF��}^�G'#33K�E��x��E���O����/ރ�hRo������^[<_�#:B�+���k��֍�К��$�[Z~��M�r�J���B�K+�LSP���fg^���D���y�������V?H�&u���:y@eLm���g H���hW��T�v4�E2 �5$*������t�P�9#m��C�[��}����>C+�AY����Q�kd �S ^(�/?Q't�p�?�;B�< x5U��kE�[Y�<m��y�Z�{{�㗼UV�ₙ��k�5��퇇'���EA��d���s�hR�(����֖<���>��YN�q��
�% TҘ�����Z)j-���e!8SZ����ec}C��^��ñ �؅tA�3p$������� ^]���x���Ub[��0�p��TU��M.GRo��{�p��@V�l����
`>4�͛d_2� �+9��B�ϒ�rbS��Ȼ��A`�+�M��@��ZYQ�6<���!�8��6�����Я~�W��oҟ��_З��5��Y�h$cv��lY���L�j�4��^p/�/8�iY���˝]�5N�?�EP����겄]�:���N��'RH�g#�43�IZM��Z�ylUy�s�ʜi Sxc-�mm�����R�z$K�3�}��a18��4��H�%k�(�sn[�A9т���Ee����Y�n���6��+��q7�����	@iԃ��_�q��Fek����(���4�cb��d&��F��j�Fay�x���;q�@�H�5rf�ė�'Bb�si}�F������<�L�$,��Ԭ!�ja���#�N���1�I�h�i����KI���C��+T��y�.���A�e	���,�
k�M��Ժ(�R�p��K�+���������u��Cf����w��)�t��=�$Xu�P?-�<�T�I�q����ѱ���G�R���y������7�l�������xs��T��&>X���(���{ ��k�|1ݜ�;b�!�������i
A��A��1��>!u��F�9rAW�hߊh���=أ������%���2]EW��U�Aۖ:'�`��4]!�C��?�
��ų\��gDw�G�f�T�B��M]
�@�O�%h�Ģ�8γ�?������nF�h$c�멛�孰I<��i"�V��|�y�e���3e�ޗ~ފ\2� >R|Ϋ���͛�F��n��l�%� H��qZh?&��%}�'�$bF�jB�����~:o�f�������G��Iu"�?��]k�2�����F���G��ik�������RZB�f������1vb�o��f֮%�zϹ�p*I�+��<yQi�T9_,�K�/k��U$�	R���,�"?ҵ��D���{*�u�%�ٹ@6e�V���@�,_UU�بg�^�"x^� J��UL��=����ңU�!-kW�v�5���#�`|�2I�.`�*��d���J��J�V��3�5�>�X�A$8�_ަ./�"���QHvF.+�/���ڊ"< t�$�)��A��vA-4}��vXU��1a����Y(����/R�Ёu=�}�ΟۖM	����6��x�j�L�2�%���s�E`���zd�陎��B�k�����@!	���	x�vh�եK/��o��.�O�Jrcd0u���43�"'*Ž������T�؎����S,���M�ڧCY���(*�`�ݦ2�7�T�̷[h��J��!�hDI�:���TFy����f��+��[��<$xdi:i���/���dV�#h_l�8
	E(�0H������~G�(\������0!��8���1�〢p_��Jė��s_+��AU-d:���ߕ�I����^��
X�)!�����%�?Υ_ó����
��^\x�2�M���P��"�-9#�uMp\b�0$��>_���{)/��5R.��uJ�>�s�M����6��O���!���
Y����*u!����O�l��5a��w�Mb&�8�0��l�3I7���=�g��G�V��M�&@�	(=�p��E!���ʲ���=�VN�!������OZ���<|H����V�~㆖��d���^���I,�'��n>�R�`Z`�'hT1g~���<Z��߱p�ic�?�(�n��@����Q�m,�q���3i�c)���{/�k@�VQٌ�� Ӳc\m�K\,�X�)���Y���%7/�]r��Bm�(du�x ~xi�|�:�͑���m�����!;�$�c���R�Bz��suu
D�JW��Jc
�����%�ꙴB�U>�2ZC0A��2p. ���V�5[����ƧF#����g7�|V��r?�r�nkd��#�-5�����e�%�?���5~��h���H`��w7���cT���a�G�tT�J�w���!k-��J�n��d�K��d�C���� ����� � �`
	�"�y��B���R�����A]�>di<@���&>�6�jg s���Z���\��,�	< �,e�
Zu#��y*���OW���*QmR3*O�\r�A��Q0������Fz�����/�s��}Yj��M�R�Պ�(����Ӊ�3��!�Y�t��u���ģ-J���I�{P���b>�0Sd��!�r�db+�N�n"Ϫ�a2�}fNѲx�\��L�h��U��`ͦ/�-6w>f5߯Ͻ�552��&�62����aѯ�B����\�Y0S�JD����Z_K��畮��A�Z��&�$ч�\�M2G$H#B�$܃�ㅶ��S����U4b�O�>����E��LD��{����Ayv��Lf~���3�+���H2z�&�(�DR~���F�;.%��F+$2���ʫh��7V�,���m�z9i�f�f�}AR���E�W�J��=�&��/�Kh��l�����}��؈�������#��W�O��2^�P�W\F!����������!D؅V���mM�n��4���s��}����	�M\W���5������ye�EP#�@�B:c+��.�[��-���Æ���-�'�`*����^*dI��cU.$,�A����_���j�1'LCI�3?h�%� KN����~����K��������G���岢��h#Ѳ�F&�V/^�� ~��#9�`鰦h���k�a�|�C+�~:�L�:Z�������:I�h I�'y�.z���m��*	tU�̵Ր~�;��%s����K�g��r�l\ �<�&N���X#��,���Yk&�h��c��v���飰��i{�^&$"cK�I���t_m����c�3�a�շ;53XS�օ9�8�>&����W[R�{����8G^���t<�Z5��d�uv�������'X D}��1o,�Ļ kr3�O�`U!8��2n���J�wQ�
3�D1�_Nѩ�ʚ Ư�tN�D��xsq��g! ���~j9��^��D��?r�!��|�Y��/�Vʱ-_+ ԟ���P2�,��8/q����LX���ҵ+��B�'�,t��T߈ϓʗ2�Wx��g��T-��!s���|;ᒌ�����[��y��9�����ѿ�ҟ�����P��k	��
ü׺~gA�iZm3 䖡%�k�������jU5��>56}��I*kk��IH?Fh��a�C �\J��F�I�-jM�u(g"Tѿ��o���ڦ|FZQ'�X���{Ukçi�j��%׉��Zȇ����U��`�p��VY�
��V���i:[Z'N���Rg73
)��b{ͅK0BʕȀ2��l��v4-&CZ���Uz�ïҫ/�J�|���uA����D���݃t&�甙o2z �*��J�[e)]v�	�������4*d3�P�؎F���V|���<��3�����;�zYDX��˅t��*)�D�eA|�(.��N��O����!���Ƚ���6��
p	�:�7$�y��x7�ck%d��z�C%��i��{�LG����Q|����u�m�]�7��"�>�K�	YT��cV�[�N��q���kn)Q���7i녛͖��:�Eɗ��͓��ӎ�(9��ه�N.�h��g���f24lf�xG��!��7R6vLz�(\|�#�C�0Ļ��mj�u��Z��H�x2!��xT[�ۛ��y۲
�yd��#��}�5WϴBXtf��v��ң�p�:��m��85�S{�4/�|��*�DһK�T��y�cC����M��t�7��>�Q��_�u���Wy���i��%���3�,`V����yJ7���L��r˄jw��<o�x &
���0���	�k���PGV�@Tc��d���3���7�%e���
E�������μ�E$�n���Y���|�n�8��_��Y*��"����{K��/��>H��
J^�Z^!o.�T��2í����+U��5"��0g��"���T�z�JO�|����B6F3G$�K��K���Jl�9�I�ђ�iP�6~���FA0�S�Jޫ&��Z&)F�m���,3M�ӡ��.��$U1��A1�r�(ٮ����M��S�.Ni^H�O�M�x�כ���٥��7h<��|&I:gː���r��>s����T��!�T��`BV��Em�ySd�T�CL���֛�����Zi���W���W�������c�}Jڃz�UTw�%]S�\�j�eVE�F���t*�XY܈e�U,�q?���t��I��1w�~	~�!�3��m����@�"�Z�*�՟���2�D�_(��X@�3�T�"��?e��Os{wR�`k��r`���N�uc��-Xf>4�m�Z�����+�ek7L�>3t�k����N�ѝUͻ��Za�{ǟ�e'����@��YY��:�c-[[��,XHfu�n�]`�^oBMpo����\)|sKK
�K](�OJzn��Gm���cf�|Ǭ1���8z�FV���0���˸25=�\��F��Y�����(�.��!ű����F���wG�τL����Sl��-�p�{�T�3��L,/4_�ϫWƔ���s.Cj픞�e7�K2Qn�*Gp�x�1�k�b������F�Qi�ɏ~�>��O���EP��s�u}��ZP�;�h>U]�9�-y�s+)��T��sU�,^��;�ʗ����ρNYF��-�^zds�欨�꣒�I�LR�Ƙe�zf��-� )�"˟1�/�t��^>&�}M�9����3��M�B8�U����b�z��~��%��yZ��G�#� CB�R/���AU��2��H�N����V�4�y�$��5�
��Fy&����!�k���T2�)���e��E�c�$
j��e��ZM���µZ�'W$Dt�.�e�6A�Q�}4r"@��Zոӟ����+ ��8����Xb��f��v�h�2��ƣ��������W?N[��T"d�����T@R����#�}`~��s�e�'�n���;c�!Ĺ�}~]4�3��%�s���_]���%��Y��X�q,�#y�Yרh���ҷ,w㥐��
�؟��B�!s�Q��T�3E���m̂:�S'x��!x�t�\B��An2k�v�ۃ��I�e��B�m(�<�bCX�@h��l�m�N���\�@��,%~<���h6^���@s���t��P#57a��<������в#�TU�A��>�)w�J�$Jwh����/��y	�b&�BH�ڷ7�Sb�#.��U
C�<����(i�k�q��Z��9|@�����g���x���.�iC{��s�߹���8aE�5�8�l^��o2Y�t�a� ���z˜�Ҍl��3A,�c�_m����͓�S�7��-�[Zz����{�\�ڿI)
L��j�!B#�(��_����/�A���ܚ�'U,��vYYB9:0���o|��&�|�
�AU���Q�BӅ�����h(g oF?��� �I��sM5���b%��eGj����{en�Z৲�h��'-A��g�
��_��kst�ƮS�̟d��֞��cVH���/˜�g�	�o"w��x+�<s�ln�S��X�|���8��|4��y_wh��~e�5�/]��!hr�Ui>��-;��Dw��+��Jx��"&�^&Y:�xo�W������I��Y��-;����iR�i]��\���T�@�N�Yqm-�JS87���V� �?}P�C�Z��������!M������t��N|�Z�a{�`Z��Ա�d�~�$��®e}{����/aq�i^j�Q )٦���8�j5!��ZPp"���.(����ڕ�W͖t�vE��t�(8Ψv��'z�2��#ờ�#�UK45��'�i��������g�j"��t^��Ĩ �-_eű̕e@I�1A�+�H�2��Ƀ'ː�G}|�v�jA3T�&^��o�t]���Y��x�H�hF�.��p��%>I
T-�P.?S�ȅ�L�9-�Dq�E��*��\����c����<��:?�4�����u���J����ȟY�FY�|��}�z]{�,Uz�~_e�i;�WO�l=�����&�}��!,;O}��z�{�Ϫ~K��~U���yi�����Au��ʳ����ekӭ(�o����TF�U��D���	ǖx��.�����@��i]�a1�4�˻a���Z�M]^�F�.y��Q�A1��r,�1p~��Hҝ�LٙH�qe7_�h�囼��B��y��o��t8�^/�q6�<6B�F��Ah}�^��UDE[]���{�#�n/I�6�#�~[3�V)h����#�*�H��lA]��\�X�th�����Ή����MY�QSr�[��]O=���O|4��)(���(d�}�"�3�I�@E�թ����jͺ*��Gd��ֈd��.|+G�K��~N�yj����BT�t3�D��%8��Xv���֩a����+�Sh)H��l^�>�
��͟c���t?��E!kB2�-��?�K~O B�?ҩ�x��6��e���		AL?�&���]�7���b
���e郚��]�#ʿ���B�'�m;@Y�R�w3SR_
�e!��h<毡�S�Y��d�|1kP�,�%�9��9>�&����4��~>�~P��š�������j�&�C�h�աrwѦo&���II{{#Q 9o��V�>�ᗤ�����?<��1P�
~�y��LE։Օ�B�Q[Y�$TAe�yϹ�葸��Fسϻ�~�χ�h���dVÔ����zP����H��w(������D��3
<ر�)k
�R}��ް���T�>�X����������ߧ����y�g	�=o@nq������K�z�V��?�l��g��Q/c#O�9
���nNj�}PQ�/
Zy�J�Kg��y�X����uF�[����&u�ܭ��.��a���v�k��txtLw<$����C�*W�vi�cf>��b�8wk�.���U��_����f;��Y@2 �Ƒ��Ñu�Jk�ʃ��1���EE�E���|���{������R��c���H����>uz-��<�Cp�ʯ�6ᩭ�����q���`���Y��0�{��ĢI���(��٧d��M�,21������!�0��-.�0G�7�f���c~Ju1����	��ݠM�f:F>y=�9��44���1��F�]!�`S��&��Ɖ�#p�k�%���< R7RSa�|�D�q��+d���1��z�1��i�3�'�I��ߋg|�,���e5�d!�f^*W��p3�jSʷF}>���q�#���.O�:�4+�����>��y��6��K7鵏|�n�x��66���|��ƁF���s��mE6:��x��V*��P?�I����@/���2F�m�ͨ����@�hO]�2�Ӊ��F�(��ҽZ"�Ŕ���h�?�ѓ#�ʃ�j��]g�7���x�M&3��V����O�� !��m��N��	�Ғ�5����J����h�:��E?b���}����~B����xҠ�ұjd^xU]vJ͍I��MW۩��y�g��u�K�d�ЩAȫg�@���ދ X�R΃>'t�*�t|���c[��Z�����[v���zz�U��秝s�[���� �~ޔ`��GD~������}.
���w�4Wl,"�l��V�F{v�}G�ud���Y��o���&m���ل�]ߺH�����g>�Kt��M�h����׾F;�����S��K7JxF�vA��ʍ�t��6]8��i@�!��;�����tx�\@��NY1zԃɾ���D]B����{ڭ6c���wY�-�ڐ���\���{��g�{Za��� ����`�]�s�}z�_( ���ҹ�usA��P�Fn>�N�����ږ��~���̧G�j���Ċ����g�"J�1�z����!<v�@���7��zZ�y��5Z��g��%�*T���M����(!��:WTč�L[��صߔ�v��T�y��-��_xos^��>��V�g��S�s�}�Z\T�����g�<�l?�ߧs���������dU��WU�;��͔j�,��}=Kx�P�� ��]����@c��D��"���.ѯ��L�~�U��-I�:�?�����з��-[�"�\MhX�&w�.����c�h����?�!���7�����	#�k�.���6ݹu����49.�c.Rń��� JK�hY�n���ˬۦ�jO;{�х�$�k1��Ϣ\^���)�}�����Mz�`�F�����du�C�j�_⍝�#�Qˎ>[��K�0���X��yͩjMs��ϔ���8u��V}9�=�� ��տ�}�0���H]Ⱥ���iZUypx+h����.��u�G�ηOZv��L��~�i�w��
i��Oo�I���Q#d��=�bZΜ�#���/Y��͏�7]N�	�Z�K�-6���>*Hۗ����+�}����ߦ�|�����@�{��94��҄���lD�M���M�&:G�ӹ�F 'tww�������W.҈��#�5*;=�t�U:޽O�d ���/]����[c�[���}�n��>����{,d�BD���X�cT?S�o���R���a!�y)͆�h�Ґ�i�Bb|��s�x�N�Gڰ�߻��--o@&A����Q����ʩ�זJ���!�������~����4~O���"��hq��"^8�]��z�8B���+q�<Ǳ�:Ü=[�2��$bn��,YM?����B����]'E�� n>���}=���<�=�rDƱ�|���i燀ul�pV����>�e�2E���=�4R��d�#Ɍ��L�"�Bu�O��k;J����m8�( "����DϦԝ����  ��IDAT��~��n]�sk�҅k���/~��׿E;�����U�v"��tZE���N�Ƈ��o��|��ƕktt|H��/у�wY���7��;y�l�l��ݼ|�>�3?G?�ۯ���;4ㇴ��M��C���>��O�?��������%��?���?���]��z{��]�AO�?�l|$��ED�Ƿ��t{}��~Wۓ)	�eF���L�hz=F�<WW�t��I��&�f����t,�z6b4�JgVj%���9ZA���]a����K6;<JfUb��yB�{����TyǓS2   ��\�����E&���b0Wљh�2�`Y��Ox �"&�j�z��4��<��J�f�.߸ʅ�B0�ae�@�)�M�%5�u� 0��i�u��ܫ�ǋVܜ���W�]o<��y)�t��"`��3���|�O�V��<�в��?�7|�}�}=��
�5������c�͞$����߹7���ڻ��;� H��d��,Zg�h�',9bb�~����?��0O�˄c<�41�%Y�dɖDY�(n�
"@�h4z���5�rϼ���}�{Ͻ��4 ����,tee�]���~��c0�d���e�8��ݬ���(���4�i!N��\N�VK�ણ����N=�����-����?�w_{��_�VGX�	�QH-�X�E[LwD�unagO�ŏ�ȏ�13��V_y�El��؍ڨ�q��y��3��"-��R��xУ?�j�7�^&���7>j���[8s�!���o��kaYŖv��Q�n��Ɛy�0Q.<\,G������bqa�҂�@V��P0�=�d�j�H
�:�DB+D�=�G�v���M�CXB�C,�P��S3U����@W�Y�q�4���^����A;-���M?�f����}j��sXc�A��!�)��nY��KO���`�[8:$H�k�/o�3��Y��8�y
4��\T�)
o���=���p�ܽ�7����[��w�����z??�{}��Nl{���{���=�˞���1�ÕK���}�K)Ú ���ǥ�;�"S~����8�j�\zt�ݿ�K�ԉ5����{=����zU�~4�%�����[!.�����z�X��js�"�O�y��&��p��9l�Y%6��v��!w(h�����V�cuٵ��8�X��;7P%p�	��1~��0*�G�M�8�ēB��@M�OFbJ@��'>����g��lݻ�*h�ƣP�`yiVz���������#M������dL�]i� �ΠE��;�K%Y��KD�C-��y��S}�Ϟc�Nk��aتV�~��8����"�hf�5Hm�:� �
\g���f�w�x/��^YzL5{�s�Qy��q���@�E�<��:[ NM	%f֔��Bn�z ��m�j+��i�\��HcU+���	�k�$�KP�P
�����v���yT�[¥*�}�|����޽5��l��[$p"z��4j������l��<� �T�����]8����AoЗ���m���-����plڦ�pa�P/����K��S.9a��>��!�`��_��_C+h����͸��`s���/,��Ňp��qܻu]����p,A�^itty��]�,@rdiy��o��vW���KI�j�bR���'���5q�L3T��H�l��A��L#y�2�Eg���j�IWdJ�w�턁-pĶ?�`��(�{湼�E����'�ֽ����pz]d����uҴ�y�D��~�́	��_l���;��y��A�����vW��]�&��v���UV�p-�E������}����f�]i�pܬ�\���l�"����Ε���:G*��krw�S'��'ǭ��I�J=X6�3i@�g���<~B�p\�F���	I&��;��HLw����F����
;�t{Cb���YIa�յ�8s�<�|�@��*�"m:b��d��͋�cn�����nK}�~<�.�#'"|��_��W���A�]Ā�i�3Do�-c#��-�L�dk吲2� �S�������>Bb⻃	������T�(Lr�	?HU���T�N�qeůo;��1q?{-��j�}nɚ�b&��Ї��`��˷1���׼�ebУ�M�CM�bf�L0^����� q�d���� GW®=���i,u/�}/��vν��u(qZ@�{�gr����\��:v����0�6����4�6�jkS��I�ok�e�ю�HFR`�	��0��!�Z��TKbP�7f%h�{��:=R�g$��w��d�q�_�{��=8���D�͍�z���L`j�r&�א(�f���K�5��\��K���v[My��=��W��f�Nk:��f�҈��@yw:Uģ]{,�⹆��/|�@���ł��n�R������˘#�\o,a�����[{�:�3�
1p%U��!��؀.�|�ӟf�66�i�f�nBYѽ�QIo��&��B���M�{@�;de�L���'�C�`���0B��1pu������o~����G
$�a��9�\j�_ &���86}��ݠL\{r�\�G�&A�u�u?a���[��0O�Q���5��u�`�ԍ�I�0Q>8��ҿ�;���z�Iͽv��^����2��d#b����o�"϶$"���h��+V�c�&�,��K���|gN���Vnv���~׮]O��*��Z-�����~�����x���Zմ�e#0�E�K`��＀O>�0�}S���X�9*~�)�$O�mm#��"ླ�������5Є��mw��?����JGN���_¨���	�Ll"G�Q�W��2���Fo��K�_IHmd���ir���#+��޺u��=���67F(f��%������;P`f��s8��=������;E�km��?�;|p:���6�Z�2$�K����Z6&���gƂ?�k�y��N��ߴ����c^p*���a��y�;��%Ȝ�`�g����0Ӝm���N����H@vd%����8�lC�����vY&l�K�1�:����k�n�#O�e�B)��C�ڤV������t:�N�Ql�ip���+hw�x�����KQ�c;q��Z��,�.Hv';���cL����Ġ�8J9ꍍG0M��8��X��-b��'pk�Tz�  �T���m	�
U�^]śo��"I�������w�:J�K��&$f��Q�8���`yn��mb�E��8�}�I��
��ئ��s�$��C��~���/eb�=ODS�"�8-wjоW����9��I���9ό�_Q<�A��u�1©�ymq�"�Mep¯�eKW��<�p-�����$�sO���>��暽�d��<�9�4֛���4�{�3NX��6�|��^כL�=Ȝ��	Ȏ��1�K�y*�j���Jn����jS?���)���ҭ����7%�T�8~���N���bl33%i����|���Jj)3ԅ�EI]�>���۫�r�V�����T�Ҵ���\+$6�����&��_|g��.��J��J�,E�Ŏ:hcs��[w�DL�;0B�Zp�7K�n�@���c���ξk�v�:N�XB���r� ,}k���u/6�@
�̠�zX��lo��iJ�l��4��`f���՗��;��*ǹ|����"nO����b�����2uRE ����;P�N���"�����"��r=��8��J֋�<�/�f'��Tzf�l��-�LR��1Q|Y��p�`!���޻�S����5k9JMb�����Q�ulkz��R�5��]IK��k2����-�8��ԡ�0�$H��}S9sg�v����S/����F�;�e��ܘ�������0�����?�3'N�k��LZ�Zڤ��\�	 yF~>�iH��صL2�F�5��b3��D��I)A)S�{��.9[M��2V��se�����l`�9�V:��dc�]k=ۘ2S��ۼv�t�a�oݸ���:��:.�:/�¶Y��Y`�$��Yߐ8V.XSo�a�@����kW�&5^�7����g�38s� l��S��Q��gp��[�m���1G�e�Gz4�;��YV|��v+gN^l���6m�M33U�{},-,�y�}�ln��~!k��%�3��R_V�6����1P���t�Cx���[�}'.�G�Gk��G]"f�uDÑ�T�9�!d3����B��Z ��m�.m�wӅ1øΨ��h
����4��lbS��V��$�������*D����hJ.��n�r�7&��T�i��,��ٙcC�x��J)H)G<b�7$�L���}�s��ͽj˶����K���X���r�@ϲJ�އ�Ĝ��ON��7�:��鹂|MǪ��w�(5M���l���؋��;S��t�U`�+�jV^����}7{�d����p7Ӓ���Љ=�'���:Y�..�H˞���D"M�?�\6Ag<����zA��[�g��>��3x��ǰK r��5ܹuK[�q,���f[o��kwn���]�#v� ��[o�����{���cO����P+��`�	|k�w���H���~�.��hh:_j��8�!"�g��+��·����
�{luZ�qw�V;��:>�c��?�����e|�����fՙ
�g�w��{��	��g�i+��jz�G6��c�v�h�h��I��r���d��J� �X�? {�i�d���X��[�4�w|��.E��c�Ԩ�{=H����4��Wo��B>"L=�|����r8���֩캆�l�~&2$G��+�oώE��Tׂ:1���������.�,3��D`��l:���{��W3�Z�7�
#������y�j�q�|�2N�3���c��YSHR��^ǕH&r����Á����t�IF�+�h��jiz��2�_�'L����Z���K�귿�o|�kX9r��_�\��2�U+�Wp���Џ�x����5����% �J��Bب�n]�/�VØK����R.������Ս[��R�I%�TX�@�@��屈	X�aFCkT��?���g�ܝ�v�2._�nm�E�]�#g���Ï��~�G��#�c%�}��O}��gp��z&%���m�Xt�RA� y@����`����d����@���C~�?2����m/o�^��{œ�u�:RU�0G�|y��^rS 7��Ű�W���ʱ1m��M	�h2�A�� Y��/}`"s�m�����J��$j�kD������6}�̽��Q�	I���0U�>`�3I� {�9]:g�NHۊ�6}����yG8�ާ�p{W�8��<V�����J5��)S����s����O����abnq�p&�A�������r�?"|�0_�b������z�*��^#�+J$��e��֫������y�kmB�KI�����W^�:>������V�V.U�̓�Ux�KA�i�*�����Cס<�s}{�Z���ʤ(�,��*�O\>���]V�K�7,�ĉ>��ɍ����Uh�:bӍ��^���#8q�,F�!ڻ�v����띝�mn�~k�ACҍ�&Y�k���-��=���H� \���?��@�U=w��Rsd��eC�{/���O�R�|{:_����35|��y��$� H7��	�h>�Ý����K#\|�g�qء��T�t#���O�a��81K��q�����x�]n����=��̵��S���˛rP���>h�A�UR@L/��e�3'!�2�f�h���V�<�-𳧐�ַ�6��e|��3B�M�o��fb$�.a��JÔ��"%C��>1��6�,���wu���|�RT0C�{��%�oL��%`���x�qw�����f������'�4P-W�������CDL��F�!�N�kršS�/]a��o;��.����H���^'�]�;"捷߽���'���2f�c�ry�*v-6mp�ma���d}i�%�|��������u���@��v����V���}��?g�Iў I�ܦ�?���df�t$D���IL}�!	������N��M��h���M���tf�Bk�v�ScX���݃fϟ���@�gZ�z�';p��.샰2��ԉ��&(� 0��xM/:_3�L��D��:A�.\e�Z���j'n^/xEOXc��p��~&U�����͚svn�ܱ[�3[-3��Z>�Zg��7d��ߝ��uΘ��33�h�RC� :��n^1e���)b� �>ivS;��>x�G��X�i*����i��{���w� :VP���`2R��0��R��tD��;��\�j$̲�� n�۸�y�n��^%#�cV�q��Ƹ�Fj�s�%�"a�zfQ�mvИ;��l�Ւ�Z�I�4A�\��u�ƌ|fH?,4X��J1���:M�9=؀R���ô:\���qQ[&u�>e�ǟۃ���s������%�Oa�ʂ	;P��g��n���v�f6�CC��G� ���<�c(�Uzd��g�H���i��9a��)�����3Q�2���;w;�Y[h��+������`2��c�1[����#�JX�4��e�"�?y�H���.�{A�*�S��&���\��$<�4���~TM"�T��]�u�~[);��O�B�������G���\��4��k+��{�}�>̒u6��	�=�{\���lgr����Ц�T���lE}��K��v�G�`��40�h�_A��2���Ka_�.*>O�l��}b��=�6sBZ#���@�F]Wv�rmW�Ru� ��ۜ�f$U��j���B�T,c�A�CI�0���#&�T�M�G�>����;��Ip�'Kpj/ziJɥ�Y ��]��Ȧ���������c��~%#�Y5Xݡ��Q��c�a��,����t���ӏ�M6a\^��3��y]N�J�]%07Sj(��r��v'3������ň`Z��*w!��V��N��k����k�|��6N�w�#cT��p0J��L��ސ��3J�z������Oi�M�L��8�Ĺ�tJ�i � �.b�:���R%���Λ�}	C�f��|Ʊ��.��1�:��FCTS��A�65���gB�7P�N�	'ўH��07gϩ�D��e.��@O)[�T�;�x"~2�v9H?��[����c��,K$u;�����P��؛0$-��z�L,�����kC�X$�ؘBi!c�m�X�l4�J�Z(*�)�-�E�Y�ci#3�����EI��J� �,���������hB�v��7���ޓ�lɛ�̂�)Rn���{�*2��8�n��
�h.�'9M�5;58c����T5��0Ec�%�d��\Y�'i����yml�FH�}�5:���{_M�EylV;��pXa��¡�b�� ���~x�s�7W-?�,��̺'$�%��_���y�X,H��V@��j~f���=7�v,�'��9y��i�s�1XhJIS�G����>�9�v	;Nv�]؁M>HiS�G"�X���[*Q�$����&�(�:�u�-�Y�p{����G����l`kȳ���I���'FvR��)�2"�� �]���QP���T�d�i-A����e�H9��􉭽���u
����1$ߟC���V��T��
� g<�6k��k��N�7\��������f�T�?�C~��I����#�g*6!#����:�6 Q�L̥��61��8H��)ㅳ݄����Y�ɆuZ��*�_z`�,��e	��jB��v�z�.�yʺl�����e"o�i�2v�D�S&u6p�ܲ�D6�o| ��l:#<�� �H�8Ʊ��2,;G"T�KR(�GH��]YR�iՠ^-����K����e��M=���"|���@�����mP��  �}=���Σ��a��2Y͘H<U>�O�^bQ3�
S�i� ;�zփX�#�A��YŌIA*�[ 	2���ā�����& �3L9�f��#�M��z��E����33dy$�?Y��JPV�o:�&��n$=���ɘ0��6k�ܱ��+������{J ��pCk�P{�8�K��̚��
2�/��g��T0���]܁�$���N>������AbY��%�%m욑��)Vm��U��-� ;̆�L�.�K�Q�3�����P��
.�=�_tz,��tb��P����eU&;|��;9�E��	!�1�$�G�͡����(�ls3uW�s�4
l�<�sx'�^z��?26����N'����0��d�mz�ӶR�@�ӡ�}+��>#��#m�U�ρ(7;���ə�7(qrK�$袘m�%qk{N�bo��OjL��̡ĸ84hh�-J���-� J�;p#��6IҵD��8�X'-' 1���{RKa�6'�)d���wH�g[k�V�sv�Tg�k($!j�'*�5���\�[�ό��fI�����r��:4b�l� )��ו���f���''�9���T! g�-͚��2�X���6}UM�1���w2x�L��X�C'��I�Yٱ��ٜ�,1.��l��Y��D�����b��<$Fק��)��,��P�}�6���%aY���`4���n�1�(�42�B�yg�!1ff�c���ش�_Sn�`T#�,c�p����T�l�]�)�6>�A�7;׶e`��v^�|?�S����S��F��7�3{�9��#����ޥs�]Y۬�t���x��t�%�J�``�5��Yc"�ӊp/p�������no�{��N" ��~Ѣ2G��z�m���8��za4���k�U�lz�D)�����5ܨ�R��D�{��������t�(nI?�!�W.��qΚv?��	{Lٛ�$b��U��	v2���>;��Kt�H�:�.~���Vh�H�=��	L�xw7cBc1�r��	Q�e�9I��8Œ�H@�nl� B�TEXu�[��ᆕd~ܢ� �]�|�*ѿU��u[�_<������zX\�����J�>;�A�27mU\e��CP�H�o����bd�A���I��b��('��D;@������DU	]�3�k�1��l�B��r�J\��EX4��ɲ���͝&��
Ft���ܜ�I���%F��ܡ�����+��0���~�B���J�ϳX7���n^�<�ōc8�l2���ʂ��W'�$`1�	H9����Il�\k�1[E}�a�ǂ�,� H"q�ܢQ�g�u�hߕ.t��C�V�#�>���"]�!`J��h~qQ�|f`N8 /$�L��(8I`SH�I<�ӫ�f��u���69K@~��TI�.�*(Wj�r?5�"l�]���$n	~�l�Gb�:}�^�	�K�2=��L�67Kc^��ءl�`fMY�isq���&�|l��� �r����h�ے��1Z�&�Hcɟa�� n�:0���}&K7͛>�#�>�Ū���.nyˤ� ʃ)Sf02��$s��Nd;������eb�=RCXrpAl�b�96��b)�drhWU�jw���eS֎[�p�+n�2�"\�PՄ3��NG�8��6�����	 ��Ł0aV�yk� 7,ܴ%�C3��Sm�h�߰e�28���앙��U$R�f��cɔC���̚Z8�vnqA¼����K�䰷R�"�cҭV�K=��PƑ�?~�}~�9��h�\ښ��s��@����n|A/g���Q��c��͚��&P�#�E8EY�@�z�ֆ�c�jX�;�����ڛ���Gщ+R�Hb��ev޼^Lk�������O���\�T����w�}�N[���?��'N�,Ӻ/��n��*vL勣�Уq�/�~�^�Mc�f����?�[�o���ui���C�T��1�$�I����P�E��N�����`9V&�ҰF-����y����L+Uc'�-��VGI
�d��D�����D�DY(��(_����{�{�78�gq��Qq�qߵ���������O�v�(��dcx�5������=o�qo��`������ҨpL,�������G�,0f�:6%�8�Iۨ�-�"ag��!ui�~g���,�~�)�9v��`Y&a�1�c++t�L����w�E��p����z��w8
hJ,*���}�84��Swآ�0GbF�Κ��~4B�E�J*_1��}*7��.����:��1�W�X9��8��Ʀl�/�KtO,y�[��f*hw{R(g�PFcaI�g7�ML�x �5�j�{���W%l��l��*�����ɌM�D�XU�ƈ�S�֔l|e�\�\�����rl�����vWu�Gڥ�������_}���&���Q��k��	h�(QE��f|�J؍��[ 6��I l�0!�߹��v�/%Ay�3��j{!�i�+�I:H��S�bi�Xsb��l�!f�v�f�������<�/�ta��SV��g�[ ,��o���=}��w��;@�<u��1[�;�|{3�3���ԓ
&0Z�P0�_�W�}���G�Z*��ɤ���I��=�����O���¶1N�f��#Lx�k�G��ADlH�N�,wX�+�`�zI��`̠S�H��0n<��Ȇ!{�iqq�,m���G�����,������-z.�����^��/~M��l��S�O�FR���%�5��Ib޽;;;�U���G	���� B��K�"�M7xveG�fIr���X©
X^9�}�c(U�h0��`c��븷~?��&޼��8���ñ2�Xa�b�,�A�AQԿQl�[�G�R��T�`e���|����EZ�s(�����Ǹ~��\9��#�eai����E�k^кrv� ���~'�P���'�-���υ�p���ȕ21�-���;ľv����Z��f�̊k��E^v�Q߳E���I��`"L��2������Zf-ji�(}�1�ol�6T5a\�� 0�b��4$@i�����X͈�=�V�������2�z�!54x2d��6��E���7�	�k(�����j�(�/ym��KG�1!BE�a���N<���:���e6���ve/s_S�(MiI��죉,��9s���_�D���������o���5�iGj.�`�'�:���L��T�y��.��8���k4Xunj�7Cj<�BTh����������Qq�V��V��!1��2mc��4�$m�\�"���q�;�������������6��]�c�6�mH�|H ���,5
4�rm2[��+	��mTf��}1�l�ԗ�ԣ*�R+qa�-�lP���hg7�|gz��c��tn-1��8���%�>~'��;W����mE��l>9��D���4_n����b&��̘~>��sX&��	s�t���A��^ 8�[St��w]*�_c�w5��	���%.�䇞�r����N�o��I��G�]��u`�<�i&Uvh 1�W��K�uGjl4U�(�+E�
U�p�� TF�&�u�>��X�*g7�MW�	�Vs�>�,������v�s���We��	���&�7m}��,�6�8�3��Mo��=9��e	�z��;��sRs�5� 4X:���ېz^��֊dEn@k��s�R�tä́�+�np)gM�چ���7Y�niJ#e����D �#���I�o5[�`j
��Զ.c$�X�^T"H̿)������dck�4�E�>�Ui���JG�h�l*m�څ9�I��J�QD�B��W�~@U���	<���j�����[I*j� Re�F���&u{���W%`����ܙ�E���W����  ,�2vh1�$p���'6\�j,�jh߉�=8?P���`�>K�^E@�mR��U��;$��;�Q�;M���0�?%l�*�ă{k��G�է��2�$,*�ޅs�퐊?��_�ah5񱏟<M���?6͝�a�4�=z�#t�MR׶i�q+�=����w��#�ry�B�
�P$�!�
��"tN���c���ͣr�q�Dh�;	���Ga�a�z\��F�xø�aVI�S�y��\<v
}�Y�e�YE�ָl����]�M������ZmL�gB��l@ϰ��.��R-�ُ>G��t;����8{��.�>ͣ�D���nF�ڌ���Y{�_�E��xe���Gܐz��'~XNgj��ԥR�w%Ӊ����v�%3�6V�;?����?�㲗%�"'�pQ|�z�b� �^#��d�5D��<Ǥ��]i�4����'?)$��[w�r�|�٘U0�<&$3N��4�P��I0�L�:�Yz�/�;[8}�Ν;#$����b���w�t�0��1� Ό�m+<R#F�⍐-zq�� �䄜b*����@a�Mp�Hx{R�-D��b�������L�9���^�X�#��g?�xu��?�����*a��������ig+�]�{8{����g���	0����)�V�F�b������H��]�>:)Z��|���9�rl�0{C���Le���"f��V'�,�h!
cy^v�4���+W��ׯߤ�h���ai����&��Oט�%���m]^A�����q��(X�Ug�&{d��E�����X���w���2ۨ$J#-��/r7Ǣ"�����%�c?Tޚv���ǡ�{��t��r-E\k�83`0T���UeO7	�B��۟��ۍ���1�^j�I%�S�����8�1�I9�72d�̤}���ݕ^lO>����j��KWX�u����{�\H�{�@%�`eclS���x���3c�i����j7�ٵ�N�ج����Lov�D,y��b�tZ{5���:<H�o~p��%�l<?�J+��-=��X�>p�q�6�*�=2'r5����Id(f�X�q���1u�3~6��/� ��O�rX�{�ocS�M�>k�W6=�H�h%l�售�pm�M'N㙕�-R{%��k����1�����f��W��&v�M�A�x�����F�M���d!1	5ꓴ �s�;�8I v���A�s�����T�厷[(ժ�7j���Ю"����>t�T�Բ 5h<�khn��2#��aI��V�q���z��M�\{�-�-����s�m�;���Q�޺���e�޸&�q
��y��{o�6�j�� 334�Us|$�I�tF�.s�'��'��_���}Er��Hm��%�m��/�O%�f?{ӾgH���fS�ς�J�e��)��)�,��4��Μ��?.Q��aـ��0�p�#�t����e>χK���i$�y�$�=(M~X��ӳ����:!�^狄��0�:1#���E[�����߃o��u����>��v�B9�Ps�2�yTI�0�����RQ0B�����We��L2�3P�&�E3�uV��H�M&�8EH�GZR�\�]�'�@��9����|��q��iZ�!Ο?�nk�n����h�nI�lU�Y`�"��1׵w^��9��
�rB�B�����@,��FwH���m<|�y������`Q8�z�(vb�hP)�Kdg���%=�ҿ��IZ=4��޸G�]��g�c|�&�� ��n�
��7o�m�k�x;-DW��K��RS�x����۷XϜ9Cx�@�$�A��Ǐ��v����E)��6��Q�9���| ǔJ��nS'Ǔ���QƶѢ�11�0Eqһ��ʅ~4>�zC��l�c�3Q�����9�}z��e9��
� �1�ڹ��](S���*�3��ݵ���'���U�N�܁��j�^t�7W�1a�S��c��X+�Ik��s9k
�p��B>��h��}�Z"�}_j1�
<�U���s _Oj.�6�E!a�H�]ʌ���yn�����ݥ���AXL�Bc�إG���G���ǉ�JI,?vo|_a��=lm����A� �H�u<�0�����c�{�ⱋ�qfq^l�Eb��b(�2(�.l�>u��9��ں|�R.�E�Y4�w��8r�T�R���=�b�x\����nWjzr������W��s�Tè ���^�G1.?�
��ܐ���c�u�WoJk��V��m�����ĉ����0�jK؅��=w^q�"\�x	'N��
}�k�\_[�N4��Բ@< t�K��p�N���7'$B�ٹh�߫d$߻���5㩰��@��,I{Jl�ܞ�����F��Ν:�����	��A��Lg~2ϢҸ��cc�t�Y���)�N�LG�>��3h��N���|�{��W%��g�q��"X�"��{9� ������݌c}�s�M^sHkh�����8mb�	�H���"�t�} �l�Jn�;��[Ӭ�&�Y��c�ֳϊE�B:���q��iR��87����J�!��}�	ܼ`q�fgP"���}�}���>��"u{Ub���NK�pp�żk����c�HG�zOYD����Hp3��6��[w��HLV-��J� ���@�Y����I=�J��R���$�R�5����	-["�Hb��ۥE��KĔ�J�J�G��^��߮r3Z��޿���?�.� z������u��r��1Q{���^��p��	�-��u� l�M�����L�0x�����W��Brk����A���N�d2{�*q~������+o��ի��%��?��H/b��v�5���S�󄚚e�����Y��+�7�}�a#��:l����{f�ib�c�]Oe����s{�Nf�dy��r�C���g�
͉�����Ҥ�܉`w�;��9�����	�>��� �d�	�J�:{&od/�����ӤTh�y�9�]�B� i��%��W��O�ħ>�W_�:�t����u�-��
=R��77�j�b��+R�#�0�;���-�{X�,����N_�����m|�ɏ@�Ć�]�:W���6����,�>����=Ie�x�F��>*��o����{���eVp���//����P�@�WA��<J��~���RIh@l���6f�W�|��OH�Dww;�[��E1X��8~\�/\��ޠ-a%l�̵��_µ{w�v�V�Ob�Mʔ�p(��F66p�sd<��[�߳������I�������l[zn��C��Z<£���)�<�l2jq��Ml`���gt��mb\S�^6�y�|M�i��_w��5�v���Ю����,�����)'�S���C�Y�l���N��C��'ә�!�$+`��9��ľ��P�����.B�?k��+�a�n��CJ�fw���%T��I	<!���������W��w_y	_8��*��>"n�Bl�Û$�&(������@˳��������[�����&v�F8�r� ��X�E��+��k����x�{/�3/=Q����(��3���������mT
�LG��W�_����/<B�ZD�0���6�� �t��]n�S�P�1�eu����;x�w�g�yrN��I^>��}�)���ˤ�����[�s�x}�A@aey��X��4��07=2����^����i ��i�O=	��'
}��́�a���T�7�jW��"�%�n8�%%Ҕ�4-T���1������$��e��ڟPa]��{9���>��Dk�� ����K�d���,����H_��5&�Rd'�K����SS�$L�����ƹ4����{-����x_��g/qj�3!�1���e�f��PX�n�?lS�Cl�G?�)�T��ZR���C�+�~�o�b���7_Ǘ���$1H��X�$R�;�}�N���bv�@��ޘ��Sg_}�RH�q|aNj%���9s׮��w߹��v�@p�G+B�����:��{��oa�^o��6fkc��r�Kȥ�x��4����N<"��!����{Xo���cO�g?J�t������{bt�&��j�=���#�Rk�94	Ŀ��oK$�믽J!�����*���׿v�]ܻw�q,1�hk'���Jxgc2�ȷ����gʿ�6�^��,\��v����J�U��}ʄe�[�T[ݍ��tz=�96�M1�>��Fe�Ůؼv#aÞl��9�L'7��kN%�?��SEM���	{>�4*�ӓ�'����{O���)	Ϗ=W���H�q��W�>�����cz#ni��Ï0p�G��ZsBVΠ�څ�%��1��Q��d ��{��{�����ҷ!-�o�]���Vc�U�!���rr]�~����B�e}*�ِ�6k*�f@���'�@��8+�>ũ�=b���۷�V�CIW�x�bXg'����3���k�������5R�hE�-n>�s�ԣO�P�'�"��<�;����?�+7oKH֘���9��
�V��{���?�u:�6�-�HJ��6��{�m�tv[��7����VV�ӿ�y��R���i��Ѽ��Ja^ɘ���W���}A��K��Ϯ���Sx���������	4���2��#��P	0��y�~�[ߖ�s��f0Ŝ��7�n,I�@:�����rg�Q*�B��Dn����ð�i�̑k�k��7/�9X*[�%��Jϡ{�<)k)�Ӽ����!'�	`9����Ye�|63p}� Q�CP�z�� ����)�Z�ʭyq�I‒��ia.F��J�yW�"��T���f�U�kH��O��Z
�k�0����R�?N�͛��<��a�='�Ó�1ړ��0�3�0c�^#3'�Mn��5��6�i\�r��׀r$��,L�qe[�H�t�� �\sGsf����m�2�V�g֦L�z׀q� r^g{�N&�T2J�f��;�雭�pk�&6Z�X�+��:�U�^��k��y�R�J��M�#����dqsEE�g���r�\r�6[@�y��A� o�>}c�
�m����Lc��M�n���1ʤ��CU"�8C�/�����5n��(TQ$V�v�:��<�M��=5p��슘S�<�7.�C?oc@ל-W%��B�?����_�:	�Y|��i��·����Z}�kb�-��O��[��ݖ��El����W�B���F=�>'��e����t.,[	��	�_YV�O�:�F�rL���Y+F��S�6LT�N�c3R|*�J1`Ig��e�S�cW�[�B��|Ω�	[�6�DԆ�YX�y���fT�e,�j�|>Ύ6���G����)Kȶjv����圳�f�qCΑ�t��H1����k�����|v`����=�S�	��R��n��f���Yͅ�&�H�u��R�L�	Q2h��6�Ö��[�){vd����8I�ލ�"�]�Cʹz<�OgH�/���m����!~�g~���I���۷����۷8�_2��@
�/M�0��v	dzR��o��f�p��Eܹ{C�]?�5�>}�Q�KL0��v�����Lbǝf��*-�<��=A+�1��1�Ao�asb�b�'Ϟ��b���>SS䅟�K�������&�\��"�a��X-�-��m7w�g�C������!���O��{��ڍ[���&�L�G��?�}�*�F���q-= �%�omW���[�ӭ��$����T���9he�|�Y��]Ԏ}d��Ԋ���AV�ݴ4}$}��e҇ �8�jd����u7�Y��+�Y������4 ��Si������}��I�P.�i�yf�8m������s�R���Ep��-1�$�0y�n&�9��y�Ml���?�g��;�'��<Ⱥ.[�཰s��a�K�ɦ7k�l֗�'�YQl�,� �vf��\n7���AZ[7��r��/���;��o�]<|���C����3xs�M�h���	��Ի(�E�ap��6^}�XZ\£?�h߸N V1loH-X�Ŗn�6��"�CKO�!��!��Y���Ԫ��v$ݖ����[�z32*�tդkV���P��V�@:� f�`l��8q�~�~�ZCڙ����"��N�^��������X�/}����`u1p#9���=߀X�@�{��� �[=4�~��"6�u3�E爹�ddM�b���� ^�
�.o��t�Q�r���Q��K�X9{��1���<�}3(IW& ��T�� ����6<[I{u���u=�l��^%P��au�ס|6���:�Ek�7)n�Ls��M�T?)"�A�e�Y��� 1`�`�M8�2�����p&C�u�թ)Oq ���N��w�	���Am�ۼ�m� �d������4�`��!y3�r��w��d͉M���&�+8i�(�#$��8cS�A���B�1���iM��!�z�$z����M���+��?��=�1�޼K�M���Q�+��2��)�O��M'��m�茇h�z������揝F��-�J�T(�_;���=�ޠ�A�*g�~��\нuIſ�C�w�sa..��V�Xw	Cb�u.,�7"\�b�4��²�|��}�0tO=�è/��Z�\�G�?�
�1����[�&6].��o��o���+'q��1ܿ{�X�ڭ�؈�=�61��w�cqq���*V[�?���'&.�14��\'B0�jQF�4�fF"�����Z4-���ld/�0� ]����Yl��p��̤~�� K� �a¨���qZ[�w:I9?����zG��0!�)evsf6�?�y����
�l���ЕЛ&˜pL^�wE�:V-mZr'b���@�|zʵُ�Ȫ	U>�Il���[b�tjw��:�*��aM{>k��'�#7w�&N�,1�6%�U�?�-����*6��x�,L����j@���.Ȁ��\N�������c�n �	uTzW��K)5��j� ����~���R�͛x�� *���3���Fua�B�-�07��qk;��"����sP���k/�����q��Ib��;�֢ �$I�������=oCls:��<J�"1�Y�=jiۛ����3�⭷/���gp�����v��樋�f ��"5>,k"��~��n,�c�+��Ɛ"%��B�6��ϟ�
Z�U=����_G��£�L��6=#[a�t��o��f��B�HªG���{�6�l��;�zJ�U`�M3�����_m�5����w� �$vQ��4���H�Z�ĴƎ�%�w���`��fə���.�N*��G��
���Y���%�٨���5vQ4I��ʫ���8��X����M=G`s�M�jN@�P4��{�ZȼHl�F~���ʚ1|Pu&�"��E�xZ��s�ZI��H�6hq�~�R��#N�
;���D��e8���Hj�
�H]	m���-��#�Z�7�l��;ȘfR�y�	Df�dѮ��?6�@ңˁ|l6�	ja��z$�q�Tgڨs\���,����k��WM_�u��`�O��hH@q��ϐ�o�����F�4#e�z`T,6ݑ*ag��}��mz��bET������o^C�gz}��ub��(CRݻ(-T1Pcb֐��onl�
�����"�ҫK/�Ko�:V���WN��]@L�|~~s�x��[���נ�3آ{fv�l��[�q��=���쵀�sL��+��7���1V�oag�COG��3�p4}�ja,�
R�X���q>K�g#M��4lz�Y6&K�1�=�	�ulǲ���l�3��c��|�ɗ��Z��M��u��)�ykoU�:�����Y��Fx����u�Q��'��l����Rg���4�.���%�o^���̔�~~KۊX�M���T_�|����S��9 .P[�⏶�
��-tȇ�1��˝{����z����sk#?�Y&�W������ڔ��G:z�%���k��B�8��%��A�����^*P&�S٨��À��V�+ǎ�8-i؂���4؞W��S�����[+F�prnn�=$����FX����n�Å`��Ԙ�'F��ӿ}��.}�
	c*�����ZT,)˼�k@�.��oݾ���JN�áO;ƀ�3^`f��ڼ�4�j^�"�-�gH
��J��w��Zci���x0��lnKQNl��:�N��y�9�m���GO�j��˪>I� M�E�>`�L`j�r?"�'φ܆�!c��L�V�b-�m��:�Tn�E���(4\�g1�X;����{�4o��NA^+��y�1�(���b��; �$��֪0��rn�����1�E�1?X@u��`�����h� �'O�CدeUbW�?���e��lf��<�����
�1���۴�#�&�T�Ϊ�F��>W�����LL\�^�o"����ɹwG�LhʛC�e�H҄e,�}�׍!�~VP��N�g��t���p&����\������l��~l:cJy�6�IRn\�YR]
����;aRH���M)��R�E���
8fR]��yf�y)��7kq H���-:���m�o �5�!�����%k�+�Q�B���q�:��OcĶ�2o�P>v����À�ۂ��=b�7w����E��&�Ml$3����#b���	��
�F�
�F:r!�>W+��T[�k������.�2�4�Q�<����/��U�Ơ(堥:Y��\�@s�7M`=�����JdӪ9/߻tSQE�����v&��֎e��]n5�cq�8����!��m�Sp�?���K��|ʴLa�0����0�
mM�u({�)8tDd�XJ9���*k4_�\�>g T��F\�g��6�+�$#��i����l�-^�;R�z$��M'��[��q"���mk�iD�4܅�N�2,$������3we�)�1���eV������#{
������{��@j��-�I�8]7#m��ˇ?�~�-w�ʚ]�q:ϼF����=%M]-I��i���MUď�p)���y�0�i�~c!�(y�dץѴ;�ڟg�v�Eq��veu⅕�+��U�d��&�ܣɰK�c��Q'���A.�����y��{q��a
��x��{�3���H½��(s���lf���y`�k���vlU�H&2L slUZ�=֑��T͈`�5�e�p�-6b��4�(0ōy\w�ma��Z�8��u��O(o4r ��
�m|��[��;�MM��rM��������ݔؔ�v��|;�RV�N?s�p�Z�g�"=,�H�X�_�L9�!j��2�baua�<���=�2���bY/E%��fɻ��i��hf� �:��g�H�$�j�1���v�)ﻣ�LFyG�>x����G����S���o�����]�7'��=��Ӛ�:~����� p�Q���������ro���a�q���,K�c	1kT� ��26�/mp`Y��X�B�e]�����/l(G.}�ڙ�JڒD�1��#�*�蒑L�Dc8@�
�p�6�$��
)�_m�Xۓs	��ڐ���j���F����՗�_�l03k�V���Z�窅�d+������}"��樋�^ZIܺOsϢ�i�9�G㆔*0��L/-/�Kk�Z����ڱvf-�@sH�G�T�s. ]��Z�m�)���e[�^ �������hI��N�À䄗����wL3[����:������(ɚ��0H{�œ�²6U��0���#n9���h�J��I�0��\�`l�MVN�I�?�l��7PZ�k�?�|��_Ž�u��9&��&�!e���h�i�������EO��.%8�iE�̓�!���;m�]��\14��#o&���2{�Me�
{������I����8L1�h�!w���dU�gH�&�~�i$-H3Y-kr��Db(�]��E���X�����3x���t��/Am�&�Cu�
����������W6Wi�z �|�)����b`��_�5�(��f��[�����qt��S. �j�*��ٛ������W�g�ʔ�D�d�݆���e�hB�SP�����g�c����˃��l�A����A��׳��F�A�v>B���6f:��ĉK�d��30�-��	)�/�}��׷��L�s2e���]�����1�
)�q���~��:��Tq�;�\o�h wa5����
m�$t�hR�a��\��+vB+4,���
�&��́O���J\���c��\y_�zdlh�T�7��Le�U�z��\�^��C��$7z��/�E�G��A�ρ��5�q2M��4����i�qΫ���>�q��O�4Μ<��ƒ؝�1�_c'd,��вkâ+�Y�q6�F���Qe;}"x��@x��r�
Y0�p���(�;��� �s�����:�#67M���{O�1c8�����Ց�R��^�͏�^f��*-�a��z�JZ?:�5��s�9,S�7?���~ǃ���|ޑ+�蕵l�`�q�~ZRŤ`���6	��c`#k�[*Ϙ��h��0��7��D�l���}�܋T^ V{�l@���q��jA�RE"D\g��z���s�\�c�7�?K��Xk��7n��;�Ą c>P�Ȱe,���� ���ٲ��6s�f�����k��x`��M��*��X��1�l�QvFL�����Қ�|����\����b�"NA�XJ;�9X1���wUR\�7q���Cf���r��_�;?��}�3X\:B���S0�J\Dxp�3��Ġ�f�5,�.��,�8�<Q�RR`�s�8-�$�ɢ�ܟwn#�]�_�F0F���;X��:N�� �'܉"�H`mw���r��q�C�vz��v��z$B�R2uxͺn���5��$���T�#K��]@��s��z����V����^�m_͌�[k������@����&�C�4VV��Ê�Ry}J�\�.��-�0����&��Ms�w���5��e6-���*Z��<舗/�
I"�p;,r݁�n� �+V?��afŪ3Zb1�R�-ئi$�z�ia866��+2� ��|�3.���=�\S��2c!�M�T)�����4�es�q��u����V�����W�a$6�Hj�i�	�1z������q,�e���A�G�[��t;V_�O������1��`����	�f�IcPD�~�&X�
����:�M���L\fʎ�S�`���������̜@QV������_@�ۑ(�U^�x~��3L~6�A�櫗��o���`kؑ�^��N"�7tll�.n��Gfj8�x?�ٟ���J�_���m4�����}�O���R(j�<�E���	k��Ԉ�?������DfU��L��z��rbߦ�]J�2�kϬ+�7_�I؍&T�:"�:�z���q��.B�� }fw#��q
n��t����K�;����0����&ʕ�Z\���$�)bX�ɳ��˥�Y=�ޚ@@��>E�H@7��ؤ�}����6E���LD@�q���[����3p�?��r3�2m�2ר�M]6	0�fO=�TָMy���`��p ��b��.X����ȟ���:yY�1&!�̓Ϡ�X @7�g����-<����W�"���/�>��3b�Q{���h��Fm�1dbl%�m�c��D �D�yu���KL��ݩ�☴Re�*i��f������o^�g"����^]��D������G��
F�V�A���O��2fI&�<��-�H��OU�bne^ƕ��'�α����D:�l�W��f�]"s���LcǓ�;LhO�MG��ޝ�?�>���U��(xZ��,���ͷ�5��
����o�I�O{L�XsD�vZ���C�,���FS��<�<�E�)�Ur��_��֙㾢�)��KS@�8z�z�1�zQ l,�ɑ}�
�7��*8�Z8q�T(91��0/�\,�҄d]�k��#�H+��'ǹ�!�mq��qw�kW���}�1�X�
����v��"mD1*WضH�c�)��mj&��8��8�����{9MR���@���3�qŅ�N-.���S�3�ĄeLq�����|]�1x�fJ&n8�����'vO�]4�w�b@�zX�>g�$�&h#�������5�@�DU�����tz�K�/�3�����"قڵ{k����_�+o�DSB���㹷�'��0=�Q�y��4c�R�����F(+�� �`����ui����{0�=�3ˈӗ�b��yug_��wQ��#� ���8�S϶`4	^��	�aM��T�ӑ���\oC�N�;�!���o�zk��t �th�^0�"�F]YA�G(DJ
�IkQŲ�U\čk��B�b��b�'oL�\`��#�4If���UY�,�klc�Cn���lAV�%�)*ٻ����K�o�8+���M��h�W	^�m��"k��v5�!��c�J��Lg@J���	�;^#���z�v�I�Nd��컑,���G���D�"���2�'�hFr�����C��p��tr	M�nwOlf�dL�]�fm&��I��P0cN2�w|MJ)߻:yL���.0ذ1	�1{��[��2����E:7m���$�SJAI(��KGR�96p�Рr��@�0���я~��W�� �߽���^�
6ך(.4P�d�u�#Rs�v{u�X4�=�L��z���iиV37R�9l��n�����E�s�L��Q-�^&�4��ł���Ʋ��t���'W.����J_�t�ۿ�;���{�_��ڗ��Ee�:ys3�rs̀��=8�B��6ۥZ] a��AD̖��N���$�Ieg&	��ϓ�AUI��p��.�g(�W����������K�Fq�*��b��a�I������ji*Y�m.��m>U�����{�&�<]���d1&Ϧ���3C�������k/���'����
N�:�j�Fs�C���R-��*�"m�
��Y҄�=��6vZ��;�Ĝ��,$�����׾��;��3ܥ���IR7����Aي[f/+	j�M�Ƶk��/~?�C������ϰ`�)�D�DRr����gq��Yb��aʾ���^Own��=���$��MP��-���l�:"\�8�����{��4�P�<�2��o,�7
b��VI�*�3qX�b�Mr�>j�Zr�+�}��48[���ב�L��pF籅E�K3p�>����$��k�Ü�-���������k�:ϩ�<f��Dڸ�jsw�� ��^|�Ul�v1"uw�lQQjwWN[�3��|�ݷ��o�<~�>r�	%�����&�S"�h/򵀤��#Ʊ/�ǔ���ky=�^��m���Yǀ�d�`2��>U��dp-Wb\��+�a��bUbmXN�X-���{��� 4��k,�;��i���<w�$��-�y�
v�o���X���W��4��@f櫒峽�%9<Kc�����T)"U�H����������+�i���Yi�$��|��3���%,@���������ĩc������">����?�s��e-솔[T+5�����t�5)\��>-`	��7�
m����B�)q�;��:��t!���y���"m��}A4.�wg�*�
ة7�d�p��X��3P��-�I:�*2ʕ������'YB��5M+vi�X���W��Н����1���x�-�������,~�3�C��
�(��V��/���o��D����n��@%#*�HF�������e�86���-�?��_��_�*�i�rg�:�D�p�����sv �=���_��$MH�$%,�m��ę�z�	��] ����I4���|�;��?����2�eg��I�>W��(3�f��6��b��$�I'UR6��s�v�6�9G������^Qv�י�w�͹r@
U�D$�D�	�")�
�,�V�^���=�3~�սf��t��Y-ǖ(��H�")fA� �S!���Vݪ��9����s�(O�X�ֹ������=�"��,Az6�.'��M��G�Z�ց�{�ֆ6����`u���a�[]���*�!��/�c g� GId
#Yq'�fW��9�g��W�{�
�] ���H���sd�^���cCx�ދ]����Ɓd]�dh_��)��NF�Go��x�bu14:�+S7qw���_�u����8
�(�,j��I;���x�8��"DHb&�J�7
d�����h�@��,A��tP�9�R���j�o%s�p��ݹD��NX?	+�g�L��L����>��y�_���B��HX7�����[�6�Yi���C�͋k��|2JcRּ���%���b����%�_��o&t%��n����3*�ҡb_h�K�L������h A�������&Ӥ ��� 
g���
A��wN|E�՞�B֨
66{3���kF��#��^�����(���Z�|j&N���$lR��~&�f�����������{�E�>ǻ�^��ɚ���yi���:vQy�}��J�9g�Z`Y�gvœ�=|��	�<=��U��.M������P�ӎ�M2��zՙ�ub:��"m�&�\K���̀���,�gxI�3�Q2?���	���`i��^�d��_/���m��^IJ���	#�()fFs���[C.??��*ϡ?>���ԁ�T�Ke� ˤ(d�A�J`>�42��� 6�G'�e�զ����*U�A�y���{��&+�%�\U�ɦw�4ӵ�;8u��x�Y:�,�/^�(h��o����.;�.o�����H��{?SL)˥�#	�ɟ�d�-.m7E�4ٕD��D�^�Y�ʒ�#v˽ǡ�	�����x�=�w�3ᛐ�٬X�ξr@�GU��2M ���G7Yޥ`M
l�C��u�텃��O��j�a�aU�������M�0G@�2,HX�!lP��0���Y�]� .5'�G�����逵h��t6�m�ؓ#�x��WI���,��s����e��Adu�I+��4�ʑ����I"K�6�7�����dqɣ��!B��9��l�i!i���FB!aBt�ʆ�3���zd�p:����[���oѸ�������-��B���;_frBʹf:<n&���nq��!ev�B�~��{Q'�Z:Ȕ�q��)��$��H��H�����Ю�X�6elU�f���5$����鐄hN|0����!�*��,��^�X��%x��I�,H}���EߍX��:�gΙ�<W��XYrV	����GN�c6�/� ��$<���d$d�|���.�֎Ep��{1�&d',�����;�8��Km��e�"�0N��>e	�����u�SS?���+��Dr
�������"T�Q���K

��I&��|��"��Z8%��&��>F��]���3sI�kJ߬��{��^�254u��)���eV[�{t�P|^�Fr�6���s���ط}�#~+�}zzo��&��ϊ�Bފy����\����)Qzy���8�.B�\�I�(���H^�.eQ�:��i���{VY�,k墓qM$����=YH	�ʍ�����ywF�x�*�D�G����E���.0�*���L���f�r�>��5�\5��?�z_[�@yhp!NR'��&�9@B�W���>KH.�>��)�%g�����N"j�IK&]ɐVf�m6��,w���H��t�"�C���I�D�B�_�X���Q/!����5S%�Ca�$8Hȸ=���!A�T~dg�U�;�� ���[&��Ԅ��n4}��E*Hp||�����ic�Hy#C� Z��+n��5�eT�\Y����
�|_��t.�����>�x!E�G���C.�����
G��
��j��"��+{�d&0x�HP�&gy�ظ�˼����4d+BX���B�wl����b:��35�޼������r��_��w^R�s�ÂIA�����yI���_ޭ2?d,�����J��ne�5_)[©A��N�9�/���E-��lg�ZY��/�[��,6�
�	)t٦@^]O�O�}	���]6�-����,M`�R��.����'*�_� \�U��26��\��H�K�հ*qe��RŧTP��F�bל)�[.i/���ÎH���>���wF19=��hS%��)A�/_.)�Ê��}#����ҔՒ�WE������g�epdXP��F�s�v䬖mt���4����<Zc)���94��rު������HA�7��Q��I�GY|��L|g�t��͒d{8�BMe�c��ʛ�K�q�V$g3�cH�+"D�r���.@���I�TutT&&G���	�">����B�C�/����-��t�!i���\W�����qҺ�+�Ll�I�W7�X��/JW:*4��M����~>��T�ИmFP�b�]�����зd�ͭ8��;�2�Xb�!jw|�"����bs=�ҿ0�����c	Rs)$�xh��t�>�>�[rV���J��"���ڪ��Υ���rن��ޛ��-"	ZbA���G���+1��Pf��A{}3)���v5H�m�6AyU���R�iCm�����u5�:�nڳ��b||�9=�������5��*G
6�L�jc����t�i�fsid�� �}R��R]�p�(2���>3uь�J7*}�t��bݲt�^�zM��t��_QR>Ƶ�7��=���ݢ�% E��F�M\��Œ��Xѽ�P��ĒL���,2^��vY�5Y;���3�����˵5wu�욟U��F��K����t6���!������b_�<P���r�w�,�޾(��~*B��o�9��ꭰ���t�+�J�	�|2cxf��[[#%�vg9χ�;�腭PUMr(g��汶��|k^#E��n��\�0	;�0���e罉%=ش~�	IrbpI"~�[�B:=C�^F&�Fw�r�/Z,���O����K$DKd�g����#	LR�-��)<~ЄHHG%�m.>*��p����bA��H�l�uv!�@�h!�˼ݒ�葲L�Ǚ�������(�R���[�԰	VV�)�͉��K�� ��9,�l�ǫ?��(|�Y<���\�y�G'QJy�5���\W`zf�hM��4��h�o%���بX��m�Qm��J�8S@����3u�֮�0��9i:�Ǧv�L����>\�~;6l��7�Ҏ.��w��^�	��	={�-*v��8�5��1�W.vY��ψ���:8��B���.y-+�� ]>��u1D|��Q�4lz��B�Y8�Ǌ�<��cX�҆R�	z�� �fgp��	��P���γeA;��ghm�N[KN�����t�Uf����^1m%ũ���gR�;�n'aD֒핒^�|��sx��Wq��ϰ���o~��]@Y2��"K�L����B�))�����Ebt7�A��ҾKU~'
��Ѩ}]��N�'�љu{��@J��ŋ��J!8������,a�3q��Y�w({m)�g�������ֱ.,���%l��EQU�곥Q�x�V�La���v����؂��EQ�*hk��Cr@ԚM����deb���+7U�W��|߬�/��̠2�Z�V>]νdD��孆��&O(��u����ɆOL���u��4k/��"fI����%���V��޳���a�}��{��ܷ�#�XҳABZ�>=�raJr8=�.���%Q��o ���y�~W���U2'�P�.��E3q�Q������W�~�)�i]���E��2]�%���F=�Y���$�}a/�c^�rE�����"�Ќ$]��$���Ȩ��p��_y�P�LA��*%����֬Ý�a�y�#A�V�i��/uM�7�0զ)������AN�8��1�Y�ARV��r�~�ڲ��[M��]
/)��%
:��C�3W{e29��G�m���y-���{��k}���__��%"_V��rT��M�2Y�X�،��v:C����=vCS���5�t����7�����M��h��Y���F����+p��Զٓ[V&��P�0�U.�|Yaŕ�����,�y;�z`8e���:k,s:�U��VE��`��E��ƮZ��h׮Cks���K5��������W���`�5��D�QU�4O��e���'ȧ��B�a����Aׂ�JW ��o`�@P�}�VYe�X�i��~g\�x�v����%�б��8�����HA��ls~W���8�I7�>\�cB1�z��Q=��5��8$���,�����f���]���~�Z�CZl��'*�Q'Z�,����־���i������Z�Em]���AC�M����,(~���d|B�6�5� ��Α��=��b�W��-|�~���Sh�E0|��e�g��Ҧ�Ӛ&[,fe���%�i,��!4i��s?C���-���9r`��r�8W����^�'�������X����-F��/�k9��"�FΤ�(:�I`eCTR�Z	�����@F0�CSK3�߿�4�/�JB;*y��=wr|���d�����s����"\���������Jx����*v���.W"(��b���2ڵ���	a��x��Qt/_�/?xH��P�BG�al^s��K9��4�jLg����U.$�2c+X�����x��!G�v;(��]X{������Υ�x���o������~�{xp��8~�c�kF��W,_I�c38���R�F�ϙ�sq��*)?:3.ZW���WR����0�s���
�ڦ��`�4�Ơ\%��
6Aq���$f�\��}[v#@c�E��Q ���g�6/�IJ{uě�37��.�%êPl
�q��ΊW|��@��E�YX��-i�Ei�NL@��+�;F�_��Ew�2��8(+�˃����}��w�и��;��Ѧ���'���쨉j�ʽ�w�g�Sէ|��_��N�-�vͽ���U�^�{4ۚ��Tk ����sX��@�ݣ�1��9��rJ;u���cX�u��-W�u��FxC!0��Þ�'���	�f�M��s�,�SH�� a��zl�����q�)�U��a��]����!2���Ν"db�cҦxȼ(e$�Z�Z����ic딥K���A�6s)ӎ���eB1��t������5�pЌ#�%K�V��B��lr3�ū/b}�bĬn�=�;�N���^:B�"/F���6�G��lх��5u$%t^��E��.��	di-����!4�@�.*��9z��'�������Nݚ�*<��p	�˙�K� d�O?N\��9���/�˖f-c��D���'�:���1��4r>)tQs�d�&5�^� K�ϧ�,mb"!L���&_��A��C���Ճ�K�ҟ���]Tr���֘��#�'/���������@Z:�R5���5k|�:��ؕ�**�%�e����6+������\>�|�' �3�
��*��[Sq`���Ң��1��04������p� <���Pt�w���w�����ڿ�����$Jt��n�B~k
��Og
�~-��2�9��2�����tƂ�p�߮�;sV�R�+���Z��^E(/p{j���?�ɨ2*m�lL���4�UO�vF�<1Nca���4�5�si!���0���?�Hpqr���$Q�rs�'QGhCr}>��!�Z$S�Y�|�П�_��*s�d�<]��4t��k��E\?�)B~z��6+�O6[�
�/�M�TA�+�d�Ӂ���H�+|T��M,*� !'e��<:ڻ�7b.����!!ǉ�6�`�����2+&���h�w��WvJ���_��N��s�m��az�xw��)(v��
S�q)���	��W��B����fs�S��gT�A�RI��m��yG�U�mK��+|�$Hǲ�����'Ϟƞm`���d�Ɣ��ST��Ql,.��ˮ�Qf2s�2t�m1�$�b;(֨�����׺�>ј���O��kd4��Jn|)\��(���Х��!��c%)�c-�U]��]@,�M^黉��|���=%AR*��ǖ4j�U9�@MΪ���
+k�n�1�J���@�<ڝ�����'G�ӗ^�o?�mD8�Y�	��/ȕ��dz����v?e�:�V��y;�P�-�޸��H�Z%.�W��ކb$�qNON�O<��'>�����8����T^[��+�.޺���L�>Kw�Ђ_�j�"9��ݕ�	Z���(w���.�W�[�(TGJ��\�������K���	ޕ��5XGؕ�Q�0�е �cn�"����ML�ڍkh7���uܷq&G'�J���Gg�"L�c�����a?�� ����`���H)_(.��PZ�~F�\�\)�|>	�4x�+��4cIYv#��ѿ!T ����SM�N�+Ҡ�jɦːf�\��E�7��qZ٢��J$�ȗ9:1e� �����'p�� �z6��c�x|v�=����F�Py�.��al�a`dd�1�&�ͤ1N�X�KP��t��7V_�щq\�qU�M)�D��Z�"܃�����0*BK��ݪР`�
�<Y�?�O{ϡ��m�-�����°DQ���~hAQ���D9`HɩӮ�br5đF�._��U��@;�@R�f��~7�rh41�#�>E����]G�-aK�0�$�4W�ŧp��Y��13�o�����2_5s��<t�\���wC�*c�S%��}7��|o���P���+~��_`����-�#�J�A8	�*ٜ��l]� �+�p�N/rfQ,DqYh���mv-��]���B
P���\��C�3�ĩ��r�_��&��؉�3p��5t�,#�W�:2Jg���?� �#(�8�ِ�<�G�8��*��-�:.��a�h|>�Um��g�Ԗ��%���<kkL��3�w��J�W�Ĩ?��~���D�K��oêy��Y��˭�/[*�T�<��T�������BBq��K�T:�E�XJ�r3�}S��RZȔpY�h%���<���#��I�CX������i�<He�H�cI�"�>��U�*��dri	Z�h�3)B��<y�h��2�xb����#�õڒ�&|^���.=�8�
�]��X�N]'�ފ��v�?g�{�޹�^FT��I�Oaj:�4	�x|	B�h��H��1C��MH��k#�j�I��3���KD�PR���*h��M_+�l�WTb���\�e����2w��*�>g�16zW���⛤ �*V
�lEק�]���[!����-�èj|���#�̅��I+�ZD��չ,��ϰ� �U����??�ϯ]�}�֢�֕���իeL��@��+�q�P��1Z_�����rA�#��=����E4ST-�2�f&P���u9�i�����ڍ��[��w�	Է���g��U��W5�l?/=��ef�:�oH��	#�j��9?s�w�$�{�T�Z�sV�Χ���J!�0.�����N�oz�Ʊ#t'�شr��Ju^���?9AJ��I��|Y*4.���	W��E��ru�g�v�ڂ�ι��٪
-��ue��\��?זI�j%�� }�s�犐u
,�N�Mh���e%I���ҵŮ�I8G�L��r����F�������+�s ����E�'��ͦ��ŢRI����'���&�.���ϡ��--�$A>Vߊ��	���m��9A^R%�*!O��:0���T�������g�{Č?$H�ɴIs��ׅ͓���M�r�I_�hr�:D�>֯!tv�Dp�tw�Ĳek wu�
�*�4��������7%5�K�n|���/'����y���~L��º4��Ƶ�[H�`�Y��Ջq/$X+��YQ�V�AN.'7��#��c����" ����+��P����r�2Y�A�9L�aTMG��U爅��{�dk���è�]����m���L����4�C�t���HH��@�K���k��LqY%�c�T����W���Z�#��\
ʰ�֕EE�D�?���Ԙ���Tn�f�x鈫�5���`��YN^��S�Y��ρ/�.]l�%[�S���k�b|�y�k>�]i��x	]�L��KS�r����:�����i+��}��h�zB�Y:�S$&�3�<y��,ə� {N��N=�����B��e�5j�zj5�4��斮M'h����Ϙ����|��_�'�(��㵪�R��n�����q�*��>"i������v�����M̐������Ё�%M�ʵ+b~��o>�Bb��^�.��#�-x�.���װ}�NYlR�hj�B��U8{�n��!C�q��2z�l��$
z}����굫I�$�<L��k|rR[�����W��a�ǥŉ'H&i|Vj�M!i.��	c��-��C_%�'�Z�Tw1N�I��b��?2���5���`��͸x�<��	c6�A6τ��5�DO�x8�1#0�B�)Z���XPE��<��-� �C�c2[u�P,�dy͹t�$"�.�G�.C*�R�
n�C��+�q*��6T�����EXp�+��v�6���㯼��䲰��ݸ,[�NB�B/����xzZ^瘀|t�d��s�%)���M�^G��)�W,{>/�]6�~�/��2VM�!�p;p�f.�6h.\B���Ec��$}�tu���Լ\Ps`j1]u��ײ��������V�V{�\����TX���q�x���[�m��;I�*���
��� �Ɲ����i��:�EG�x����B��t._B��8z,�)��vo���wL���YT�g��6��Ҟ0{� W�3��[��rU*��!o��㻨H���΃�:�� ���p�L~�b���C�;��3c��̧hnh&�5J'�Z]Ӓ�ʄ8-�f!?�r~$R)B�%��*�0��qn,߰�H(|�Y&�G�v�0�LK]�H"�$���/��������d��+�4[�H�d�fQ�x̠vM|~��>�<rE
��sy)��hv,\�][w��~��I���HI [8�ȄS3S��_����}=��i�IQXҔ�.U&��0�޺us��S��g�1[H�&%S�+de�� �s�]s@j�T�Yi�j?9�O�	a{h.Q/�Y�Mh�������(Bሔ�NM���ށG:��7o���u[���fE�������9ޖ]U�&�s0U��1�R�5&vU�C���,��	01	LN�^�܎:H 1�!��s\!�T�MK�~�Z��:0���Aa�*i���RȌ����UcQWW[Oɚ��4�r��V��V?���Z�Q+'ړ ��p�,�@{�"�x]��+�_\~���&t{[;V,[����ݺ�D.��,�3+���L-`�.Y�W�����5߿?�c�"@��{�(��Gw,���BH�AH�j�ڔ˞��Cɯ\t���yŅ�d6-��5#H��iR(É9\�� &pl!�pzn��IN��ո;*ယ��X��q��rv�kv�r�Jи˜���^lq�n5��Il��E&6.��Ga�������O�#�js�+���c��*��[qh��O�'Y9��:_�:F���D�.)�{�f�	z�A�hs�$�d�ee	U����Ӹ��O���%�o3�1l����Y�s9$3���=�p��z��P^�W�oe���dnAoL�@����5lBH+� ��";;C�X!#@6���V*݋�;���U�q2k8X��Ё'��?�E���2��,��#e��%U	�"���q�iܷ�o"P���0�Ma23�$!��i�g�Ad"	�v�����-�])�����#� �wk(��Vn¾�{��{9��:��i\�y�.��dÅ�E�E���"><�}[�����A*��Z�S���1<=!��A׀ր9$��F�:��V��9���R�0�c��N,�3�i�}5�F1U���.Bck��ي�w?�����aln��?btrPރs�q��G煫�v�݌U�V!�c�*�:�>���a:�D���&]�%�M�IK8Hip�Mf�V����aT�}m��\҈��R�8㍓؅��i~M�zt/����k����hmmb��dݹՏ��6��R����c�}x��Ct��#��bo/�'G�;؇��I�C%��^E=�R��9]Q�f8ЧyT���Z2XGV� �-�ai�j	���Rf$Mg���h�{Za疭c�t�K׮���,H����A�H���Waώ��'�8{�3��$���_C��3�i�|��::q��cƮv���TlkAe;Ӱ���E�R�*���@���lu����qU�P�K��,x�����`W}�����j��H~�O�f�+&�ᘂv�TꇕZ�)��.L���E�5�fP��_,��Ğ 4�������Hg���a2a�*>�z��/�/4�ꄡKDHIUqz���y��>�D/~�~�>^8�V%�	��+�H�C(h�����p(�x~9]b�����9|r�"U'`Je���g'�	3'��ڹ-�ٹ	�Bs>i(��y\9;A�Fď9���dqz��"�W���u�AY.�6���D(%�Df;�1�C�Gi-��voٌ�t�7�݂h�Ax59���ʍK��L�c�b�F���&E7=9��/��K����O|��oŒE��}�f<���;8���p{b�0X�n���X�2Iʓ`�CRRE�W��ǚm���G��
���O�բ%8�� V/_���V45�	Eޝ�!���K�sn�CtT�
�PHpݾ����3<���ز��پ��n d>���*��ꝛtf-x�P�T�s��F0jlC��E;5h��R�qd6eUB��a�%Z���߇��?J��X3����o�w^��W	���}K�t5��~��qp�oَ������I�y����52�_��U\軆��&��t.�$����mW��SN</1�6GK6�-�\��&<��y`j�MkVce�JZ��t>��>0D������s<�0I�h�&&�'`�e�}�F�ixd��W�L�:̒�dw��
qR�Ȱ !1�3�Yqq{˥���b�\.J���+Ō�о�U$\�l�%h�J,J��t������>ٻ>j]��n��X!U�pC���UÈ�K:9�4ms��)���Ӄ،�!�'�,�,uD��V�����	B�c��"	15����$�;}���}U�
9k�L�*jd(�MB,S�,�J�BS��)�_�i�����S.ݮ��<!(�t��'�l.�H����� @;�d1;Gd���E+�\��~�g#!�p�굅��x\���� �X3�ݢ�;v����m�V	��qdh��>=����Lv���y�i��xٕS�q)��&d�ӟ?��t�w�E�����˱�c)�l�M��	��՗q'5���Y@rd��XeG�.�@U���RpjWm�mR\~�Y)胻�aߎh����D}:��ǟ�����ӣ�$Ę8,��l^f�9A��q���$ &�O}8�fB��,Ǯ�p��8���G���k�����KS���I�s���D��>�T�Ps��sX��۲�����e���FL�vl������{�Bbv����eD�AX���L�M����y�W�#�Cch6��5�%A����d��Ӝ�� E�J:�Ґ��;�D9��U��5.�ܔ��q����`+/Á�`��M�����Iq����w08���7�>��X�J�Vޓ#�x���ok/�i,]�Wl�#;��r;q����3c��16�>v��m�*�˛`�U�9�aT\�g�T1�*c�}��]�~����vWV,1K�"��������Ul�{mŋP#d�MQ�+S�1R��-�=H���*KA���e�L+qk[I�
��z�J��2�$) veA����+_H����gåM��ڴ�\��N$�\�vj:�QPR̭����� \H=��R���1�3kV�'G�]n�G+2�e�$�8�&y(�gqX��S��
���N�rH���2�i&�@���ֶ*��K��tac^7�v.�#�û"+""��S�B�G>9�7��%�K!2��bh���業:w��F��:�H:���9����ȥSx�����Y�܁�?�4֭؀�x��p��E2Uu_hN+beh�k�UPe�rZ��<�z؆1�k �s�5x��/c3��\�Ϸ�]�S�x����滯!�N!ԅbB�.�U(FJ�]QR�gI��Iٝ9�9�i<�����JB�G�o�S_zWm�+o��?;J��m���ՠ��W�Pu�j2��ξ��8�a"_B�Ʋe�|�k����؝�*i��	ͷ>x/��r���+%IQ�ْ��d�Y	�1q<+.��R���$~���=��o�ޠp��Z�?����	���?�-.ܼw,�D.���y�k(���OՔ[��*[�-N,�I	.k�ēǗ�����b�Y2$S�Wo���I�n&m2�r2���O�"���+z�Hg��~�*���7��t�w��Ģ�.|��.��/�q�|򡌓���^�X��]��;w�kmz��f5eK� �UsW��T��&��0��VhZ/���!�Z�¥[(8�FE�����	"t�4tZ5u��|_��6w��	ȅ+YE	@�t)�s3FSO@_��c-乆"͖�R�r��S����+��[gA�����h>�~z��_���q�˩�%d��q�uQ5����>���sk!���E�**�v-�<c_!�)r|C�ͬ���u�P�Zz*7�a���M@f�W��$(�����u��o}�ݤ \$XmN��r�E\�p
ׯ]@��@GS[�<����
!Ivn��9�7Q� 䡋1��\�|�LNN`ߞ�ty"d�r{��������~������Y;+�&,-[����8��NzN�>P�٦Ҳ�����xt�~|��W��P3�p��+7.���q��e�&�h|ZcA4�7!=���!�K���٭�mQ̑UAVF�?F�3�Df
���1F&��c)��X��@�;��?�C�ޱ�/����ۄ�~�*�`7�}Y�ٖ��t�e*fPVݖ��aBg��'��b"�M�-�7���[�č��:� �z�������gV�U8�%DY���L}�� �J�W~���<L�<�
��>l�Y����3����׎} �Iil(�T�����	3��str_Lfĳ&�Z����_y����F��@2o�y��{������x}��loSE64�t2��n����7bbjqB�EZ�_��<���S�Z�/͓o]������M;��/�r�5d�K��"ʥ����K��8-0�+�厕k�}rV�+���� ��>r�t=@Y�:��]�!9���IjX�^�Cޠ"���ui�:
Y�ɇ��.*������V&��}Vlnq;�W�T[m�UdAK�W�����**7&�`��bD�y�,`3��[�,Xw_��tj��34c���:Cf�9t�Gł0��"i���&�eeB��\Z^�R�iii�g�q����������ښX袱U�>��29��n��l"a���~_%3��rEBK�"�;ro��&&F��h���V_���FBF6R3)L'���\��t��9y�B��s��֚K|n��>:�	��M�F��7��5�V���<�[�*��/?��|RRØ��hݦ�İ�h�a.�R3�I��P������_#AF:[B�^w��˄^_#a:���:S3!���ې�ț(0M���Otf�HJ����vs�M�������u����C$�W�,g7vm�NB+���o�+n� M�����^�T\�����pY�rI/�c���|h�.����A]�Q
`f�Y���Gx�臘�#��C,`����u�g�M�Z�f�]	�JP��\��d��&s3d�����ŅWQG�y�f�o	�:��?���?~��	9r�6>�>�3G���+��w�����Q�>��C;&3�/ ]�G��p��g8~�fg����Ѐ !ҩ���U����9����!D{�C@�}���$��'?�ν�c���떯��.��՛��މ��q��g(xX���g���X�P��^M~�Ӷ�!|qX���۵�_˃
��QS�V,+Yڂ�/d�h����?�w[:XfW���Z�9@>
r����SiPAB�(2M&�$�)Mfk���R�!M�
,D%��!!юj�1�r�Ň�Q��7S�ɉ0* ����WTTGe*%����>�Tn"��%<" M�� *n�Wk � �y呦��"�6+([�C'~��]����s�	A&#���@�w~�x�����;g����^zG�B{�E4�����Gc8"-���D�����ˉ��ȇ�6s.� L�^�J~B�a�����dr_��_�wܿ�~<��t>=�{���'�_�d*!�Y�d����R����RQBL�H���;��������9���Wq��5�G� c5������'15KJ;�	K.L�:By�� �H<���/{�����ۣ#��1<<�K/���G���O���潒~��~���7�:r&	si�c+wͼ�	�.�ݑ/�����O|��2|��	a^�zϿ�<.�^""
/W:�� )�EM��[��h�8+�������DI���RP���%EB"HVG�D��<���3�R���k8�{?��̳�0V"D���̇@�������(UcĲX^�Q��+Q:H*�ǀ�(%��~�7l��
y���8��k8{�s�=�t�@�HY�P�d�a�K��-	�Y05"3�-07G8���6�P�H
�K��'El`��H�>����J�<��4��w��������"�S!}˺�/�^�֩�3M�aAտ�Ȏ�e]��r�L,[h9�G�����Q):�٪������)V@ŵ��n�`;�l���T�^����P�L�2w��nS������.S*k�4�3�eS���[]ڌ����Tണ�N<W�]!BK3�U��Z�?�+�sЛPI���Z(�;X#`��g���t��Y��q����{����-�����JqRm-����"r���M�J�H�jP�>L�l�Ғ��OOz����,]�ׯ�_��ϟB}��b��no���X� �T2!��[6�BK}�ϟ��3�C���E�b1c.d�'�_���s1::��TϽ�s���/1=3����G=	�6l�ˑ�Ko����q�j��	���K6��n؂m��#�*b���'�᭣�b��IC8(9�A��%����c{%�]0����B�O�Kg�L\n��f(���t����]��3�<f�IL����~�;c�x`�twt��u~�������b >N�w�UUr��ڎ�G�2�h��a˪5X�l=2Y�3c������"��D[�\�B��$������Ȝ��n�����F�AO=Y'A!V�J���[�}p�S��L ��\
oy�^����=��0�L�nۃ��I���_b�0'y�0��7E� ���r�e�����cՒ��-͎���cx�Wh����Z?A� =�9֌�/H�����nC�?�K9t� ���VL��s�	�u��	5b�\`pyKx�͟���x����h�D���?������}����4;�]�����@�:.�*����>��]�oއ����^H_���)\Ј��:Rj)����cPBV�W�����2D�x=L�ͭ0rR���O�''��.�F����/� !؟aJA�x��WY��P�u��]��,����WS�Y�,9�/i"P�SY�Z��	�v�M�)��-]���\���I?��aB��pI�R*d-P�A9�R"��A��GY*\\����l:�,�D�Y�H�o��r�9�iIr�;�N5�̉��Жz�~���x��!����|�������~0�sO{V/�T��bA��²�=+�%�������
�������l߹�����&l$��9y�c�ę��Ǽq�6�?�G>>�㧏K��C>$���Y/�ʫ���tB|�rn�+���%8Y=@����k��@|&�����9���J&��+���K�C{C��!�VHd��/�~�$�#���J�Aʞe=���Jua������	�v]�׹�����t���M|r�c��U���-%S��G���^;�2k�����U2*�!�."/!Ff�nܿi!m?&F�x���q��c���x�d�5br�h&�b� �ˌ�3�}.+�������r~&Gȷ��W�.B�3���<�h���;�FV�DbN�7�q<��O�b��;��ص7�p��Ii,ɩ�FE�8`�;D���.	��׮��e��K��w����\9�Bq��1����Ҷ6���B�_����{Q#�'�$�MխĈ�M!�E�������$F�h=�m���%�	��|�*\�ҋ������}�7���{���׾�9R&��<~���b���]�_6� r���&�ei߬tfv�%�+��B;��N�BS�O��L��5BVi/����$�j}8`[�Apb0�{��[0�����ӥ
Z�����2��4��H���!�Q���V�	�"A��G���R��d>/M՘UK�Y���u���X�q82���E�┩��A���M,���tᴡ�;jlo�nC��K�=��ż8�͂�5pI�mUz4�S�#�)�n� ŲZ�2�9�����~��8}�m(� ��V"��PֽޅÖDr1R�ð��R)inS�ڹ��s?�y�q2�ct�ܸ~���_~DwP����MX�сB&/m�c��v��A�.��	:�	quHR6���Bo���ܪܥ9����7	U��ڵhM���ix��i�|�m$���;qkhs�sA)3�F|d=�O����R"N���8I&|����y�E:Gt�����$�`?	w�ҥd�^<Z���<�S�/G�GƦŧ�z��f��+<�'.�f%�֒7���Y�����G�C�ֶ��]"��/\ �>+V���35x��� ��*Rf��n@,Ҁ��7�'{�:3ID�B(�t<A@�$�tY����u��T(�8��:M�^��ŝB�
�ᣵ��R���el�rh�#��]�v�S��/��>���E
�O>�8��b8>D�-�J#D�f�<�t����ۼi����ч�g/���B��M�ҝh�o���6����P�J�x<�	�x_[[ŒP�Vn�KvW�������#5�&��G]c�#���۱��}�o����o=��ھ���}�w0M{w��yD.����tj����xLU�-*�Өp�Z��N�1�
JuL\[w�q5:����-O�&AE���B �%hK8�0S�*��Q��t���iTO�aYZN�q"����t[W�D���H(%Ix$�06���O籤�EZx{iӊt��&��d���C��u�A�n��J.i�h*
��UqI��S�z�[]�4&s�Q�aq~%�³@̑ ̊�u��A�n!є���B ��M0��+�$��"Y�2�oU��.{$���ׂ�' ���_ؚ���[ZY���C�`�����������v���cc��?�k�\'o����{�r�yFK[;�E1i}��H�3���Fe�|NaU)��T\~�mr<^&�b������c�0>5� ����V���m�=��y�a��|�LJ��S4��b�J��I'��;�ۂE�FF�z�:�\>�l.E���
hij@'	r�B�b1���bu����ɤŔ+��(N$��CBv.��1�E$��ǜӡ�LD����z�M��rsˠ׏�Am�p��O�)~�/clt�ǆ$gS|�P]F��rIK;��y=��I�����8��1z�׃663��"��,���x}�<�`��L:+��c\M'A:��RPư�G¦�-C:��3bA=�c'�''Es?�A^z�5qc�߹=����o|���lV��R���A!�%˰j�jIAZ�>��ֹ3t/��}�}XL���aoH�~p���?�,Z�.�������%��ꯉ�)A}��8�mۊ��.\8AJ�'����n$��͢�����ϣmQzZ��Js������č�Q��f7\ٮ2�Jꠥ �Z��jY�|T\�*���L3̅�/�"h*L��m�*�֬u�����s�辴���A�!-+�3d�v����{� 79#�X���`~6GՅ�]�c��p�9��|ɹM��n�w��|���҅`�.�_��006*��:��w�vl��WHUfɌ,ꨢ�S��� Y���18�N�ٍ�-i�kQ!�	�	�I�F�	�p�!2U��(m���j�̫���	2%�
��
�9����CڡR��]~���i_�"�,��>e~��ͪD1]� 8c�7��mB%�} �[Kg��T�ÿ��i����s,�9j��h"���Ԃ�a�-�ϸJ��y��ѥ	�fg�� lKJ�}� b�R=Ӥ�������x�Gp��U\�x�K���D�$e�����ކw�A��^���s���LB������_T׀-+�c����=q
'ϝ���4)@�;����"��&��r��B�i��++�Y@¡Ü�ܡ�P!IU	���B0G�v�^Ǽ��^;@�gN�6]�Ka�p�<!"Z�X$� )<�Tq���������}�,[ԉ|�������HO�J&�Wم�[va���`��|��||��BMa���l_Bc�a��m4��҉9L�NД����L�ˊ������jGV�M�-4~��qQ@�+GGF�l�hN�x��A�w�c\��bV��EK�A�ב�ݽ�~�q�C��Jl���gx�@�{��Үt��x��Op��<��$)Z��~kIv����
HL̢1JkJ��.$���uR3�z�a�0#��E+�u��"����S�@�ҥX�l��_�r}7o�$K��CssJf	7�J�������ϰ�!��͋��Ǿ��z�1����ɝ<,A�:��vʡ�%4횯�uIk��Q$hmW�!A~ܕ]P�'9~[;�$]ef;�D��@]����؇)Tx�R!�FnLh���c8�+Jd��"��3�3���K��ʌ��"m5��E:�f'�U�]OH(`q"w �z��KDX�����؉���s2n7r�'7Z��^c#����1L&R(�xS�LJ$���VN&S=�kS$���,!��iBG��L��/��Ҽ9������e�;��8Ahiݪ��^�S������B�ܸ���gy�38��i�Rq�F'���:�C՜;�^)x��a���渡{%�Gʇ�f�B�����̕ �/ ۣ$9���+�v7ã�#���EȊ��&����xB�
�᥈�0������9Z�H(��_B|r�N~��_ڏvRPsl㽏>�Ԯe]=ط�~����ŷ^W��$��MKW�G��?R�qB�l�N�ĥ���.������K����ut.� ��mAzY\�t�;W�~qv��X�.y��_��b��=LcL�$$��M>O�:%���Q�H�>�ю;��8y��e���AlY�����gΐ`+�\|t��.Y���ף>ڌ	,0�O���l)Қ���у�N���FB�y$�	�gfS���-]��dDI`�O�;B�d>y�2�[G���T2/	� 	j�?"{=x{@�����8����Yc��y��\�!ËC{��˸39Hg[sV�?&�>o�Wm�l��O��QB�3��`I�/nh@#�t�xI\bnMIȎ�p(F��K
��p��ΉW�X����FQt)�<f���%�y��-�ݸ���zlܰAZ�KW{iZ�/^�)�^Rz���%���o�ЀC�å�+x��di��'+p�Q�vM�� F}���?E�$�R�N�����U�yU�ڦDt�RQ���K%��6W��4u����gb�r�}A	]�ͣ��d�J�bJ.(3:�RE)!��׋P�
h.J�`�&S�b�4s<���M'�����k%Z��0Nf���|17\E[J�<��İW��I��f�y�Ȓ��O� �\SW��1�Еt�2������q$�,���h��O��^���}ŸD��n���8�����-r�������IP�>G�!4�ZE�u`�&%���𜜋Y�x
CQ�'������)��������ڣO!��1:=�O/�&%U �nc!�.&��w@�W�_$�1���p�-� �n�PE��j�*�(|v�"e�)B-dbӅf�Y2Os��QO?�^~�0��6ף��N!��	||�!�Eh��㉇���>�HrR�H[���-��a��m�y��s]�5=����܊��q�s�JZOva�1dַ�\Z1m���#VD�l9;O��։��@g�KȈ91�!>r��O������w���K���е|)Ŭd ���p��El޸KI ���� w��)�qR�sXҺ�<�-������������t�KB���֍'�:�"�.�Mc���عu+N�8.�z,Z�KWJ|�]Z7����Ĩ(�n��>d�0u��W�'���OI��pޛ�W����'F����0EJk29�[#C8������,·�x�ҏ1=7#e����5��c_AKk���9���	'�5��c��]O��OJ����A{c��Y��0|�������h^�E�7�|&)Ap����h�|��-����krb��c��v+h-�e��[7��k��$wmہx"��?|�,��ؾv+�Cux���S��`�4'V��4���=��,�����|	߃�p\ �X�V�Vk*r'�^���.�+~�NbK��\yϦ�A~���"l@s�a_D�:G��t9�ed��� M��FF&�Ȍ
�����Uk�`��D�v�5:9�CtY��$
.!�f��-��	Y��)B�,,	�L�佘!�%�GwK�Y�t�$��+�v�d��4�|�_0Ȇ���gHk,�b���#���ǐ��3��t�":K��A$�<�V�_H�r��<	�hSD����D�����N#��B�ۏKJ�+K'3}	S	m?����% P*q�����bhb��Z�$�;i��0=1-B�[~\�|U�<�;��J�˺'�Jh���
g40o)�y$h�oG.�%���%�[ D��3O��O��^u�-�@`r:AH�8:u��G���˖	����H�a7voނ��m���52u?"!�.����b��LD|��4m�4���)�e�Έ\bL~b	៴br� YM��T��Qd��Js��g�2��8`bof]��\���ML�`ZA�M��Hp���C?	�%�=��X���<��?'��-�7�aRA���&qⳓd1��;�����q�L�ׯc��U�ʣ����ӂb9�f��ho������,	gW�ٔ��
�s�rϙ���O��g�9ګ��%�\����]�"����!�����Շк�·b��-.�x��]x��w�#�̈ Lw�5�����������������#X���zV`||��<A
��Э��)٫��V2�W�}XA��� Y�C�b�Y�ӹ�8 [D����y`t_��J��z��ٚ��w/YJr����;�L�v`zv��I�.�q�{hUw7Y�q��)X\�� ���eּ�mx��|��I�� �i�"��2��y�Ǘ�L_U.�!uE��~���D.Ku�$�HR2W�0�t��x`�.,�X����t)2"Ӌ�;*9�����s�����.��T.E�@��÷/c��
]�BN��L��mn��"��	`�bѥX�z��gG�$� TK]H�0��%^(�$X������P-����/� �L���,H@�&a�cJ�٤�@���	�p%��l���Y�JoJ�\���qR<>a����p4�h]X����s���qә�0q�[]%��NK����6PvaזD01ʽI�ӥ+���qa����I��0r�B�0�@Y��㔮�
tZ*�&���*Ō���	
o��\H�"	�0w������߼A�҃=���O�cQc��1<1�>��w�o��8�]L/���Kh����Kh+���R\�/�ӟ)�|��c(F.�Y�*��<Ü�/
�M(N0�@��Ę}??;��(�0��N�+dr��T !�E%���O�:����}7��V+��|hoߺ�c�Nb��d���g�ŧ�!���}�>�D�ݏw�H�#��P=��-�t"N�ٌ'~C�#��z�j��~�0�S��t�D2���U֤������	K� ���Jd�|��m���Iy��%��%$�s�JaӲ58{���p�������a��?�s�����}��0�Ź���D��,����kFcK#�����PO���������a'	����}�=91�`\�B�1�p�4W�2C
����=��7����1ff1F�K{��~ϐRO�k{�m�FL����¥���҈����4��;d�ޘ^��us̚���?>L]��ڄ�zA���òe�L�'�c�z4:wl�H�[�*k��7���s��q!�U����}X���Ϟ�d|R̓��$2�9�m̑6fA���p}"$<�6_� n�^�1:��iuB9\v�hL��Yb����D����>sR��tQz����: ���%�a�,KJ:3-��Z_
��
]�b�+y��3�I�̝[� �O'�9:�ܶ�D�9C㟙��MjzR���a�o��##�]`rਭ�+H�pO/Ι�c�����ނ��7pm�OȰ9�M�Ĭf$n:Z�(�ݼ���v�z/�sq�t����P�gn9�e����)"�/Х�K&��As4��d�e���{Ŭ�=�?�Z7��I�%B�}7n��������e�Z�B�ٸd�����b�I�0�F]�B>k��E�l�
I7�>�(�X�[u��?��W�d�u%��o2#�Ϭ̪,oQ @ �!	$A�ˌ$��zM���gzz�׬5_�1k>fuO�FӔ�$RC#R") �U�{��{&#2ܛ�Ͻ/2���T�P���{�9����>��&��&�J��G"����+k�fS%7n�`(lԝ�V�33�9HV��wL�ù��8sr+�B �tK�8�oO_�A�٬D'Il`�8p�����A\�rQP�q�1$�pxx?Z��8~�6:L/-��wޔg��&(F�Q�{VW�do�O}Z�{	��\T�-��t�E���;���<�K'�N��ß��UL=S<���g
���Xz=-N=�?�֤��/�#��Ȯ��7���&����p��y\�vOH��� ў8�s.�ܥ��Td710؍��N1�-�;3�bkݲFSSZg��ʾ�A9�8�Ϳ�Z�)�c)����ܢ��67�Z�e��ۘ���d$�Js�I�q�#'O���~�SMXK��?�?��?ǩS�q��	�8(���aL��k�y�N��7}�7Hѫ3����Z����o�2��]#��A��BRP��8��1��Fִ��-�J���n*H��\Q�G�L=��'�h�+_�����4g9=5���%Td��s��^�!�C�k���DJ�X���skp�A6����mAbt�������J��v��-��Jmrt�-=��켆��`D�-��L�C5d=50��B	�3+��zf��jT�>����?L'WUmH�oOK�גQX�u���)�w��}(��������3R�|"&��U>�$�< �]�����a9��m�G��ٚ���wK�IђB��S�N�"F#C�ہ�X
9A!-��9�,ϐ���*���VYG�6�n��FfA��)((."���T����yc�RE[`�G��v� �ՂbZ�V�g��30����X�[������(R[�a�۲��D���T7����KdR@D�A��vA�-b�V�7�h�����ƴ��3-�0M$��,Z�a��qD�bI��;ǌѓ�ɏ��G���A%����+�56���U��T�D&�H��%
/f~�Y�Λ׮�1A|�bh�����.F&�c�/��z��)�͂Ҏޭyxw,�#�N�������1���zwn�ñm:�EU�R�
NV�4F�Jق�� h�G*��j]��w<���jT�z�\WF�e��>tv����C8{�F��ý۷��ѫNg��Ӛ8AJD��<'��;qw�$2�g'���i;UY�n��s�t��a9�F�*{`nzAMIL�E��ދ��vU �6�,�V�{�3�#3]:ڮ�T�n��5%F9/�ae"$v����ı]�q#�F��H�|V�?�S%�KYͻ��S��L>��j���h��j3 ���Q���Ӵ!��Vj�е�,|�1����!`�Ú���`��x52�
�&�
��<a��^��XR���n�(�#�[Z[䠵"*F��-�Q��NYߛ4�p&�������#�C�"a�䨈*iP�?(��p6��K���V��%Tkհ�.#媴#�f56�rpsb�z���_���̒��=*6�E��	ŢXʭ��|���r�I����c�d���}A.�l���D�]�C�{5�0'(g||B�SZǁ_����>���gf���K�*w��cO���],^=g�Ys����4π�tF���<���,�MadiS�W$����l6�퍍�1<lk��/U�Q���g����ƪ.��{�c4�)��9F,�t�f1�]��(��M�1������5A��|k	7�@<��g� s��MW���f��5�����J%4�~�g���=�\����V9�E�Rp�0��Q��.;Θb�Q;��9��AB�y�T���d{��_�L��!Ē�)�C�K� � �XxS�q^~�ŻO��iA{�*�}��-y~�GZ���c~a^+�Q���7��bX�@�8��:���uE�O=���'��������$}ŦiXa��yr<EL�艣��jŋ̴����t�+*�Y���AAñ��BH�$�����'?��W.i�ߚQ��a��9���w뵲�t��5�8�KH5��o�tL�=��gmz�Q�Q�TU�ͮig]Ti���Ҷmz0t4���}V� ֠k4_m!�A{O�\[6�95�6cX>gaqA#V� ?��Gq��-��9z\�5����G���� �@��f�_���d����~�O���v
� ��zz�[�
�%��t�ڻm;�����K�LSp�k�FD�)�1���;,�A��D\�rd�KSb�dA�KP3�s�s[U����R94�R�L��<o�ׯʁ�Թ^�.4�:H���c�6\~�}��&�,�����K�1\:9�O|�i,.�p��#(�Ɂ���.B��r�]�8�'��[o����P>�zB*�%R�T؞��q��'	6댣-��^^������J�2M{g;wi���+��n������(V�k�4<(db���f���y���5E7C]�8$�;~���z�0Ҁ�tW���ss�L.�S�R~�x��f�]���=���C��B0H�[V�;�;(��HF�K��zݝ���@�5v�C�?�n\�)�vG��c'�Ʌ9�S���cŨ������!A�3�:��9G,#g��Y���)�����cE='�H�Y�!�0!��5ܓ�ĵi�}�ܘ��6��8ʨj�yd�P-.,*���4+a���Hw��kJ$�J)L����Ȕp\ֹO��.���l{���k;��{��X$�3oݾ�Ǝi��L'��=j�&�#Ҽy�l�6�" �	���0��g���p2-�-�016&�ۋ��BoO�8�Qu�\㼬�7?;��aG����(�'F�6!�A�|��ǣXY�@A��O?�y�Y�|��EY6�4ɟ�e,�/h�K�S6���rYK�tk�'�;��T�N�WU��q��X]��"�����n8q�F�lp��+�$����4/Z��mp`�M�6*�˪6k�����Η��w~����x� #����zGô��o'U[���e{�.�#9F��	nnh��Q�"V���_a�d{3[Z��� �:��/hFB�� ��|�ܞ�ET^��.QP��3�g��L�7墚>֠x�*⭭>َw~�R��0��^`�#:v=���S8�³X)�07uO<pE�YF��
i��ʍ6
����f!�;����z�Z����������lmg������9��l�D�Q�i�؁�70��+l�mL5iVmYU.%�S�$�#^�|���+�hk�P��r���M	�����x��'y��R0�l��4g&���!��&�䘷$2st�-��c_ǹookE��(q�D-�"���kXYZ�A���O	�[�_Ķ���X*q��򓟿�)I	�'��`�n_�#�4f�:F��U��Ub��fP�=��.1"�F�\6�@=� QbX��r�l��uw�s"��2��T�|F	w����8!��6�S6���9�ۓ�b+C��8�eq��O�Q�
*F��{ �r���->rL��u��5SPd�ʂ>R�hH����AȎd��'�Nӱ��x�nU��Z3�|����k�U������g�V#;��������<��>aj���+"̀F������ݍ�;�)ۇkJ�O5=r\���5�+Ə��YY���u�;�,�h,�-�e�'T���iQ7(�!��P$�`�Ȝ#j*%�LH��Dw� +�{X��իה��Ԯ�K�ʩfV��H�����t?��7��,kF�A�}.�V�5��C�lCB��7�昚�D$��q�&�PUcݔ�����ȑF��H5!Vw��6d�g��5|V�� ��4�$�&�?���i�n9'�`Z>����`��U,�����/9W���4Ju.���5AX\��T�g�\a4����;��ֵ�h�x�%'gd���RY쑩9�r�e��-����!f<�Ķ��Ř�4K���*�׳�]uM޷AHC\ǻo����E��� "޻j%���vXɳ��r=�w�Gөb'E�s�}���� D
���{v�Ɗ�	洌PJX�w��ip�mp@ך�z�j�N���1AZ��r�Y�Z[S�P�	DQ�D J�������DGlItOt1'��{��-VulNE�Q*�#��St����.��&:ь ��Җ\k9~�:��V�Ibomm��X������v���L)}���%3�(��w�����(�:��fma��T+N�e�{Z�c�#m�F��n���h1EA�yGK�
:#o�~d�Y��f6���(�ΖO�x��]gW�2QwҶ\�Ú:�S19i�1����$2�}�޼qQ�k��#�m�[�F'N��k��D>�Իm��&q���V�����
!�ı�q��1��^A�}ؿoXSB���7���lmD�,VŐ�h�?d[�7$��c��kU�
y����
#���v�޻_�i�̦�^ȡ������}��g�TưD���Rۡ�]U�G0��"�P'��/_��~D����!����`&���E��|�SO�ҙ7>B}�r��4�3߇=�9]+v����&U{arJl�C3:;%���&�B[2Um�Qm�s���e�:b"l���L�,'m:�i��}���W��(�ܽ;��ƒ�^���g0%�PWT�s�8�Y+�9	���lxh�Vn�{j�<�x*��j���
d��G�ML�L`�7%�-�Y�)G-L�de�P����[�41:��m��aw�[���֭�܍�h��Fx���'�I�;H�M��ƃ�ȱ87'#/�q�]��ˋ׍NH�<#�^yM[k�CU+�\絥e�t��!x�C�j�r+�V�g{w'����2��J���{tcl�f8�]2�M"
h�F#H^jE-%H#���������%�Z� m�!�'S�f_;� QCg�zJB��Ck�EN&��[K�ixp]=b�%�>��̖v"�9�Q�7(k�N��u���K�9�`eeIܚ"��v��}nz�M�3�/�\(����+��g�61S���LH�=4,�]P�|�.\�r�l���1L�0u�˼�.q0���^'��C֍�~�H�� 0��I�פʲ'X�Sc��nPVŜ;/hϳg�"V��uj��=�S#\�\.��>*�Q���cG������ݺ��cL
6:{���p�c[+N�J�R8~���e�$Bu5�R�+�	NH�� M�9��y׈a�����̏h4�yYQG�[P����D7���yf� M�L�C$�&0�ajvVS"��gf���g3P8���Z3ەE��T�����Z[
�U.k^�iZu��+V�O�Y�.k�>(%���ܱ�i:�$��>bG�yY^�'�se14��Gp���8���Z���qS4IX2?;o���۬㴃��`Ŏ6:�U��Ż8*�uP���&�)(�j�PI,߷d{�3���Y68�0KY�S,���N�l���I`j��
y���sI�7̠R�ac.�F%���w��r|7�
���Y5��" ٌ�N�	4����@���ݠ����C:�� ��W����Q�k���Ȃ3���~S�����4����>.S�l�����!�����wiX�F�ݿ7�^GR��$Ԣ���:>>)(���;,��͹����s��kH&4,'M+&�'?�+.(ReH�.���!2Ԥ��Ɵ!}Z�pzsCy�a'����U,���.�7��/�C;���f1Ђ��&��WiœR���쌶ò�F��]�B&''ĉD��֪��X��*]G��{�_�������S�#�������d��SO>�9ErY�_�V��d�����3��M��i��KM;<�OC��U$Iun�*�LNjaҳbL����_�?tN�����r߰֜���ls�2|$k^��cd��C��?j�k����8�444Y�i�wM��X�d����[�n��_\�Q����QUw��ϓy]���D!�DJQ3�]�o�z�HL&�SD673�y��l�!F#Qtt�ɟN��+�eC~/��A��*ڱiI�c��˚8Z�G�y��H�A��H\Sd�E,�>�f���^���ܺi%6�X?Wπ���@p��ݶ-n�������F�쪙��#�Y��l 7�jM�n��UlH(��z��059�C���ы!����yP��q	e��S�� ;4X1�v� <mLx��)�xh�=l.O��3�"��i"p*F���y=�;� �5�\'V�3YѼ'�-GŔ٭W�Z�dAˈ6F���Ωl R�`�}�����O�>GP:��rFca��b�#ޔD@<t�^�Q�P
2�-��W�6k$c�s��Y�('*=���E��!d�Zѡ�;o�F�4USN+�e]�9<\��2�4H��J;��Ѹ�4����#�������%2���2ʎ�TF�����H�2	RMͺ)W�W01:*d�)q(�ul����B��c�d՜i�b��Ҷр���	�J�AS4��I+)(2��͜��������e2?��.�9EW�9PTћ�I�U+��T�@ѐ��4�!94M�j��0�Ïqԉ1����c��)�%�L�fYC]G#��\#Q����1���Ѩ�JyH��O63�W��'�i�f��;Nm3�9*�E3�_?�X_�v,C���xL�A�d���<��-m���2}����d4�87��!D��(g�+����3�8y-�1:�����'EóML��e���)s�TÚ�"`�Bc'D:��^���&"%�VMڃ�ڢF�!M�����-V	dhp�S^qzr�4�D�̳��Qg0�Z�Oذ_S�����p��Tn-���p�VY�?LǂQ�WDj��/��n+r�d����nV��j�P�@��gKs1X��^C��9\�z=-=޵W�/8Lb��"��b �F��z�b��I�XbXם޾q�K8���W���PT'�f�	�z����"�l ��?�C,�L{hF�e�,v1ɵ�͜�v�8�e5G6{4��������H	�	P�E��Ym&��ؕ©�	s�4�0�����wP��jkA�l��ZZ�uT�<s٬>�\�4���\��
|�Z�!'FvK��Z9�cH*�;���M��QwTB^#��h���"
��������$
Y��/�z6���{ M��вU4�#h���4���$7�,+fj�ڟT!#�^�"��D$S��7sy�w��%_R�.�$(�B���ю��dŉ�EU�Jx�fJ�<�B!��g�\J9T뛛����C����}�JԖI���k����b�.-�C-X|�j����ye�PʏT(?]���zUR����fs�ʀ���4K�٦��Ui��DU�YXXԢ[��zɾ���V6�C��*
�,-.
���޽Q<��bDbA1��&�y�SN	��Ю;��-?�yqD��ł��G���\?�4�[X�PH�H������,k��{+j�A��-j�e�)B�Dw�eV��'"{�p�Seg�;(���5�G0u�6����Ygx��+�iO[Y��Ut��BNv2QTD�k,睼qW�Y�D��ig�BV�ޔE��#�!J'FCL����f���|aUӑ�o4�%C��X�0�C뾰��ikA� ^U:&�,��f���Ng���7�X��_�r�H�}m����?g'��[q"&zӲ��A�;�w�]��a#�oC؂ ��T�Չ�)L���vAc2����Jg���A�����haK�x�d�������w��ǟ�؛?��(�+��,a;�3�g�����[�0��YF!A�A,��3�����b�X���xeq
^X�U��X�����L�g�[Og9�^6��]C{q�ģr����r�tζZ�WN���j	�K���6Q��ء9'�b
|�QN �EbT��n Ƕ�xyy��-�88Ҟ+=PD�e��`~�O���eU��gμ&�l�EԦ]{��N��G��DC������T=��}�H���:f���DB�:P���'?�dK���g$R��w]�!��`��Bل˫K��d�hj����-�9QS1h�D���Kv8%y�$�id�A�YJRKH��P�Ё�8v䰦�VE_�qK�2y�V�F(`Q���r/aq5�5���Se+5B����E����#��$�`�i.�JE�A�F�C 5��L6���Mi0���<b���Y�wu�W)HD�ҥ�>��T��-}�d鄢!wu���Ĵ##�#v�b�D(YYCrdW�PƓ)
�i�dX,�h�I1TT��m�Z�Ø�l�R�D�d��,.�be}��XF��6��!��BZD��4Y(�}��_����4~��)ڑ�ѱ%e{mJ�>SVLQ�&�I}�ܛ�\�6aֵyҀ�DBm4�ca~�g��JI,��H\�E�E}��}��v�Y��>��h��j3aS�N���e��(\Ơ����|9��oB�֥<�=������Fo��\6�*'Jf7�K�B� �"0���Ǽ5�U}豎� 5�ng�	ZI�Aa�eI���Z=�:��54�ܝ�r #:�ӣ4��*| �Eҏ�����������4!���򕫶Pc��-�÷������1�)j��ϛ�����W�{�|#Fe�v�ЋjSq����,�5����ʅ�
N^7z(��j\	lf���V$t+�njFj !�V��z!/��E/φ����ʁܐ��.���3�E,O6���4:[:�M�����(a[ދaQ��=rй��<�t�fgg�07�m�͂��Mx
�xn=�Fڍ����6���������X�Ѻ���=��(�1Ϝ����}�$����f�lWB0)Ws��)�,�,봂�����T�1ǑgJDg_o~�Q�����;��ޝ���u
�Ya����)e�oy���Mr0S��Ǔ*�^�7���u���`iyQ7L��1e�y�`P�>�"~����<���(ttu��[�*Sղ��8=�[�4���,Ƥŧ>�i�<b�Y�b�'�&%2)Yc�5q8;Ӗ�gn�Z�zI��v��7���^7Z�l𡴥�OZ��TB��2D<3�^���J��*�0��ᓝ�?w���ռuy��ū͍u5��+4� 
�[�����)����^�g	���er�ᘉ��o���X�^���(ȭ͘1_\���m��=�f
��NP�	PS��C��c��7�6;`�<|�[$� u�3�hݑ:�$���꒼5�o?ͫ7�;�c�k׈YT,�]�Tt�!OS0�־��P\��k���!1�-���d�Ġ�.	��r�xh�DC�������\	ݔ\#퇟4"l��ܙ_D\¿%��p����x零	��O䣡��l G�<��/e�R	���51��*a{�YDc���g?��W��(�7բIzv��O����KJ�v��Hcʅ�� )G��⩚7F$�����`�H@E�s��se����@�)p� i��F���F��.�Q^�i���tt[j�i3e˫��C$C��]��Ě����9��{�)U��L2���ïhs�<Ф�0,����cc�@3�WCOZ����{;�Ko`uqA�&���,�U�9��9�C,b4+��b�<�rh�?w��bxp�8ҐR�x�%Ax��o�5a����12>%�,��N,�4���"@Mw��<���c��MC	�_چ3J��������r>�,�ș�����TJY�	A���D��G.	�"���*_[j\f���5��f����R�mhikUg�٥�9�lQ�4���7:���z��9�]����>q�$�We��D��x$�kHcX�2��Y��n�D$b���?\�xԬ����(�s�����(vaF����<�5�ca�$٘ԳO�#���vCC���1׋Ə���)����s�}}���3i���t�YH���[R��
 �/b��gp��v4��L��j��	�/?ZoX}MX[��Ӯ�Cɚږc��|�	�:�2;삺bWM����T.d�ϻZJ��wu�g�u^B����0C�϶ AU�֓t�$�I2���H�ڔ��O̅��VPzC9���5,d�p}~L7�4���b1���*���h���<���Wϫ��]$LaC)Pv��6R(SPg�n�[٬*^����Xmp���W~�-���OB�'!�����8�Wj>$0�!�*�-� ��	�HX(���
���qtv�_T_�j�Il�A\d�Ԫ��~A��_�C$�ҍ+8,H3N.����f $�UcrP��:�jC�C����E�;e�rcm*�.a+�SC��h��������=��r:�gtlW.]�����E�=�P�����~-G�L�Qikm�'>�">����c�S�~���)t�`x�\�{UהHkfaFյ�\F�)���Ѯb-�t�氪s�ȿ��'$d����i0�
�_8�^�&�i�7�jo���bT���{�E��}%���"_sbb\�Z�b��s�ڦLJ^L�^�Ա�:��֙����gd	Y�%JZ��M�c��9t�����c�Y7Aҝ
�hWT׀ΐўg9���hV�}@�{��Xu)$�8�w��F�0[�j�6g�Z[ZZ����٩��ajz
�}����z�m�CA5���1yV
:�Q�x��)���9���F��-�+Ӄ Eօi(��Q搓k#Jg��l`׀^�8Lq0��(PUGE0�b�(%��-���t�[Q�k*:�_{�ԋ�9�j�|�Xml&	BL��qM*�-��``GK�t`DQ�?��a���?�0N}����ja�5ήc���5��Z�I҂43�خI(�2�%A�ƅ��)0צBjʗ�n�\}?�K阎3�;��U����f�-ÿ�,�ge�L�̜τ*1Y1I~�?����fv�g�l5��nR��7���L�4ED��"E#�|�S�%_�##� V	!�9�ۂԱ�xj�6�g��}���"��������?�D�	�>�4~��+ؐ�y���ڽ'�g�<��_�~��uܽ{O�a҆�1�b<��FTy�Fʱl��jlä'�q��Qݰ�##�_^V�9�2� ���LAL��c׮]��X���K��1"T�b����⭷��`�6������Pg� �'IB��ДE�������K�/c��~	÷��믡 6�2�D�t;�a��2|��R�amcM'�F9������̊r�Y�Q��:t�"��T�"v��ۣw�	}��q��w����x��9M뜻x/<���(ޔНU	"gy�۷nj?>?k��A�T�jhj�������\���kOs��fxv�^E�[�sb`�ݹ�{1"jR�����U�����{z�a�xHևF������f$"�%��蛼gA"�[��`߁��Ȅ\����0��t0���*P��'�K��5Ȥ3��0�����r��Hoe�����t�pԤ~xX(��(G��i�)ۧO�<��O�Td�%rB�@�9��AJ[@IU��ʖ���5����exuF���\5�Xnp��R�*L���)>hh�_��s�>]��`�vU��_��6ݴ����)�Nͨ�� _I큢I�W|���MY,��͗�`�� ٧�p/#`���c&V�$�]ߟ�q�ldp������� L�ϴ����am&w��%�V���LB%/滪V��(�0��"�gϟ�a�������Y��I��X��c��c[�� �Ÿ��s�\]��[W��n��/�ԡv��.J����6ŀ�1���Z9dEGu�RH�+Fc�����k!"e�X�)�.��-��bKPs�}�p��Ax�����C-���X:L ��ݚ�.*�`R����BY�l�>eqB��IF�Z0�,dD'E����|��f�n����+m!��4��Q4J����V���u�8��k||\[yc��/�=�k��c��a��TA�4�\���U�<�m��1#�8������]Z^����i#AK�A����F�����q<&��\�k������o�^]�1�g�(ly}덷4�MU���5-~�*��4���՝�t����9[��n�RCh"�R~�(α�O��{��w�"*�oais���5�Ԟ��,�������DƉ�&FƱgz��8�;���Р}4Z������J�(ƞ�ڲm�(�4S:��s$��) �����i��Q*���{�iK�d�I{dC��m%�/�c)왱vK�"����l��A��m�����YdƐ�޳�8[ �$�\]��;����6�����*cNK�3�|4�Xzm�oF��>L�	�75.�d��/�M
"hnV����c���@Bm�U��G��l>T���݀�Wf��3��j��E���N����3���)�~�����6�1�BCV$��i����ҩ���A�}���
��ڼ�ks�N� �MO�΍�7�O#.ޞ)���b(˸r��	���8`�*�^ryض�Mz��/I���&���>9���@-����Ɔi��(�h�ac��I���}D'Y�m�u@n��4$�3�����l��_�K�99=��5�;�{`�o�������	�?�0��uh�xnvA�3�d_	��[U�w�,����j�m3�sf>A�yZҶ��%mq~fJ�K�DJ=�-:~;kTܤ��n
�L�1�w����{��.({#�)d(��a��o�#�b��ﾃ��U}/��Q�$�UE��*�5�~�t������mw�
Ce��<��΃�) S*(R,���a���+)����b\9���I���;Y9T#H��tnw��U���ގ��A���U�����3ￏD8���%�>��
z�#'��ld�ư|�l҉��E�ժDM�\�\����Z�kς/�[��L%��NG �S���u	Ũ�:TrjzL���4½.�C]b�%`�j4=c`=nx.�(�էf��D}��Wͽzv���(*���F�{�>�U�q�c;���3τ�~᫖k��6�G�XU�����8t:��V�=�O.�	f�P��П�4B�7� E�[����m]4T�G]��|n̢y6�'�u�"]դv8�����Ni+������'���[�#(�O�8U?ש9��-g��}�����	�S8t|Y����N����*�[^����C�O"i��>�"^�� �M,o�blv��-���Vu4EC#ċ�)�rH�bۗ�!d[rT0�����;jH�&x�l-�>�@2�c9��Ϸ�o@��l�
�=sJ��,�.�xN~Xˈ�lK��rgǦ���������Yt
R������HA�D«���M���M��6��8���v��T?�.�4�Y1N,Tiq.��K��i��ŢYȨ���O�xƖW�J�oD�D��?���1�2A�72>��diH�׳���f�JK�e4,&!�Ʊ����w�Ʋ��#b�:��)������K��S�K�4��9B��G�j�]dE��֔���M�n�ҌT�T�v1>3���G��ϡ�Н��hxajａ]��qx�A��������v���hYmDcsڛ�06DIP)e:��#E̮/"%�9R=,No
��JU��"I������e��r�
�d���i8��'bߴ��L��,p>ׇ���8r���j����a��u�̎�g�[�Ж<��L���v=U^ �(a��Y���:��Z���L>�v #lA:�VL�Ts� �کu��Ր�1� +tM�R���yG�f�k�LmF��z��(����m���v�UZ��SQM�� <6g�P�^$�V�F����ذY����@|P>��7F*�k�~K.���_�3���J;&�=�d6�m;���ǃ_�5�~>�7���x6^�Q��z���Yڌ��3׿M$��G�Ù+��{��2�
Yt�q�n���ZA'�.�-"$Ϋ%�@��lU�2">t&�@U�ޜL��`��LM������ˤ�����Bխ�:�<��]Cp#1�;��?�(b+SPq���%5��{w�{Dؼ%vI[-�lJȼU̡7¾�!	�GqwyB|Y�K��VS����(��g�#��C9Y�خ<}H�gS���;G0Q�
�˿�:��*��q2򝕅9�S8{�
�&��%!,�yLc����p�Y7'F�!�W�r_�R�Ǯ|':[�tl��Љ�9�.L��JO�#���"l^	��N��y��Q��5��jN� /?��7VhJ�dʔc�Iv�,Z:V��1ȍ�Y����V��И��&����]u���ЕmV��p?a17�U*�Q艍�
�W����E`���|I�%����6�)��(�
Y�0mj�}���͕�|y�����9udu2frE������X�	����ò���M� �
#��c�(%:���2'��:���V���ϳQb�����k��NNְLT�M���kq��xf|�9�;ů��j�=�v�������N+Y����_p�p��v�����f��q{յ�T� ��h��������*��F�W��s���՗�ޭI��R�^�����u~�W����W_�?��o����g��-���������l�����ŴF��j�{��3K�b���=���F��羈�}篰&ޝF�-�R�O� �����=p�lb_	����i����Dt:�T]�=jv�ҥ˂(���مCG��!~��WpE�ݼ A��y���YܛEW[+���U������:�f)��������´�{oNjuz3���(`��,�-�X[�d�����lGu�m�	1�A�BCNb=s��*UՎ���dU9L�kv�����X$��ۘ�-p�� �t6��9DyAQ�g��xp�>㾸�&a��<W3&��eХ|�CG�aqe�x��E��V�H�(,�[:z�mH��&i�R)�Zh�4�Z�e�]���3�S�0HJ�O�;�ƙ�(m��Uz���'�?d=evw���ynq	�*4�������H:Շ�13��S76�򶱲����{њj��ǔ8���T&e��r�3� ��Z3b��6�룴%���-���M�� іL����w��P\Z��Mɨ�,J����O Mj���g�㿠Q��+�Xd[����Ӡ�O�d	ktZ�H����?}�cs�~ܱ6�O��~#[�W��c;<��tme�7���s}�|_�5If�w�b�������J�+_V��r/�F/��>@�����ש�Y���/�S����3�T�M/�����3�6$�������g���{����e�s�{����Z,���<������𢡄r"��=��������IgT�-�"�уH�I���c�ib\{P]�][��l�c7��ɦ݈�bX��Ez#-����ն�����v��9a�A�𥈃�9讄χ���_KQ��<6�[@,������55I|��0�2��W/��an��o�r Ux��UU�hy�:� �c��@��cw���k��]\DI�t-��������*�����6�ah>v}}�v�CW{��M��.!�v���@�L7m!���?��ߺ�����RH>�G5_����٨s��*����UuDP��`�6�f e�
{Z �����m�]*֜	��
ח�nc�#*�rh����+G��Ԥ8�--�-������GO`����ø=vy���s�Z�^^�ݑ4��!�F�*jyaQ��m�7�+6����Ց�<�l�`���,�Rs�*Gi#)~/o�<��R!L.M�ڵ+��F[��w�&?s�<r��!Os�&�i��W�@U�JY�6�X��4�S���"�������S����_ٱEjN;��A5X��<";�j��Θy��׺�u?7t*��pO���!��͟O��A��P�ը��U1H�G�N=�����8�^�~ԩ�+�b
0Csվ����zP���A���[��_�y�=|1��`d�˽�g飿Ϩ��_���7d)����(���w?�%4����翂	�.O��|zM�Q"
��3��%��aFxF[45��Z��#X�fH!_:+�f�r�U%�=zDf�/�ǂ���V���@��Q� � o�.���8��0��۱���� ��RVS�=�V҉�Y��|��Ǿ=C��'_���4��@�.��1:�O<�,�b�����$�]N&�o*Y^�78FR�*g�d����P����;�x�hH��Z���G�/�~Yͤu�dJ�5�X��4�w�C�<"(�k�S��{&w#�y��f�&h��]��x������X㨚XLXJ�/,S�  S�IDAT���ͷ��g\rTH�����Lqة�2���9fj���?QX�ILH�C�U���23�� �g{�X�,�`\�-��s8`Z����$��u�`�|�c*�����[�u.���эFJrJ�@����G�37�	�ʊ�Ӵ5H�Q�ye"s�T-K'�G^.�`���T�!z
�PՋ���(��fO>�<���q��{ʣ/��t�X��^Yu1*��.SN4�|C
�ƈ���:�8�H5���um͵�A�������~;�/~@ŧ/XZ�^ygc:V�_�`��2MSZi��-�i,�F��Z����Z�L�u*�I�J�����p��=*~a���0�`�joǲ��1���ͳ�;�ў�Z~�7�Z~�7}i����tj���7�5{�N�M���3~��?�s��j�E��.���������'���=�C��������&����0uxhђ���hXS*:^.�o(���Ϊu,zJo��!-U��^ ��hii�R
�s����r��v�RŲ��U�����ѓx�'��ݏ��37�`bu�P��b`����Źk��_D_������_�|�{�����!_���H�����ަ{i���+�s�U��rT�3�םc�� 8]!`�*�,�Sk�Is��l�<��G�*�bS�qd��MA�0{ԡb������(�|�)m���/��-�So+��l�H,�m1v��Xn�o��*�� ij.��kS�ډ���b�͕����3d!X��j"#�PCL��)�H����x��g��ԆiY��o �Q	��g@Ԋ8��W���ǟD��O��"Ff'���oj޳-�@�rd��eR�p��*�(6�h�4��8�P�(���]x~�õ]x�����������Iq�R���~��G<�����Wϼ���M����m�S��0���L�0�Og�5N�rh)�S;y��/`�{5�W{T���Z��;5����55s�Jq��q�_��Y�L�y�c���e�O�6�AP��~/�Շ�NM
M�zצoM���m㘰B��lnӳ:
�o����TT�l�#��V�7P~���}����r�kl��A�c}lk����n��k�Ӛ���ACoG����I�F1_���������&�<t�����XO��^e
�=�ԓ/���k� �7D�!1"�t�5�P'�ϲj�ZHY4��K�>U��Ȧg&����MkgSϮ��.���{{��Y12�w�O�{o]G R㮵I�t��eM6W�֙S8����>��Z������e�/�a��� Fd��[S�Ӎ��P3����V�y���	�l�3�EfZ+���Y��5�P!�|i[߻���%toK���?�ށ!q~��O127e�N���X��}x��5�z�}�i�E��ǿ�G����w }��7�����{i������H
���Y���uO͎t}�Ϧ��OY��=�x�'�g1;+{��_��o��K."��O.�����2,�Ʈ���k����k）�y�Kh�����;�=�r�&��S:sh`�ݸ��Ξ��?����K�A�>�%�c�{F�}�c緋���&���x�\�#�Ke�Du���tv�������#�U$� 덷_���JayO�A	��� �;����Xv���fR��h�9&�`��1��S�p�6�r�ն� M�~�:��⾜,�T4JoR)���!e�F����@e�|�a��1�!m�3�_�$*�;;B���McMK��S�W�Ö������P�l�@"�;Ƨ�W�Q�Q?���+����Mh�����P�˫��C��,�~d{��|�3������۫{m-���ג��G4�;#�_�1~�S_DSC#^~�E�]��o��x����i�3[�N��B&S�nft�65x� 6�l��l%��rXc��r��HS�<���Q@��Mb�b�8?3�c���/��A(ތc��֏~$(�@��}���#K� ��͟c�� ^z����A�쳟@wk;��7�&hl��^=ê����5�I���V����� �`�\Y~����e�&���$_(��8���UqJ�H5'5�������<���ڵU���n�s~E%/��W$��#�ۉ7V���~[~w��Eok���m�;u���ލ�b	��9l�ªN�&4BȄ�t�%�ɏ;*8�ۥ�M�����|\��;��R�������7����/`@�ɋ$���O~��{��6�BS�!�����F���x��c�78��������u8��T�8k��Ņ9�#N��O�c�=551�c�(HΜ�W(*/���vp>7uzjXLJ�Βч_�f	�uݸf�xk|�}�8r��<�(�b~)�⇿|YW�W�P�L��*u��3�pDS�kЫ�к�s�2	j��>��Ca�x��S�ɔ��q�����z�6#8�1�I]wGy����6�k�1�������Z�NH�D����4]���F��4�Q��ر��Z7�mT�R�$�a{�����\�^s��N��O#[�~�֣Jc��{�n`ڃF��%<�U{�Wo"�����|�}O�B���L�7����|��~�F�~��;�p�� *(+�{���C�����A�/<����[!!�8.߾���ݪRU�ʣ��	QꢺF`�tVUz�mH�n�YW��i�!���E	�gfTm��������i<r�!|��>��C���%TO�Go��	�Y��L���b�ڲX�|^�\�׿�m4�;��#Oʽ����GLF��_����+�)`O�G�(d�
�YN~u��^C*��	�W�` ���ek�|���6�������f4��*���ݏ�����H��������B�~�u���Tm"}K�bfc������=m��hnǿ��Cs��tN�a�cniE{G0:2�d�It���-I���:�=o6�k�&5F�":-lf�4$p��%�8~�~�+_���K�������[nE�I��Xcg��gK� �|����=��9��{�����ox8+h�;������E��}��طw�ʟ�Dk�<˓����*�/1�쫡*JA�a�,e$�9��fbk�Af%9*gtjR�?xPl��:�g�]�����KI�VUk@�ju^�Sw�!�PR�\a�Y�k�|�v��Hh�X�l�ô�u
���i@���)�,4lV�����F��8>9�t���c�S�*��&�I��
��(g��#i��۶��4 }_h��N���d�3�b�B�
��0|H.����+U�$o�֖-��|�����Qq9��U�U��Z��|#Q�����!藭`���������ߨ�]s����Ϳ��Sg0����>!�ܟ��/��Z����V-�S]�j8���&����D��8����<q�Ch��$���Ĺ�gq��-ݤÂl�9e ��Um
�4r��Nw����ֆ)򹄂�h!�Q6~��G��G[g��ᦠ@��?��'��3/`�{@n/��|��������Q�@'���?��7����=�O�/���눛�GO謭�O�?������wpw��rj��߇8�e]L�{F�QDq�/Ķ�*M�G�'%��N����J:�-J����&�E���C'��Sϣ��W�AS����o~C�4�N^���Z��݇�)r��U9�.޾}�������c�+�����7�3����믿���Q�+��`Q�'EStD'�F̔ �e�L�5۵U�Č#"י��R���h4��2����~O|�)��Ƶ��������Ť8ȼ ?'�Y1k�rS�d+�e1~���[?�����:��ػk����;�����[o X���Z�B:�C�8���˴�io/������m��耔]N))�1� ��Q��m��׊�56*N3�b��NX�-�7Ͼ�o��
���c�l�A�ac09�đh�c�Kh��(��!�����0�r=t��#:>JLŬ
bS�r=yF����B}�{�)΢>����$�$��Z�.�E����C�<a=�tբ�bSVٰ���|X��7n9Ivɯp�}$�R���@z���ʴlP���o�f,G�a�6{�iˊv�s��0�\Bu��x�Ns�'��ir���9>��L��qw� d���ҳ����}� ���o ���-Z~ �GML�7�}�}��D ��B��o/O���������ٓOho�C������/>���NcvlM]x�䣸{�֖V��S5��`D�AM�¶����u�����-ETI�qΥ:�'�xR�aW66BX�e�_�����_ �tF��b��>���ԕ���<��7�+���KA�'9�O<��^�{�=���[X�YA���ʘ(p�a&���]jq9����Z�<���[���E�m��[P��#��+7��N�sٿ�0�<�F�g���/p��e�Beq^!m��a3<q?wjS^D�ˊ���_|W;����-�Z�I|�˿������ϱ�2'�˕��Wű��2w%��dt
�@o/6�4��X�����Ġ�Z�R&S߈ ���%��=��GRyΊ������(��U��FCW��TM����-�,k��7/������Йl�Po?���k�����4޿rǏDGG�MM�s`��#j����0�|	ꈼ�]�mhZ���SI�ӱ�E|L"�t&�����i(Tۻp�&��Ə1�^@!X�n�PD� %8J\cP��G!rY�8u�#�%�n����`c����{W5TJ�l9i�R�Vri��/����I�#'Z_�L�Sq�tD�6u�vГ�����Z(B4�f<���X��U���Bj�$J�&3U�G;1�Ӆ�T+R�(��!���� }%'�kikc�Leװ��u	�2l���T!�Z*��8nY=[U�[1�5�}�,�7{ۈ���異Su-[Z�+��W���_G�}קo<X����W�;G����HL:��_��k��Ʃx�0?�t2������aia/=�q�T�p��g_ĉ}�0>2���1���i�55kΪ���wj�:�B(�L9?���Am��{�n�P�Ι�0�?��?~P[6�w�EK�EKa��ɥE|����O�}]�����5:"���3�����UG%����$��_�?��O}	/~�9qa��B_O/^x����cZB��մ�Rklf[eI��ᐉ�6�6Q�Hw�}#mH�7�`5���!��u'�?�S-����jB�	Q]Q�[7��}�]C9^��1v��ı.y�j�֖��5p�{:X�k�Q���/�6��;U��#~���\�tV�7��el�3j�ʥe��-	�fȝ�z�v.V�	R���M�Ȭ�q0�|�3��̦��jjH)�$��������.M�B!$F-$O��jځ�+����U�T6�t�϶d����ϔ�/>�����qa��g����~����d-�QΖpb�A�v���WU�%&�E\��+�I5�I�@[8��VN�͋��mo� ΞET�=�^�Rͪ˻%����g���I䶂<�V������$M�iE�SZ�mM1ٻb�;�k߅�p
=�mH��"Q��k��K��&:�
dEW�[��o�� �����א���#����T\N�`��#��(\6kY��N��Q�g��m��T��������D�p�78�;�=-]�6�)��Ƣ��T��x�lE[�p��{z�X����2���Yټa�����f�<Y*�l��[�����W�}�_l�v��]mzݳ�sv�:ne͸=` lF���+�������7464x�[oE�;�٫q[��ǘ�������W�������/����#"n�wz{�=��aj|a��r0G��T����-�V5��FZL��h��m��j�~�g�{ϰ́�y�~g�˳�������e��H����PX��+
��xە�)l|}_��_+{�^���-A:r8�z���=�C�O���]ܹsK'@���ؽF&D��L��*��/��?�Fvt|\�n�Q˶���2���]7��ë���x�r���|�V��c�+�������6�nӂ<+:�37/"'φ�v�oH6W��8��:�rYP���.#%מH&4�^^]Ո0��A��/9�M�:�:�h5�����sOah�^&!��Ģ(�=�_�����?���]� �:��$�+�L�A3D���0�Mc�ܶR��<RŏO����?�wd`Bb>��c8|� ���aanN��:;{��E����gW9]b���� ��FX:��%u�d$��98�q�L��X4�ϔzɿ�t�
�ݜGI���D
1�D�4�Q���\�D[9�&�i�ކ�Drh���M�#k�����Lqjz=`r�q!r�B��܀��v�l.���=\��bY>#2@T�O)`N~�[_��y��E��7`$R<��W�l��ll���oAk%��h+�ۏ��{�;�+�F���M������l�̬ؠx��X34v���s#8-~+����Uےk�����=e2h7ϾHve���Ϭ�b�����G���L~=hd������ox�}F��ۿBY0(���w��%�C����f[*z��a`�+��;�0�8��=�)<���r@�e��l�Ǟ@����Ξ�	��0�xD5-V�ٳ��dx�M���ցT{����=�nհD6%�z�6^{�m���)l���b�"%e�hޏ�р���=�W����6�/ߙ/��W?�..���������� ���".��?�z�����*J5ڑ�ca~.���zZ[�����)	��9t��i�F^,OG�
R˫��+��'l�0���mM��V	�� '�Q�?!ʵ5\��ʟ�W��ƌ8�e�"Ab�N��#��1���v�=}
3ӓp�1�O�<����N"��x\YcCR	�caJ䩧�C�����FA���̣�x��Y��/_ǜD���(k%�z��Ҭ\�V�
��d�rp�L2�!�{�"fĘ~����G�B��	��vkF�hY%Ϟ;��A��4����X���6�Jb��51E��:	�eM>��'UT��*UOE�Y�������㽻�VJ���TW6B)Q�}�Cej ����r����L�Â^;���hooQ���&�
 Q��m}��5`�D�b��
[���D�L�m&�S�c��K�GZ� ����Dl�Q�j�y5D�oGĚ�b7t%��j'���އ���W�kB=i��43oȼ��Up�(G�3)�������܄��n�z��.�cUB���<P2m����Nӄ��m�@i���P7�
�����3��1��ڑ0{���W����������;\<���q�s�~��GL��8\3V��(�M"��Z�w^�!F&���C���`� �hQ"�)�3����F%�
k�(����0��[7��ÂXN>�%4Wz���0*ɩ���w�����0�4o�U�3U�AEY&a��oZL� J�T��������[8���:�a<v�am_e=<<���W����LfK�]�K˪��� ���Q�����a��}x�gŀ���XA�����{��x��{c�J��*�3t$e���+������������oh�	T�˻���_��K7�L��O|O>����dR�-����̙S�{���(��h���TBg������1�o?��8����=�9/��(bs��%����0����J�qF�E��L�-���Z\U��Y�:���/�Sl}��;_WJ�g_�4�t�#���b'8C��._��A��R�+kX[_Wu1vxQ;#ݔB��}�߲=��?�2�F���ϯ,����\����w��n���W=��$Q�+�'m��#�R�cMx~�z�D2Ԁ��A�c	�Vߧ~ڂ�]]���t�y����/o���;�����Y��EQ\D�T�ݴ,Yv�r;����#�*��S��R�T*���q�؉%��bʒ(R�D
 $@��`�����{���~3 �3��������j�,�؃�Y|�k��}��y�l0��O�HW��Ը��֪��;��}L�l�U9Zv����|�K���Qϡ��*Y!.F�PDT}wl�B�*%@~�tLϫ��햰��o{ժ?��>��2���$V�3��9��(�UI��eE/n<���7�LM)�s���P����b>�	=�y[�x��Iw��`-���#�R	�I�sמ��6�����7��g���o|���/�HhQN����?��7ހo�巸b�xV�d�H��y��?����W_����7�ܥw�������:��o�]�� z��D\])���MC	w�e��Y0R�Ip�����]�������s������S���g�'������_�x�W��ٟx�5+4q�n#�om��������WU�ǻp����r޸pΏ�pu��E/���x8��ab�mK�j�<�LV/�&�L\��a?����5� �G��_�����~�~�x�s/§N`��"��[/C{mΝ;\� �NEIS��x!	.u��_�*<�%z*W� b���D��o���Y��q�^�F,�	�
�����ʞ٩+Ä�q�lV���@�3a"K^�����_��y�������8v�(���#�����'p��wa��	h��y�0�:�nl��˿�����^����^�.|����y/���O�꽛0D:�G/F)u|���z-l���������L�_��s��SЫ�p��1� ��hQ��e�Y.��L5��N�`Ed-����~�y�\�������]�v��E��s[Z�C� 5䣷!
	��cf��	�=����1�	��Cp
�~���ERLUj�A��U!�9<G8�܆Us̋P�c���^MܡD��j	@���#�n���0������AW&96����4'��=��g�Ty^8�N@Lb.�4��5Ԉl�\�"L��@�+��=�a��cB&���U����V��-x�̧��/}N?�8��,\�e{�E`ޭ]CQ���*��~�]����m/]��4K����W�2���MSPjEUUW�A�Ό��^�X.<D�J��0C[�-pA�7n�o]��?��W��W>�ex��������R�f����/�܅��UA}��{�󳿂��MOxJ��e�
�c�Kh<�,�e���i�h��c��Px�_q�L˞�{�#!��l޺�^� �wOz��7�~�@c^��g�K��p��/��d�ᆗ�{p��	���~�9n�ý�-8w���֛�`݅a������O��&xy�<��(�#t<�%59ġ'�'���@#q��v�K�[^Z6�������{�����+߆k��~���˿�,w����۷>�W�{�j#�]�1����s�='��l��ks�ݼ��}^���pgwZ�.8Ē�뎒$:NI~�Lo���Ŀg��T��+<���>_>��'�Ga�oΕ�U�B
�N-é�<1�����!Ĳ�ҍƿǳ�Z4�4.��>�	J�ܾ7�`1jq�b �(]�o ��Fn�'ݒ:�垝A{V������I��~ά����f�����⧇_U(%2΅4x���^g��Ȟ���)����@��ynL��S�aX��/^~�Rr������oXt�H�{���L�)6WUS�AJ��!\�[/��k�1����.��������(]1P �D�d�C�K�����T��l^���Y�s��2����8��.;�͛��k�)d��"Ԫ110D� t�
�w��?���2ln���O�]i1���M=Q�	9R�U٦�-����&(i�bSh]��T8#��!����w� ��߷������'̾�i����f�`�`�h�y�o�/~�]�Vv=��]�]��cZQu�; �
'68�[�!���J�m*�T�����f�"��M/�9oC�0T�3�7����r�b6�qzu�1��1�m��������b�ݠ�UU�tCÈ
�EF��U��L|�� �
 �����
e���z��K;�����.�-��妰�q��?+����#�b?�&_�N)�����*/Lt����OvX���Z��-r�ּ ��5(�\<�L�od�$����.զ[�5Ӂ�n^<�4h�@Q����A�:dk����񴖠�"�(@�DI�u���Lե|��X��w.����窓�p{�ň��~!��Z�K��O.��7�}	N��t���'�K&�2դ�;�}�k`�,y��c�{�ȫo�͹~�(�`��+�*�(��E���@�T�W�PTڃ}=��}��H8X05�>훸�Q��������{_'oWad�0)~�Yq6�KSJ�*/��L%E�*p����X�*��Sa�+�b�d���5��T�Up1li�9�̶�	5G�&,"�"\hw�� �� m蔢�TƆ�ѣ,�g&�DTHTD�J�_Z��b%zڱ
*�?�Ѽ`1��"!@�>R�4�:��8:֠����đ(���bw���@r�D��G0�Ɍ�X۷(U�${������ͱ&Zk��@�r2
���LKV0�X4�\:g5���ʟ6�d�a��)FqDтb�5]KN�m�Zv֯�=�Lesf��a�B��n_����y�F��Xm�:Q�=�Gr�8�=SY�0��u���׬{��s�=�W��lk�=J�f3g���i�����ܛs�I{Q��J��q?�I8iݏ���,ŕ�/�5e���	9g�s�5��x�x��c�h{��	�k��G�L\d� L���p�����KоX�ݫ税��q�%��MC�m%:B+Ǌ�+4p �����:%�M�	�����CjXJ��D�������x� �@(�yG+�tn֒�Y���ID�G���F^}k$L*ǃ��>�� �tSJ��`׃���l�%�at����%)���H[.�N#�*	���f5�4�'W�=��`f%��t^��)��M�M�(�i`]ӡS�A\ْF�Έi%,b�5
�Y1^2��275�Ez�5*g��"Y���D�8$��R�J�.�͸G]�9�\��V�<��1�A���y0�v�e'����YaM.�+D7<����(W���["7�Z1��3j��R�9������AO>��S�Oª�����A�v���k��ϏJ�Ț- �Ҋ��hw>w�1����U$����j�p /q�E!]?�O����?	��w�e�	��y�g���;��� ^<r� �~z�]�ă�{KV��c͆{�
q��N�ʒT�Rt�Q��N�Y���U� ��*fU��� �g��}L��#[s��С�&�U�x��+F:����F��"(h�Ǹp�U���?W�z��K������g��Q�p��!{`�N��@�~�U��&�0�����+-|)dr洜�@��$,"�;�
�,��A�Ҷ�4{��q�3U�K��,�^IZ7Ľ�8h����V�c��̢��3F��*�^�>�D�J��� X�A{���J�1����m�Ugy/P�����@s����J94�t�$JЎ���!])Lw
h�&"�������x��*��CEf�C�\������0�-��<���u�`�;p
.n߆;f'�bQ�kz�����~>���N<�18�;K�7��M�xh� �5�d����t`i�j�/�'�<�w�®��s�P�Q͢�(gb$êm B�7���O&n�UP�=Ci����
=�8����7եg��C]9%��<(}"A ����f�[�\��H��PN�7�a�%�j�;9EB@����X*����H���:)����Y5�@�t�++�@�s����U�����F�kޱ��z(�TZ�"	Q��	f��n��q���:��$]������UEB��B�U��hchu�-�&L˾	`�_:�I�Pe]�[5���u�U�P��⬈���yT�]K^S\� c�x��4ٶ��%S�H� J�	4lg�K��7'(�+<a��i�~�ǽ$���nn�
"�GD���`��墝(~�P��Sq:���1��t� �@����CI�w�/�=�8�	�O���(F�1�>����DzA�
��F��C�+������Cn8�7�PN@�օ8W�(d3��1~V�MT�ssC*Z��A��|���(Y��Z��J/@Tں�g���J�B�����py�Q
$���� �B "���D��rY��i��_D�d<�q�A8ҧ
������Wb��I���Y�* �'*�qb��pvzp���LV�$�L+�V����BpPh�H����-���� ��A�B.�'��AH"�F/�	������$tx��4����eӾ�U|1�[i߰���g�5����iѺ�>�X�&�~�Hy�l��v)	�0K��ˌiݴt�'���:x�m�Ո/������j��ce-kaq6�Ǻk`F�#�Ţ03�<$�`�WD��
x��q8E��[$��Z���/�f�(�Q�Y��=�C��M�壢x��^�B�$����r�x�CL�]u��L�K�s��9����+|�֐�C(�Ȉ�S�K۴I��C����ϸ�!mL&5;�Ap�!�m�h��S�������:�T�T)'�H�)�"���%rn��7%�W��`1��!��$��xU킉"�ȅ��R�|��S�Ә]5�5$ve��l3����#2j���O�k���M���ԋaf���Dd��m�d!��|Z���Qˀ�ԯd��(I�tl�`�f�H�z	��S�k�\T���E��9vVIJ�$�`Y!��-.�ATt�N	�E�0�M���2���J��@Qe��-��9�ōP�a'0���6y�?p��6�B�\�gU��׽�%��H��^b�D��W�{�O� ���b��	�A�f�#T�5���nN�a���dF	nl}r�BU	V�tcۤN"9 ���sO+0��$� �n������ݔ!(�	?u3��pu����Ad�,�P����*uɶNU!P�@�wڎ	��B���Q�T��l���5�BU��&�*i�s&Zp m�>3a�0Aq�+6ِ[p | ����]P�
����Kn��;����^�Ui"qVS��0�o:�3���m���+T��J8�K� �����C�n�8JuL���H�N��Yy��8
Wd�3� �--��!!G�'� $(ȊC7+H͚.�,��W0���ь�)�H/ې�pY	�,VD��@ZLoF,���0�:0���$��7Nؑ�C���C)|�0L� (��l��ť��;���V� ��"��J$� 0���^�ҭN&�Mt�L!H���'R4�$LF'oR6�siay]���e(}+;�����!���6�9PUL��6����V_A��3N��M���0�>�`�dN�y��u�$�?n.gr�:����P�ǸtۈpVEo�Q�b�S
1w��le\ ��X��(��*��\?sq=x����M�p�֔J��T��9P���o$N,Z({��rO���bL�q�M���TgJ�Kz�s��*�	aşV!�Wrx��@T������(�yfԼ��lD���ڶ\pj�'�K�k���4�>;��_�ҙ3�$L �;Z����A�BdmR�Ō�"��.4�F$�c�re2��#��;p��X���'�cR�ڎMI�EI�8� rO�I�YJ%e��T-�Ń�/�4H��L&�Ĵ�:.�"^�'҅~̚ ���ʍ��� �E�]���B���?��焨[&bFD��ݹHD������\�ΘUmv&����fPV�Щ�[�e�?�F�؈���w����grl���z�D �����)�N�Km.tT���l~�Z�0�h�Lܱ��� ����ҭ�].�$k�Ղ "�)q�u������{:O<��7�����4nR�J� ���������"X(��o�:1IJ������A�;�ԅ��Tc�o�-�*)k������z�d&h�����X2N��W&h�&�D�Nɘܸw"�a�q����jy�m���������ژ��,�����.tW{\i�`�QAf$�	��`9i2�R#ZpQ�mؚ���ުBk:e�R��j��̎�LȞ(�d�Z[^C�r{�ih�d�����_��<�P?�6c7K�����?�"��m����z��UH���o*�p�a%�B�k&Y���K+>�5�U9��#if�d6I: PS=/�*0IF�~j�)���}����o-�.����A� �L�~Fp��qO$��:p끬�Gm���Na��䞤�\&8�N���g�Z�Zw�@�Z�sS��o��2*�;�Sq�a3��*֏6\�i�]ۂ�v��&���jva�cI�zp}������F���0B��"����@*�9$��-YqN:�aY�*��#�վ�j��q։C��;nȈ%( �L7^aCa�8�
7g(L��_�mJ��X6�r��و�O�XP���c���&Ң�7��-��C
T*���ƥD��������.&W���xn
�����N	�����G���p�~䜷��J�8�/f3!�f�P5�������i�A�7����o��1�K�WRR�%b��'<��e5��+c�X��s�#���.Z�2c)��Yz��O�	�:�sLGPbY�%I]�a�<`�=�"�ٌ$X
��0�s4gʂ
�n�r�al�OBl\��	2� ����Rd���d��8Im#���w ��䟋���3���f�: Q�*�KO�����Z��|dC>WQ�S)���rPMQH<&��on.�a�|�y�L6~(*����h:髕��v��)z.��f��\d
1�q��BA���Y�2��DBL��ȸ�J_�&��=��~��征��h8�V����t�`�n&{p�X�x3pX#i�:.q�QU׊�/#;dB�R��H	�G�b���hc�&�֢fc�ww��L�0�v���$XlU���j�rQ�M��)H�-\�Bǋv��W=����E�\�o�$/�@@����a����.�/*,�?���c��#;,3	���"�X�4�;,�5Q-R��r"��, ��Ñ^���sBSۼ'z�H;�F��'�7m�"Q��3����6��6�@.�9�j�J��̚�UU���g�U��׭?�i���%��K/��4���(���<)�3@�)9�[��`�eB�lb�*�CC����;%L6���p�D+���4j�D���Х��:�?�O��E�f)���a�mR�s��)͸�0�Z:gaڍ|ϱtX	�4��R3�,�RfTie�Ma�M)��$���}�WM���(nla*����ҍ�ڄfU��������<�vn�~BO"�?�
��x��l@A4�2lX���Md �D�FH���s�����Q�	271t�C���fn����K���.��(��M~���ߑy�%Y���$YiG��Ԯ���?2����6j�z~��v�����Bk`�i��AͨQN`C�3��n5
\��aL@܆N��ʟw��CW��"&!m���$-���i�&K"3�n=�X�~�O�8f�G>C�X��GØ(����%�hg]�Y���R1YT���=�Ma�pm�l²�@�mC����
���c��$� J�=م�M*#���!*ӌp<����/��ß�#�T�j.e���H���pbe	~y�u�uZ0�������^���h���"���d�5<�	i5Otc�C.R<<�|ue��~�6���ε\2����sX�x��"}�~]mb@��
���4U�{��}9q�]6?��S ��D������I_��Q�Ld��KU�R��j$5�=55�o���4]��i:Z�Y)����b�DV~����h%�|�3q.�v�><,�0Xppg�ۓ!.�tb�~RW}��kL��5��߄��:�@��e`�XZ(`\:�5��d��j
����=�AZ)C��a�RF�D�	ܻ����M�t�L�3H\�nl��s���;%�2����m ���ov̵2SD�N��s��4E#��vHd{��{�Yڐ��fb���fOeJ�\j��%҇�j�F�7�y|�.�~�a���r��=�'���q�D�g�FP���O<*�ԅ�t.�	)Ι���ōaB�i�3��E�4��f��K�Ĕ���6h���M����� ^�r�>g�U��\��H�(���l���ī�pes޹v��YE�'t;��1����}�{����BU%�$:��n������I�* A\b��
�5p�5��]��O���GP��"IRj�#2Hv�(FE�-8�,z�I����A�M���)N������P"�Y��v����~YE�;������/�f˷�o�$���@Ą	��*y�g�0=�����]l;2�*�>ZVUi�U8�WE�&��˹�B��!7�s�[�Dec,(�����g�8¼u��K���];wZR:��@��D, 5=���e����f�5��Hz�˾�W�4�`Z"�W{$C
2<�*�.�y��*��B�zG�*����T$U#X *��p,���7^�^�o/]�1F�mX�/�D�*�b�ՂE�AT^�����3n�&���K�����ѓ0��g�2�r�2˃�>D��JoH����O��s�- E�oFp~�\o��Lk%�)8�p\I�ہ�&?�m�������OAkba����4\�t�G ��(vD��Fp���~�Y����밋��$1�Z�e����$rn�p�ro�l�]9%č߃@+(��
!*šV[�6 �*f�$w���F\W�3����׉���ܽ'3��7]r�#��f�i� �Xc��Qs��}�\J�i� ��*x�"��si)����w'L�_�����~7��$��U�ĥ]Ԥ����4�=Pא��	fbJY����Ϭ������\J$��:~�j�QM�TF���R����57_��H�4�|׊�qR�+��Gp7��nʥ}�m۞0X�c��`���R�	�:P�uX��� �<���R4���!��۰�i��]�kU�������2�M	�n��˾��n݀�C�C{�K��!B��M�t� �V�{g����[p�3��+�B��)�EAT��S�M�`#�2������4�Lm�MoDb�{�6όe	�Q0��	MQ���d�a����R`뽈�~��A�����0��X"�I잀��'U?�U�W�[-z�;����g��1 �$u؇�W3����~p���^M��9j�1d�I�	Mƹ�(��(
��h��~������˲��Qi��^���¥�6_%������Ð"��x��f;]��omހ���aqm��d���#M6,Ef'j��qM?bF���c�va`gpn�&\m�d�]Ո�uyVi̢�*D�wp{�o� �{=x®����"�jP"�R�~W}hhƻ;p��(V�? ?<���T0򜡃�ex�_B� 9¸�&n�8g)w�L�fv�D�QT*2��+��L��rU=e�Bb-�a��Dns�ė�mi;���x��$�r�!�O��� (%a0`kj�k8�Mܧ�O��ɦ�R Q0V�!�a���ΈWf�_����R�ƞ�5.'({x�����O��f���q�ET��@�����Rgl���2��	&��SKWࢴ������6E��i�uB���%Cc�Ph��N�0��r�K��Fp��U8�^��n���Y�������w��x�Iާ���'
�z����|;-,"ZR����R��`�8��ș1��wlÎ���au���>�q�m��ez�~�N]%�ߪ&p	��Owp��i�:G�OϿ�Z�V�xm7�TRYq�{1j��7+óCLT�L�:'Jr0���a�±N�7uX���D(4��)����J��3F�A}
�MfLbǬ2i=��G ~\��hk-��;������!���f�λ2`�J�}Bŗ�Es�(�I��"xٔ��o�t�3�	��s�P���R
s��k`����AiJ	�}N����\3�߰X?�����c�q�0=i_�-[�l@M*��3�XۛM��)qS~�D`�?�Y�/$�
�FC"|}ߙ۞������Fu�O>G�WZ�.A�rx"g����"�+����#���p��	� ��ރ�]������i��y;�.`�:������O�/��z�2,����o�ѱ`��=U����߹�����)��뭬Ru���!�b��5L=w�q�#���e�&)�9�u��01'4��!h���LL���ҋ�D}�d�Tmd�8�[ik���+n�Fy@�U%ܴ�����lHt�U��'����G��g³� a�2δ�F�n �q>�դw��;�0���v!˿��}�;����U�Ev�a�q�~��^�������8��^�k�F#*�>�����0_��"�&�=�Ɛ�k�W#���!��A|G�E�F��,s���N�7��>OeϿz�q8�r�j�9,��Wf;	�Ʒ��ހ��-8?X�m\�Knv-���̻1tR������x.��3ۆ��>������-��ɧa:����X�[��&�j������f��s�W��Wv6��ހ�޹��-�x5���Q�;�AY��O��_
�K	^O��[(���6�db ����Q��F��j���ĥT��{ZQ��f���PY8�Y�R�D�pB�]�(���K����y�V%���u��ɉy$ ������&��6�*2�(��d��gD^�;��z����TI�2�ZB?��XWӳ~=�H�Z���9F���M��'�M�c�S�B�@�tJd��ØR���ӭ�'�5L��X�ʵ3-:�������?����߁�O?�U�a�Ӄ�V�`\ST��1R�+�T�8XO���!�/���t~p�"\�6`���1�dh��&���z��fI�.U��BаB���n��r�=���g�ع��@\��6u�U�)W�
%A	޿�^����>v^�v�{���_�I��p�R�SX��жblm���bC4��ڒ\��$-��@$㦑��ˎJl��y%R�rs�����-Hfv�o�h�v�T*I���5���y���D|(�f"P�U��BĚs������)\�x��g:?��)n� ���%��&���i�{\�Ed��/&Tf��J�^�a����F͂�=�p�*���,ٳ.&�D5T �;m}�J)ƨ�0/-+�d�iN��*(m^��Fv�;�I{�i��~��h���w����&|��x��iX.�pl��.-�����(P�����8WhG�,fs�V�=��p�ع��� n�>�(����L<qmAo��U�$�빕����8lG��;sXBcc胝ͨ�ְh�]3�w�n�g���z��0��n�u{~�8֔Ru�"omo���ܾ~���S'�����\��ߺ <W�]�ЛM��7QU�:C���P�ɒ����*岚
+[��	n"�j��F��:��LB�eʈ����R� �]��Y��:������kL�!@Z����$��F��p
Lxz��x�!�OFǝī&������c"�KI��Ɉ�W��� ґPi�:U�mY%�:㉓kC%�BN!�sc��KI��O'җ�}
��!�U:��w�N�K��z���H�朙5�ݪ���Co׸cA݋���_��祐j�hg�?E�H��*����d >����*[�M
kс)ZYC�sH}��ό�����P�P�􄐥�
v�	L;]x�.޻��^�'z���cg����#lXͨ@j+�������k�3�#	p<�w�߂�o��b�����'\�����4�21�����{c8�#`����NYuT��o7�G�ކ�^��ťP����;��y�21�~�Tu`:�6�4���K1�+���S���;����pi���.�h8�\��{"kK*��@5|0��� QG+Hk���L�(��4$��%����ya�e%��&MWt&撧N����c_�mm��	�S�.���N���H�*�����H$3�:�xܡF(�1IK�f�Q���VQR���Q�5B�:�b2I��� =�1F�`#K�F��>aaꈰGϜ		۵�d�,L2�=�{�.�߇�c\]�D�����Wo"/���*�q�ψ�9c��]a�/�Eayn��`aP:O։8#���^[�L0���v��sa�Ȧ��K���=X$82Ԫ���~��v��S](�0L�A��g�+�.��준��$&�!��:m��n�{�'c��i�UD��D{�)�l���x��[T�1�:	 (�"���/·n��m| &Z����܀��t˄a�_0��z�'���g���A
�2nf���"�#j���U���l�؂�� �;p�W���l�&�~�G�|ά��yE%��Ș�l�ܳ@�2Xw��*��j8\(�ѭs��ą�g|�K���ud��TT��釠i�d�@I�R�9J���۬B6T�7\����fu[3�[IgrK�z���[m"rF�-�E�.v)C���*Պ�mxn ( ZEr��2y�2SgHq��ES���,c�@U�zd�qGD1[��d:S	k�k;���6�*u~�8f����9;p��*!���R�9���� ]\��}���䂮�+���F<��T���sQ79X!�D����~X���Y��g��L�==�h;#�-P�_���5��\ނ&�x���za���5cOS����j��A ]@)_��M�^\~���%F���� ��<���_��`w<%����U��t	�j#O��gw���یH���aq�K�X(8��[-x�����6��?ܩ����s�g-? 3��z��
��(E���.�%�.�^���_aByn�P���q\E��H�����Ô�m�"QE)�J�*�Q�K��K%.�.���4"�N�
A���~�D�Q{�|�y�߁���$s��3�(\��Hm��A�=uI��{�a�>+�̩���D�M$�%f�%��g�C6l�����LUi��c�ci2�2 a�ɾ����iV���v,^��Y;e��cm)sL�L�NjΪ}�D����J�g�6K��М��O���)f����Z߳�m�!ג+�K��5�[;�0��m��(K�5%W��9�5�#��ݝ�8��=b�2m����l���V�OK��g�ܔ�ia�d-���?��)�X���_    IEND�B`�PK
     t$v[�īd}d  }d  /   images/ef87c5cc-d843-475d-a868-97060fb00c54.png�PNG

   IHDR   d   l   ��9   gAMA  ���a   	pHYs  %  %IR$�  dIDATx����%Wu&�U��:��yr��h4��Q�H� ��MX������:/����5,�`�0 #PD('4�䜻��sN/Ǫ�wέz����mu�������|'�[A�|a(=��S�җ��o|��于��{���|-`ِk���>g�����%\ؖ����׼���hU�t���z�,���N���_����.�1_�ի�K�4q�5}��|ǥ,��K���+��K�Z� :�M(��~�	�~y�,�԰].1��l��� �2�be�� Gdq��Jyo��W��V�7����c�"����8�ek`&���t8�
?��4�_�u��2��o��l���-�meq�z���cp���㸪lz-�w_mD�lۓ�Q�%���x°��6�0�{�XA�E0�r$�I��!~q	�|�ﹲu��f����1��ʥ�""�	��FP��:y�yXn��{�y8�2��c�1��:Nut*���������b{��/��%�[�"�C`Fê��8�,�/
�}f����-������^o����c��a�hY�h��uu�rъ��G U��QQ%*(%�k�b��p��T����R��A]XG5:	!i��p+�%�9qù$��s��E�f�%~�\Qs+��,_a�Y�Bm�U�D+ep��B���iU*%����:��!�7g�bH&���+K%Bӿ��ʸm�X��F3oa*����ܿ��Q�ϙk�U������.��^O,* 3�=�I����@uR!�2�j�Gm8�Mu]��Хc�ϥp<;���:��"�]�jr�fuEb>�r/�n݈D��rI
��� �3t+iQ�f�D!i-v�he��7�pd�Fc,����nE�k)sYo@2��l!����K�i�V�VC��r��J�(��VW���x#���it�&�`fK��%%B1}m����Q��4�"0'+�p#	�.L�кm��'Q���\�Wem}'F&Q(e����r��*��Fk(�L��l1�������ι�J���Vl����l��;6"����V'���o�pi�cq�%���s��h�����`G�VQ[�jb���6���-��]$.R��x��TrQ�>�;x���B�K!s��[w} k(���Kعv�?~ _z�[��s!�ꃟ��|
��i�.���k���9�����_F4ڀ��A\��J�������~�@�F���s絸o�=��w
:z�1����;ʶ(E=���G>���.
b�����-N-��P�a������i̦p͆����>��.��?LW�{��P-N���[v���G���g���o��k�_�|7�6��r��c�Cu�����b�2H��1�7��xw�N��B�f9c���v�n������,5��:j)%Z�j�`p@�©b�S�{W�P��~�	�!��bh�v׆�]B��ʊ/�nj�5�wcra+:W��C�i��|���[H�֠��a:���V:� *Ŋ���hB�m]ؚˣ���r6�	MZ�X�K��W�ܠ��Ќ�VS��:�X~�um$;A��W���l�-u	l�݊�D6v�������.�G-�WW]��00������ih�Gڷ�N�Q �q�Zb	��&�x^滼�v(�͉N��Z0�P#rԯ8:AuȮ�a��Xdq��xm��%|�ej��bpnۺ6�~F�NH���/?�1tpv {)�K3��q!��ҏ^}�t#�1l�^���IWh�2�������N��ê������	\/�Rx������b����T�r	��B�{�'��ŎU[037�0'W(��9xz��^����믢�Ω�/sqVRYv��[���'��[��Ѓ�������D���/
�>ZCm���=GHg�8�ڜ�R�u���R�U�ǿ��
6�^��vߍDMb55�Ɠ?�����PZ-i����ԝW����|��2=��E�C����PK+��k�?���8<|�N�Xaws;~��O�w��А��G�Ɠ'_#L�	F,�y���������(����T��e��ص�
l�m=�Z��8���}'^;G���sn[V��-�o�:���g~��ϝ �0��L���ť�q~Aqn��q���/����W2��\!M��d�#�,��J���P�Q���MBPQ�C3-b��/=��B���O���cx���	���|��'��]ă�yS��'̵\#�o>�#�R9|������8�w\!�����}�O�&�-����=�׎!$��B�Hj
���;��$v_u�<�sL'�)��"���z����;?�U��?;����H���8��������\:�KS���D�s��:���EѹF�r3�aX�8.R��5�[ą�$V�w��Ũ�_���>L,N���T�'h�"o�ؖq��w,�˝�8}K�J��S�}���O K󟝝E��+��I���F��{?F����7_�tjVWWԗ���m��W��1d�yL�̢��F�!�(q1w�݊���A}þ��x�2�8d�=������ݛ�������M�KH��+������T�L
Q�ë�*�kۻ���}T���G��P*\';��p6���ø����KY�&��1�����1i�����7�#у��V��a����C�����q���d2Jy�ʢ���~ܣ��Zl�p��=#*\vο���oQ�~B�(�v����ߢ\�D�'��Q e�ܲ	/�{���ba�Sc�Γ?F�k�~P���E^��=��;%sF9࠳�U�"���r���ã�x�k�Ggk��D� a�&T��g�`xr��OdnAY��It�6^>�6�P@�aC=�2K8[�bad�k#��޲ʐ%�j�F�f����Q䜤�!dO��2y��d�V�4�:�>��6ln��@Of��f�:�/���c�����
�XQm�.~$ส�?���m����B	K�{y݇�����W<�V�|�
"�q(�'�|��I?���o���YeT>a��D�?�G�!�hD���Xhc$����'�c[�jܴ�&B�?a��)R����^������8�x�u�pa�j����IMc����".O\�o��c��7��P�?�'���tn�lm3��G B�#��)��Ȉ��V]��P��Pr�gώ��s�~DEa��w2�u6�'�+�c��7'�q]�&�LtQ[r�?3���qL�O JS,-$�ʆ]�F���Y�q�����[O�+���"|�n���?�w�t�vu�"ٌhx���E����.�fV�v�];�`�o�p`�=�-�
ܵ�f�}�(�}�mH�7cln�V|.�x�T�1Z��k6bC�Z|�w���/��s�A.�]��+��s5޽���6\�k/^:q���<撋��9<p�=���{���+�y�u蛘����j��}�Gc�6����᷿�x~��C���"��Q��9�����N�3-Ж�����O![Z@�-i�A㐒h�8�<�Rs�,}D?��c�$�+U
�
y���`ɭ�KDӄ��,��N�.ѺS6���;�6���o�L?5�~���W}��s�#l���U�('5??��7�́#d%!���܇������8.�C�����f~y�;8�<c�F<���8s�$�)�P��̠)р����H4�^����ʄȊSB%L+N%1<5����_P��46̹($(2�$�±L�?~�g��¬r@aա/���.cbv
����$;�"s�s}B��D����$�$/%�Y2����.(�` ͸jQ6(	01�'X*z�P]������]���5FĚu<_"oK���9�`�O����q�^8�NU�����C������_xg��0J$4](�\�k�<��C8}i��. �O#,J��0=p�/a2��^;SȢ>'T���gF���_�"k�157�E2���a.��Nl̗2��G�['�`Mw/�i���ӄC�7�2Oa|�'c`bS�)��&:X�Q��A�a��"��j�4@;Ȋ#
��^�Ҁ��,犔����&]����?�������]?�NGZ���S�L�V���	/�n�ƪ*��5xxq�|�G�e�K�J�^9}g��+f)� !b!��Dd�P��]��J�E��PH#}IT���gi	_}�����[��������g�zɔ�'X�QAu�2uy��^|B����~&�1*96I��w氦�%�n�O/!D�P�v��%Z�M!��|J�?�%Fd��ۂZ�VFq���z���d�d��J���z���i�՚u5�|_`~^����1X�G#c�����9&Y�p(l��Z�2,L��
9i�8i��y�<a̯�~ ,0`j��ҹs�onbL��˘!LDȈDXǰ� 4ƿE�!U�n[����hE%�ɎM���M����,�z��|
qKր1���������3J95M#�& �!*�:���z�\�$����nhۀ��� ��!S)��.��043L��P+���eDmǨ�f����^w]+IW�N����UOS'Fg&��y�Р�1���g����~���ш.X6��t���dO;�|
��F�� c^�p)�E,Vm�Մy�L�x| -�4�z�'-L^^�k�D�l����T��@f�Hbsj%B�+DE�D�h	$����ep4��R��y���Mp�Edf��\\���φ�5����O�����CQ[�G���B�O��AEuZD�a��~��G��wo��5-X߻o�:�W��=��{�6�iܴ�F��?�ޗy�k��|
}#cxr�S��3h���ן��>~md/r�o=��fG��4�u௿�E�$bh�5j�0�Z�%
9��JPX6:�@��F%3���m�� !�v�NN�-^�I�!��tp��<�kj01��	���\�����0??�ɉ��JY,�ƶM����З�'�>æ2I�ۼn�[p��%�F	3�3J�Mմ���l�x5F��0<4D�/ҺJ�󾥤B���,�rY_(��ˀ;R=�
�N�Jr�_��a���֍��5�Z\�t�7nC<Z�֦f�
���[��\j���Ok.f��M��-��O����[�}�������B����Ϙ����ks4�=k������ts��c���SL降�6N2�	aaa�v?>��UJȭ��]+V�{�Z�ajag3}(4Q
$ x�����kv�C'�܋o�H�hl$��"����w�V�����o1>>^-��Muq|��۰f���/}�(�u��RR�U�������GN����&����g12'+U�*�v���"�]G�E�ly����nR��һ���`���� ���7[�։��^���&�
��ZZA9����RfIeJ%R˳������'98��q򮦗���\�]�v#��cnn�B܋�Wr�pr���JR���8��GUYZ��d$�N	y�H������c'��tS���&�/+�9d�2�<�3��q����s8���_����ɳS�>K�}��[C�����ɹ~�3i��Q%~�.���IZ�C?�T��=#�(m��)�b�Mh���I���]���L�����j���J-O=�{��F�`?:���j����q2�ؽ�
DBQ\"�Ţ8z����t�D��"Q���6l߸�|<G� ���6K�V�
mSR!��.tut���	ZP��Y;��5~~�۹
]=��kq�lV�����vጦf��ظi;��8���21<@�*S�T��R��^HcdtF����c<#N]�l>��s����l�>"*) ϱ755i~-J�29������E;�9?;���V��/ �Єd���c�$A��okoC��x%bɝI0��^�#G^�
��3�����61\0�}����� :[�a���������'��:���M�z�o�׮C'������ï�7ܻ�f$�t����]������ܔPp��!\}�6��Goݯ��D�z������I�POGǁSG� k!���[/���;��Тb��sx{�!�O=v��{�9�x��8t�.����:�h��ID�#��F��zGg'Ӌʖ��.�43��<]�V����I�?"B�{��o��΅�S�j��X���[�<Z��M�,+��g~](���i��\�e�!~�0W�u���76k5,Ɓ?���r�\�b�����o���[�a�&H��]WߊG~�(�f'q��9�w�=�1��x�_w#N���ű!����Zj]��N�@c]Go�JH܈:����F�P���G��@�����vvoR�|��a6����.�j�����i�7��c��D[C+lYe�R����3�ӚKJ�S�ℎ)��I2 �4Wr�.Ʃ\(K�G4=*���>*���$�q��j�N�.0�>5�.����vӴ�,tLK����&hi�д��;�Ğ];��"�U&߽c��_�2����ş��r���2!/�A�[����?���*�޹S�'@���?\�0����ѱ��s����V޻d��t��У��B�{$�&�l��T�`��-��fI���"��9���s8x� �5bR�V��W]�k���t�8jdQt%ZM��]�w� N��_WW�0	E��	Ӓ� ?��_}C=j�1�t��7$(쒩��ԇ\-�ڵb�^���z$�g�����ç��'�,�H2����Z[˝����m��8@����_!�����ܠ���^]�/��a�E��ױ(�+�6�<�ɮ����S2Eq�����XZt�l��% �RR��j<���Y%�U�  C677�Wm��+�����k�+��c�H�$�*��\�[Q;a:�R�tD�w��S��7�X*R
����܏157nzE���1�$�z��zR�%���-��w��8q�$�صM�?�����}G��-ZR��m��&lM�����/x<D�]C�"��D	�с��*�	+���p}��LJ���B��������y~O�V�Ԇ,�d���T&=��W˗ɉP��>C�����6����՘D�[�v"z�j#��w���3��(�]m�x�s�pg�r�4�;� iu����Y�0���x����wǤ��"b4�cH����5��r;.�E�
d�ͽ��{?����Ǹx�⅐��O��4����CMlm�����e�Q�����R�8f2��R��$0.b�|��|)�-j��y鶘x2mY,X���2��U?Ro��I�M�%�\���=)P�-��⋅��I$./��T�Z5p�B��%G&�Mʻ>K��jUY�4a�2�t�Z �k��{\jK8F��d��or�=�l0U����9<��v�rx�d�LR8ID���O=�4����J&R����B�,b_BQF��	R�N^o�xǗ�	B4�5�k*����UW�¤�j-bo6��$F$)��D�P �qLPa���d`��Y�+�-���i� ���$/�;�b�6�宔	�b$Ky�P��Ö�Ŋ��5��Y�dm)��c��@��Ԕ�	G��M^��n��*�PL��E�� !������9���1:9������h'��w>�o>���N�8M�`a톕�:�f�N町�����,�V���nI"�AT������p���� ��مy�뷮�"�cȁF"1�$��*eL;*IE-W���)*NT�)���Q%%^<d����*TTR�1:�K�R��(�m*�Ƶ�Q��M�m��3g/�,���$Wt��6J��dQWA����q�0�J������	�lV��M-�8ra@�A-�Y�Zס\�y3]�'��	^0�p�]��c,T���(�$�a:?
`Ug7�f:�S�H��.�����K/R�j���-����05=�}�Z�H��&�PR�(#ː���S�c\@+�5�1Ei�d/A}���,��3��4%�181���ndK�������vwtv`th@3���gg�(�N@}VgK&'�11��%�	.ǟɉ�ʨ#fx���I���b�*�H2ֈ���;��#"�m�kPb0�\@F�%W�~ㄧE*��U�z��i���d��ѐ�BE���/T�,c���y�v~�L��LE_D;)�8IF��p��PP��_Fz�`�[����;Ǡ'��h@�A:[ę3}X��S���1��AHw ���U�q�q�\*��Z�#���HW�P��y�K��!�^��{�0�\�3��{o݋{�w���/���˷��E)��}�^4���D햺ȳO���^~����{n܉�?�	%j��ˁCG��S�jzgu[���""��o����=��7�`���=�6A��(���y�e>uZ��[�ۃw�t�Rc�k�p�~���j1�{�����bu��)E�R��?x�A�"i��Nl�r�+����ỏ<����8:�`�����R.�$��3��Z��ճZ�LLN�\J���$�ΨPu�i~.��\Z}�����qcg{�883T��|���AK�i
e6���|E�m9�D����*t�X����I���.�)��s�h��J�N&�x��OhAM�ɕ[6��;oӔG"��eG1<<�M�!jo	��ﻃ~'F%���^ƿ��i�'<�p�u�y��(��I,����9�U=����S�������O=O��Dᷡ.�����&��jGG���>��Q��qܰ�]�y��\�0ЬVÅ8m�8պ�Z���X�`�݈��^@�NN^�y��)�E5���MYL�I��\!�ճfb�z�]t֗02_�\�����ze룵ZȒtICs3�G\��19��L��z�ԺYj^3!e|r������Z��<Q}}�h�|�l�55�kVb���D� 	�6�MA:�Ī�Qaf1���&*g#-d.S¹�}j!�aF��XR�P��Fb3G!��F"y�D��>I^(�q�2��	�JK�221Kf	�d��F�	bx������`9��E��2�q<u�uT�p��@)��S���]W��W_F�6��h̝�,	8�U��yDB�fS��ܵ:��%U�M�1����E���%t��E��Ke3Q.�������� �z�W���?��+ʀd�Ī�e(�-�r��ţ�?�'�}A�M{�9�\��6
[gxt���_� �����,S���9j2\��c�>Fڌl*ڏ�}	Ͽq�K���*L}}��|.�?��Re��&��5T�X�P��~�!��:��tzW]�	C$�(?�{7~�N�@�����~�0S��^L�j�׎���9޶������LY,��pCg �tU6��k�
SS��"(c�_��ij��V)�<�8Ny�ˣՔ�T&ˮ�,��l/����V����DK����l��O�lSK&�j�!��J�ۦfb�<aȱ��с��B�FI���d�%.�S�����2���Br1?���M�������4k�"�N����:X�u�GY�P�h�D�5�E�1���fLg����Y!��ٙYL��1�f�V�TNZ|&�F�4݈%Jdm�#\�-L��@?#Q�]$=&�K��t�E4���I�ߣ��\0��-��@\���M}����.}�&!���E�Ԇn�'i(�$5�~b?Q(_p�5��Z��;�ྣ��>e;���S�R�f��~����ZQk�K{%����KN�Ń��UB1	FmZ��_>���!���KV`q�>�+�?z�9I[��7_e�S�6�Ò�
:����,Q�4,)X��!�2��G���(P�r%Uk-�K�S�i��i���@���f�j^w=��7y�
���^V�2m�~����z����ʋ��ZZ��Tk�:#��(��P����R쒂Tw���Qk�WKw�M�~��5�R�S�.�7��K�hY��i�n��[��=��W��������cۦ�u�U�?}}�#�,���n��Ԃ��M�׊����%A��FM_������]1�
~�S��6�f@&y0���]j�����vj�������
�5�غ��5����S�۫䯺e�e$n,D7�Z�����j,E�U��dVUsͥ�e�x�uyW�m2��l��О;p}��>�e|p��x,�".����2(b�157��ck]=�����F���!�+��{�,j6^���9��A�N3e���=u��R�p���DK:t���Im���_ܵ+��}��7)�D��޴t�{+���t�h�ZP�}1t��A�ÇP��tݢѰ:�p �~H��R�֊&�@z�²͙�x�Ԉ4F��T:�����[�/�(���X��f�A��n�v4�E�|���׿�9�u�%�p�� ��&�yd���l�<v�.��-ل�jYV&&�m��6;"���qѣ(�dJt�i�)~ϹZw.J�SE���HO[��!�p&���|K�B��]�5Y�P��My�Էs����#pea#wH��qE��јM�T�ZÎ
�@�����}�t�6#�EI��~Y��%Y)הk�R������˿���d�����
�U�r�0�8��m�莶bln��E~�G*�m����I���k(ЯH �O$υ�#��0�]Z��ZB�����4R(颥��y)X������Ӎ!l��S�/X���o���_�׵R'[�y-��Gj�&1�ir������˞46C�F�ȟ�S1cj]#�GMƖ���Lj�Iz�jk"j�E��c��)HXb3��?�C	�|T�k��F6�jK���{�͋���{����U�p��$�猳�BKU��ދ�G����I���rrP������&-0�2!�V�!,�H�i��&I$�����Qll~Z���̰�T�\f���T-�cZ�aK+���J�22��a_�sUW�Ŧ�������M���mr5�I��$��D�BJj�$���Pv�}�����������2.Ro}]�yN�I�U�OcŪv�����8��m�KG����
.Mk�^SG�AB��� ����L�kUMI��J��dI������| �:�dt�NEyY'����"a6�#0���e�2�TӪN������$��"It/��^�q�����y=� w�0�(���X�I�\hnK���:�,��� �*�֞T:g�e��$�)k�#ԇTax��W���:���t:v�~�-7�����@S��V���M!S�kKha��0>qA����%Q�ѳ�Qy���E��"�t�N�8�r!i�$ 1�*V$�n�@$�'j�Բ�-Uj�v`����u�P|x�R��*�m:;�$��\H���5�f��7��F�(���b����Y&h�<\YX����E��(9'ΣX� �,j]M��	�hU`�ey��r��B����f~��ͥ�������^³_����ػq)k#�S�� ��C��ؘЪX�p$���B��d�%�S]8ȉt�:�|�QzI���ϭS"D���
�Y�n�g��w�갫lŋ%�@L�w-�P*��5{�sU�<z+�@д�h�M(��"�����	iR��"y�E*��A��㫤"<�KsHC���2+v�+�K�w�@���D�'��Rk�}Y�r�^<��nP_�%tG���_��`Mw�NJr7^UZ����+�J�;Fj��+�,��"��D��-�/'E�dW���թ
\Np��-�4GH��r)��LS��i�Yta
�m��n����j<B`y8��E��TW|�d�i��$�֍<́��R�:�t>F�!U�D����h�X>^=ңdXVA��`����S�%|0�ޟB�B�����4��ʅ��j)�V�Y�3S���O��
W�W=5I=:=��#�,�9eL|��WK8�x�c�/#l9�0�����Z�;��X�G�uq�٬id��J� �Ai���r4 ��G*��N;"Pk�/���9^���Ig��ԹI�ʳJ�����>���D׋�5RU�|���`T�]r�B{sٜ�>7o6#Q ��R������59& ��=���ʥ5�N��`�����ڶ��#9(���z�P"�'�j}1��%Q���HSf�RR[��I_�@��l��c��/�Y���1�@o�K���Ҝ`�	1M���Rт�����ӜsS'+���GūKXz�T8d,H�l�D%���wٖI�d�Q�s̗91����}�?/`���\+��O���bc�^	�'���%A���'~ז�NB�L�0:4��L�8q[φ
 ��#9�S�,�/�4��7![)i���!Y�L!�ԙ��굼$cy)��4	�M������@���N*G�$%���������V'[��N�1�[���=7�P��RqQ�B˴�w������U�wf�; �@��~Q8~�LPIJޒ5t}��i�;/L}����&�Ə��G�++)����hM=7m��2a��n��fZ	�KʹR_�P��B����.��*����|+M��aڶ�Ɇ�J�W|�6��6����fi{������
��<�3K�-�/|�^�T�*0$��*��兎9�F[�̑G^�����쮞�e��P$��e��xIF	T����
���Ľ�b����Zu�B�DiH��jĵ{���sg117I!q0A�P���s<��Q2�W�/�+�R��3�w�؆˯W>Ti�gI���SZ����\Cn*�X�=�����Λ?��VT��OKaZJ���O�-��C�X���i��{�C��V��]�)��.�{F��=p̉��A*zp�~=�}9�"��\�҈�\,kl"�طo�F��b)�/��m���PFٔflݲi�S��R�Y������a����uL�8�vCZ^? �e�T�WH$��M��5�=�bN�s�6G�v��\���z���9!���y[�j#�mT�#�Wf���w��BH�WȀ|�U[V���&75�,�:*�
�����Mv�"��kC1�r�U���i�Ɂi�1P�Y؊��P���~������a���
&�#ΰ�4����q3V��I;l�A֣�>�Z��������Ӕ��gϽ���YԒ��y��hhn���;x���<�Bܴ�{v_I�kNN�e�e�쥷��'sڳ}z����Da���ko��ܼ��^{�X����n?���$��=��oi��ջ���G��]��&q�t��M�x��X�x]��VN���3g�`n.-�:��S��o���xY08�'�y�Ԣ�UKK7�a�PD(ij���B!��N�ZD����ڌ˺�a��H�����H4���~@q����x����Qw�����F��K	6�*��^��-Gg�e�
�q�̈́׬:�hm��x^y{���\o�S�x��O)���7���{]�yԐ]>p��ز}+#n�U�2.;�F�N;�w�#����E1����g���#G�i5�j�o|�~���5����u�Μ���a�5a�绰�ʭ����w�Ͽ�y�S���6�X�@�u�_����KXA��@�f�
�01Kٸѝ��f���Eu�W������tY Av�C\�4����)'���ĴRem���_|��tlV�t�ɒjF�!��p��ID�t��]���0&	Y,,d���^W�j{Ñ�i���U��8|�ѡ����� ����¼��K�x�}&q���6�\�d8��L��}���1uxH��T���Ip��Q$��fMͭT����`6�h�+`:�]��J��p��7dvaSӺp�5{�&gD����9�O��e���誻$d�8*����A�����4� 熱��1��M�i�&�lY���W���������M��Mϧ4�ٶi�R��,^��o��5�A��ШF�m�mڵXF���?����6΅�"I!	�����`����}����T��"Q �U�W!�����y�|�I�i���\����wt��O|��� 	���b���ʢ�H��Q<���úrrzQצ��u�t��Ν5&�אeJ%ShZ�j�nJ�Աpf)ʔgg�vɆz	"e��/pr�1T}��q�'!�}�W��f�8�l�5h���S%
T���YLS!$]!�_㴄�X!�I���R���5)��F��k]0�ɕ�\ӭz�tN��@Dz!�^Z����:�ךNf4��%قZ��hBK������17�A9�D��M}lH���/�wQLI��O�`eW���X�e�`&4?�t���$�3�*�����
%M���t�lA���}y����#!�5�4-.���P55���eE�h�mR�v�G_
6}j���ES�(9h2!.V̢�EsH"ǧ5��c�@��NDM9p|r����y�#dkq�Z���am�Mmt�$�ie76Y���2�t��;���xa1��(ܥ�$�IBV@�5�ؠ��Q��e��;��i��&�J*�-��AL�$�&�J���A�����46�q
J�T漉�kk��؈X���S�!y

�	�XR�x��2�h�f]v�6�	�)��G/m��H��X�n-݈֬7�ս~シ�K1/Y��Gran��\�.��ʦ�����̒ӧ%$��Mmz:�2H��k2({Q�$��Z0�.h��aَ�M'+���5c��Z:y]�m2D�W��*cKw�:�=�� \���K����d��ӗ�`�#K]���0�G�����e��X��4#S���")������s�.��ne>��j@ ������ڢ�?�����ځ�K������m�5���,�?귤F�7���c�r��8�3=�Y��t�l�zµT��+%�vŕX��KǚԠLbۇ`o��f�f��o/���kL%iB�&�4����s�� ���'� ~�POض-o?���75*Ā�L���9����7��CI�H��Oۣ�����g��?Lt�t��"9&\:���8n=<Ew͑M��{�T�.�X
(<zO���}WeZ^�\��B�F2�%�_�=V��+z�G��hj�Q�����R���\"� �5�j>�Pt��F���+,U}��ߖv4[�w�@4Ѻ���b�	P�kXz�L��=�pL:������n�4�|��ud�4�6���1���i�f�F�z�����=��%tMj? ��R�ݸ�E��v������my;W]�.WsW[�]����Zfg��$W�px�mo��R�βGp >;�S���㚖�_<ֲ�M����;��K�xr�x�zt������g�*`B}ǲ��"�l�SoYh&<�8�_B��j�����	00#���b�S�a|l�:;pvq���^��HP��k�ݲ9t�K[��L��%9�7Uߪ /�4���g��Y`�z-BҪ���*F`z쓟�W�R8�~�ԋ��\����&{aڿK�÷({����1;���=�����Xz,�R�]�4{EOu���+jLs �^b�wb��p��q��9-�n]ߍ`yN��ǃ94&���Ӎ��4��������-�plx	'�C���&�Rn6)��,��M����kTUs-/�����2
���߿hYK99q�K5��&@-��ꖴ�b�/
Ĕ�%���~)����gy��}�]#�u���A{٣/��1������z�_ɚv2p�O��u���㟿��&����������kW�$�kAea���E
l!J�Z[���V�+��v�ʘ�$�''võ�3�
�U
��y��O���zf�a�	�2��ݻ��?��;̈�Z��ru���6�])�H�j�_�i�c~ib���4��u}�x�\t�}~��$�wv�8&u��$����v����ޏo}�����]Mu��������מ���ch�EҼ�qK��HJ6�&���VL��Rn?+��Bf{@K[+i-�.q����u���=��!ݶ��b�:^��țǒ�-���v�f�$)�E��SOq*�d���W����TַN��9L;��]h���>�#��L��ã�L��n	��䙀��.q�����=��[��e����3%ۺzV���ٙ�b�Z���8�
�j{:��~ij�7cx$� ����F�>]��!72��
,�M�'o�Ys�Kʿlq|d��ַ���;E-{��9��K�K3�t,���* !
BH��7�z��b��W�֒��-��f�+9p��2���*�������&ym�U8�qvz�/�M�n4F���x��$ΥS��~��۟��2Nz�c&*g��M�㭣���]�ؼ~�9�lZ�^�_(�p~v�傁K{�@\�*�KR��J=�c�ŗ#�ΪZ�i{��
'�P.����(Y^���r�`�\-\�R)��.���)�'��8&0����֘Hj҂*mNNɛ�Q����Lp�>�{���d���s�ʊr���q�b� 2�0��C���C���k}B���߲/��c��(9��B�_���1�Z�v�d���1�d�T�s�#�����1�ڂ��s,�;��V���@x�b�t��ʥ�a�Pomړ�ǹ�
^�k��S7,p�/I�%�㐀.$G3�S49W�3��{���?
),�?�լ�(1���F!�B�A[���\QBy˩����:)m)�>fy��NV6��:LC��0D3+&�u�'�I.YH�q_�I���Q}�߹�s�|-���a�c��ߔU�gm/+��\e�&GKzdk6�FF��M���02g�r��?61�Ԓ��v�=�j-0m>�z��.�-f�0D�Ptt��<0-i#�/��ڨ����>�"@�m��^�%BN��$�.�e�&GG��i5�٤����M;�WbC�L��jD.��cd`b�����F�6�����D��)�8��hu��x�9�ŝ�,,�\��N&��/���ҁ1�Z�ď�P�
}�+���]��]�G���Y����6e����3ǎk��;,�A�B�dr���4�d�Mm;�iDz��Y�h^VG��*Bs���R���-ɨS��>�w]�G��O�,�'�cb}*��9Ɓ�c��v4vaK�U�;u�C���5[p��|f�<��Ggp���������V�cT߁�T���������5ZX
�G�z�Y�4��h$<Kv�qt���`�8|�_S�7\�.�=][����є��s�	�cX���h�����\��;�2D���f�=�HJMr���kE�.v�A���b�X���6\�ۦ#�Z�r\����F�+V�B�q\D��.ɧ9^N��*,My��t������c��̐�F�Оb|���\qn5���0��Z��͞�G1��,Kv/GO��]ƎUkP'O0��ذa:Ww��#�0m4�4ò��ZΜ������a0�&Hܟ��7gz��2rF�c֭_��V�l^O�Oq�>���K�s^�uB?�<�j��Fu\�W}c[����!ˣ�FbX�q�Z�F)�9�ۮN��!���KChڂ���D�_�Mk��V�6Yȥc���Ėh=.��ǆ.F���\��5�0;�A��S��nNL#Zߎ��,����Fkk+V�\���V`�R��.��Ag� ��կ����r�7�sx�p�w�������~��w/�(�!Y�{�͸^��W:]����z��X�����V3
�j����.��ܠlR-U4��7."����jH�s�X�$q��:�5��p~��X������1�c����4/^Dw�������Sغ}�&�����\ߋ]7މ�=�4M�����]������c�z��y��]͟yny�j���YՔ�(�3c�\�f<$P���
鵣Ǵ��f���r@Ot�k��xQ�^�?��lUz�]�Z�q|n�VMxYj���dM�7Kk$��(��}�2%��u�D�'��8����%�e�i����[��E�L����$Jo�\�U�;896����K���@=�1��ԩA���_yN\���k�
�*a\�s��Lb����\�_���"�G�]6N�#�b�4�M��#R-�������/�]]��8&�)��Xq
Ք��K�ӫ+^;�n[�>+=��4�ێ��柞�%��eT�X�[��jP�u�T��=�������"h�x���<��'i����}��5�*S�G����H����a�I�.M��61.AX�(��i�k�����y�{[��*�цM�@��<6�'6�\��ڄ2'9�y��E�r��*���Y�����ػ�@�"�E9�U�/�ONz�](ݖ�E㼇�`�cq�9*{I KN��-�~��ή
���Y�r�,�zh�Q�qm�6[������YJX޶aK�����V�I��*�V�݅���5��P���G�F��-�f����;�P�mu�j��v�9U��+���}�7�}��vS�,>�w����ac=�9�0�C�g)�!,�E�LT�%ז`L��\�����0���-m˚ٖrR�/�X�:/�ޙ��f)�f���ZF�_F����'�Yg(�D4����=�>
T#u�����G6����rƺ�_;�`p�Xƪ������O���	��r�4G�3sYl�hA�.��4n�}3#��:�unSMD&��\ZbS���#�~�Ώ��k�Ɵ~�q���y����gY;�c��S���ǆ�p���L�:˶�fm Of�8t�,���?c������r������ݤ���E7����!w�7D8 }S���C�}-�{V#w9�ӳ	��aW���4� '�ɳ	�8}_��w��-2�;7_��{�'Иh1�]ʣ8�Kr7�6�?��0�Ě�����8�_z�f��{5�[݆B}�I�^��\�eZ���G�Av�n����eܲm;��v#~��eD)�����ܖ���<^:��r�<��s�r���51L�����܀�0us&�pX�+��	xc�,�����ym���b㪭��?��O��lњ#��b���ï"A�H�+���§� ]m+<�`���:^>���"H"2��/���"�q������NE�0�����o�� J�Hq��PQ�j�T|����X׾R������r|F ^Z��B�L�6$�����'qy�V�Μ|-yBj��F17���V���^��D�kWa.^DO[&.Fjx��@ѩ���;q��k�&]z�0ͅ�=��ל�lӾ8t	��܅_��~��Xe�>��$?��Y�v"�+:z��N���0�ɒ-�o_H9�~P,h�������Zŝ���B�#Cصc'���O�Δ啪.�l���p��ݿ~� >y׃j��Ξ���spæ�����ȟ�v#�Y����!��X�x���y�Q�2eE-�j����-MXϨ|n&��G� ��Fa��u��%��8ƬUQ�gQ.P{�I�C..�\���HM5�PwO7yZ=�ܱu��Yʡi�r�C�u�����3������A��#���f=���c%#}��Ǥ��|��hѩ9х���BJ`*d{Y}��1�^����u稐##ػ��W���d����v �mعU�~�K8;pQ᧖$ᙷ_���룿�E�F�eFm��@��/m�u��}��c���9e�F���}�V��6`zn#�؍=���>�O"��j;�r�hY�����EUB}�F\��V|�+�������G�R@�䈷����I\���������	�����:k�l
�\��-�Q=�~�_�{�c���N�]��Or1K��xs@T�&��%G�������Ӫ{4�-�
���L�U`��j���1����%�L�:2t_���{x����TH��7��[=Xǧ���G/(�8�	A}���&�`"W����˙9|cߏ���%����/g�����ڋ�J�/���0ӶQ�����wg�3ذz-*|���q`�"ִwb���z*�Pi�y2���g\��m\��-���u��S�}UK�w_3���o�����AIȮ��NV���;�b��+��ۯ���!�n���?��8p�^8���?$�t,/� �on��={n�v��ꁗ��C�m�u���O|��ƴ����D��6C���5���V?a���W��ދ߼�n_�ۄ�q"EF���'ݷi�����J�W(��ރ���XZU�2L2>կ��R�UHy���x�M�ʬ�B��Q9��2�l�&O�<���T��6�i����y%��PZ�>q�}������ۏ�P3]A��O�������OᑗG)h6�Zd}�ں�~Z~�����.�լAn>��'O�������܁����ёsJ�Ÿ"t�|�}�Э��������W�Y��y�#�������]��%y�	���gP	W�{f�cq���?�=[߅C ����z�{������$��Ɨ��Ǥ|�ҲCt$�N�ԧ��!�Z����hs�A���s�țc���T�X�i�'p�R���ӭc��j9�_�@�A� `�������'�(��}��_��o��~�kh	��g�$y?y�X$�b��yWm�
҂z�	��(���t�/�?����a3�no}�vB#z��׾��]��q�/�o�:.�*)����lZq���7Q��bmK'���R���c��J�ʃ����ړ�qXǹ~��Ua|�+���V�a�	���<3�<�]��z�ů�'|�;��ܔ�Pb!Ao'�<\���p��NA�9l�Lr�� i�M��uupR)��k��#d0�e\�-8���W��.���
�oO(�<�����o��m�GΓȳ��(�}��/�r><}��W��]\�?����M-5�غ33�f���4D�\�j5y�W�z7��nك7O�Ã����ۏ�}�pӦ�hkh�-Ͳ_š#o���#������O�y?��ݯb׆uض~'{��X��Fӆ`�FO��"V��VF�(�U*�G�� ��m����x������I�v�ܶu3V�իc�kѵ���vL�L���_�Ƶ[�G�m��oEi���$�	���u�@�j�pٹN��,���n@c�ZLOM�.��S޷�6<��9�$,ܱ~-��t�u�]ь�.aCov0�	`*WĖ�^L^�C[�Z6�L�)��QM�q���'C�ɢ�~�6[�R������DH��:[;�Y8�6~��wcmc�nڍ�=�nش�Z���QЇ�A�̒��h�m���L��6�݋�ރ��y�'�c��[,�M�O�!�Ok��Rl�Ʀ���֡������ٸ����ů�Oܴ}+��t�]�d�m��5:a��Zݽ��G/��fZ�]�Ş>���̺��j�V����!�x���,/Y&�׶����?}�Yr����ꔃ��?C���-�>�	�&�aMZ��19�(��DKf+(�\F�I�]��-im��x��Y71�lb�:8r�pD-��~-x\[[A�XI*G�pq���@����~
���`}gZk[��A�fm9�UL]��N*����"�H_�~c�s�.N��������ӣ3�h��^.�˲�~���b�׀�|�S�w�4�j��ڋ���hm���ǵ�yf6'tM�_�ͫ6(DI\s��n�'ߠ�.��\<���D�"��x'9(���_G(�����{�T���9$�Z�ܹ-�98�Q��d��`W�p�zW ����WT0� 5erv��1���vpR�[�b��,v�߂�+����3����^.j�T��H$jQC��{��h'5���֧��p��>�ݗ��u�˼w @㝛o��ڃ����3����V�_�n���:H��$��9$g��d�7���u��m]U�{ZlI��/��4ξ8���I�
I;P(SZZZZ��ӴC��2e���3�2a(��!��Y�8m�4ISgu���۱�}�l˖,˖�{����M��{��ܳ~�;��/^"��q+v�_ٰ[6nA>y���I	����9K�I:���E҉�|�R�75#��E&���t@�Sʶ������G��{ �ե�>�zo�݁�@�M}�:���񳍏`��B�Rd�`p�,���I_�����	;&H�Z/�����OqJc'HUѕ�£؜���i��2�a�T����Q>g>�[�)�tæ/ F�ߛ�Ei�$uA�,ny[�dF��7@����>!#c�|ﺵXB��!)^�f������Ңqӝ��ʕ����#�s��0� �������b̢��*-E{{�Ћ��X����Yt�ǅG�l�\ܪo�kNc��rA2�ѕ�"B��|��	T�
a�҃�7:��H-��	��R3�C�:�΋G0/� �ω`|� ^;�_��јg��8���Q;�f�=8'�����d0砮��S�gd#��A#��]�� ���p������lᲕ���u�RD�mn>�si�k�Ԡ��Ӂ� ��<"��͆:,-���6o �Ǚ�G����()���|A�ѩ�9����2K}����lo�����%K���hk�X�����*���u�h�E��,��=��t�IgI�L��q�<��������=������t�Nl!:H�d �ͪ�(��qL�D�B+���!�[m��U|p�!i��xd�>	#Í�:�����&�k�#�-.���M�tw{�[�J@�ɿk�:�#ү!�t������l\kkBin&��ط�F��e|SN�ᫎFE߃d�jji���s��dȑ���}ȅ������� d��Oa����kp[�=��`�1ic����A�����7$����d�����<����p &�ϐ�|��2��c���$t���2�5DB�kM�?8��vR˥2���+��1GÜ=���xf�Sp�2kXԻN�8�-"�C����h����w�ZaC�Dvn D���v�N��N�#�'��"E�!�
~��'�������M=�����.��&��J��d��+Ld�"1r���cd[�p�p��2����x��\k��qm����Hjj|S�ݸ���f����%��э��X�LJVߨ���9����^ũ5�����{�¹H5�Hǧ-��(yx�>� j�l62A4<��l����%ݼc��פOQ c,�bu3Ej��Ps�Y����!S��ɵc�0�ߊb�i�+��p���D�|Sf�����'�@e
g(�ڪ=�B�M���q�r�dÁ���ş�����t"'Q��I[��,n�㊡=>�j
���}�����B�ψ}/|�yT�:�d�~�8.�0*m7�F����@}� ��!��/��1���>�ߍE�d�M�p�3�ە�Y�x��S�e̓x��]��f�e��\�9G6��J��N^��Y�9�<1E�|�\��-W�(� N':�v�����4CQ�3�/�'���;$r���x陙�&Ł�8��4:=����g�ō	EϪ���p$����s�Hҥr"P��{e
��q�������G?zR�9��
��I:����g�㡭�ӧ�8ԉ�,/���a��W�G��'�Nbӆ�b5y�!�zn]�Q��9t�-��ہ�Kg�g^�����T��G�c0�FFEr������^�9v�6�FVv߇?��+d�2P[S��+�!)����)(.Bь��0���1��^RDv��E�����w�~t�)v��ŉvӎJO�\����^�g.���%��9������v	��0�����<CW�i]K����pU+ә�Ț���E8�^7ޯ?��7��G(����+hki&��Ӈ�!�������g`��$�
�Q�����~�>�a�u�k�S��Ұz�z�ͤ�?��l������T/-��=E�m�j������n'y^�X�zz��<�o��;%�>��ީ~���x���������݉@_���٫*�Y.��� �E�9y^k}�ś��t���"�Z;�}{z.Љ�d�?C�����N/^������H3���[8K���j�QL�$�=BQ��M�M�n�� $�����+m� 9�.����ӈw�Z2���å�N���c��P�T���0x�����[���B���_���*�����ϖ�ۨ(���N؅���'+��hӭ�¿u���_�}V������ 9Y� Us��^|�t�W^�0hW�WR�}�!���?a��ش|��#�i��9t�'�
���n�蹅���K�D�F����t�R��z�am�2��|Wv]T4�q��$��o�ތ���6&���K6�?«�����2C��N��VQ�{��L"T&�z]��j��lR���c�p��xf���'�����]��9�MS�I�h�E˥.��H5��c��x�67�\�KA��B�4:�A4�V��������d���t�����2���ن�wje�0�Z��N�e�	�ǉ��t�+�᩹���-���j�I!����-C�bCL:!�iy�ZZ).w�*���/��\2�7xp���W��R&��@lӈ
U�PvE�ƒE��������&��\��J��y��0ݓaRR�c"J����
3�(G_��5B�������JSLp����CF%� ĬN��^�!�J���V�����b�s:���f���2O>�u����a��M���Lp����vu3Y��f�"0��EE���ʛ�g,���h�B���T�t;���D�d�&N�ڻ�����,���54�����+�t5�n�0�B��	���©4����T���fD�ʝ��&)������-B����6�ϗ�åB��df#��J3rɶ� ���C��%Ver�o�F*|��)ך�5LC=v�6J�&��i�/�p����n��iX�k�0V��v��0R�� 4�v�k�@�sɘS$Rp�6`��L}��;h�)*V;��h9v�F5�$�A��;����#!dQa#5�!P��Q�@փk+R��f����N+��@�75��1?��w�R�Q�ۊ ���}�+���GE«�9�?�����z���A-�-���J
�'��i+��%\}'�m��Ҩ�5^�Pn����h�Vئ@е3�Z�VK��ʚI����܂C�t�s�+���+�N��F�[8���I��NQD_�R��p��co�E�g ۝��y���ݢ�e�$E��@5 j�#d���`�,�2��LxTB�mZj���$�������oL���@�x0`Z�oM�ѵ��	yN,��M��cKA+껰V��S�	B�.e0�i�U} �_�z8ug��$�sl ��⥜"��*X�+�q~�nr�2�����8���M�x~�
z�:��!4Dwxﻁ����)[\Ԅ��X�n�Yᦪ�Y��哛���#�}�)�r��BK��\Z��ٚ2����k
��Q�)x`C��M���r[��BN��ba.24r$��X�~Z�l)65U���&8���1Ik���՘�3C1��*NE�Iv�Wc�1
�ʬ�(�g"	��M���Zx��kiqEV�A�й�~4��c&�i�(X��$�=Sy<<ʛ'�	�-�)��9M]sA<����$�p��U^כn�<�q�'�����Yݲ�]�e�&�P�l�%�	)М�6�
�z�d3Mm]�Ko��wI�ֶC�'�!-\W������.ڰ����ڌ�� �P�nڃ�!�By%n�R    IEND�B`�PK
     t$v[t���?  �?  /   images/e2e2c934-b375-45fc-834c-534243cbf361.png�PNG

   IHDR  L  	   A_*   	pHYs  \F  \F�CA  ?5IDATx���y������ϯ�i��qa�x�DI<��D��x<j�5�`��db&;;�&3�f�8��a�hČ��Q'8:*���!�A����~[U��B74PU���������#������6    �ݼ�曓�,�'���<�4dȐ�`+&    ��K�v��`+	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`�Y?��^Ql<��vd��Y{F����w��/ʳ��E�|V,>��&��;k     �����wD��w�b��E���?���������ҏK?�
_˛{-�5������u�o     PӒ&s&~wX1o�~���J��l��~����;�<�k�;,����s:     �II���=���E�,��J>��l��/ߛ3O�y�ߜ������      jNr�d���}��?d��k�,bT4fOϙ���{��?f     PS�
&3���y^���KpuN�o1�ƿ��1��_�     �f$Lf��7�<�5��K��H��>1�8�x{�     @�H"�L�xeS䅻��������s��g^Zz{C @ɧ�AQ��������TvX,   �:�D0�=��E��>/��;o������\ T����-��'Q��~�X�O���1=    �P���w\٫�;�C���б�һ� ؉�i1 ��c��!�4P��~��t|1`��ߐhl<6  ���5�[��+�������r������l�KK���IGs�3
���������>��_^ ��/���Ē6��MS��g?	 �:�o�u�std�����ڏ�~�lwuL���U������� ;X�|�b<Q��G�g�X\:�g    ԩ�&�ĉ��v���Ǉ`��?�F^�%{m�����.�^��p��   ��������}
�跳>?˳� �@�����X2d�'E[��}"V    P����رo^^�k'ɣ��A�Nȧ�AQ�� �c����gg�cm    ���&y�V�y�$�,�i�[ HK�||,��e ��&.�$V��ã=    ؤ�&Y�3ߩ� � �����1���KG�M\�->_β(    ���IG�Ya'.� �[�B��<*�m���[���U�   `��:� @=�_��#��Jo7�ј��e��7   �NL ���Gk�qo�m�M\�~vx|+    �4� jL�B�y���������a��    �K �!��qA��O�����?Y\�?    �L0��?_�<�!�(|�B%�\�7    [E0���tv�"e�e����K��D��7[z��7�E1�d���  �v$� P����Ȳ�"e}�߱��l�s�=`��#�ֵu됍��Q(   v$� ���^�߾�F��9x��ح_�   �I0ل�=���!�G�]v�b{[�-����+�     P��i���>=z��������b�+���3�     P_�we��G�<'z�6h������"/vĲ7^     �~&��u��>4��_��~*V����X�"     �� ���e�!��/k��=0��x.     �� ���*�wVS�-�D     j�`R���٥�M]�     �n�	     �<�     H�`     $O0     �'�      �L6����-��|SSS���/     ��#�lB9�l�X,     P�      y�	     �<�     H�`     $O0�@�P��}�n�|�x�g�755= �X��]    ��&Ȳ,�������c��ˈ HDG�ϯ    �#�     H�`     $O0     �'�      �L��b��/v�~     ��	&%kWE^숬�Щ��W/     �~&ey�ߞ�{�۩�Wϛ     @�L޵�7�̓��Ȳ��׶x^��73     ��!��k��?�;/?�9�C��X�"�?�@eF
     P?��Y:cj�[�8��Sѣe��!�c�~�^z�M     ��"�l`�[��M}Dc�~�w����ߎb��.��Q�[[['v�w�����.     �{�e09��S�,���7u��g��V�ѶtA��F�,�Ύn���     @���`r��g7�^���Y�}=��J���Q     �-��`���z��5k��eٞ     �E5LZ[[��^�Ȳ�      �J5LZ[[�eY�O���     `�d0imm�j����B      l��&�ƍ�v��o     ���T0immb	     ��j&��7nt��7     @7��`2nܸ?��|B�e]ڳ$�c�*��/      tJM��[�,ۣ��]�;���|     �s�>��;�����[���m�3-�ɟ     tN���P(\����tu�yY���P�|     ��Uu0;vlyfɟl����+�bP���f�_     @���`R(.��1^}s�N	&�-����      �_��1c�����m]Nk�̷㸃����r�Z�<�Y�6     ��W��������Ka[Ǚ�tu��֒8h�n�#=>��      jC����k��~57أ_
;f�Iy�r�     jCU�Q�F���1�5ޛ�WƓ���<$��uŘ����&     @m��`��ܼO�Ow����sc���ư-�=���*ˀ     ��*�ICC���=fG1����o�ғ�A}�c{x����̜     @m��`R2x{�r��_���u��>�o��[,�,��j�w     �E�L�ۺY�hr���3>�w|r�A�e۶��5�⟞����4     ��T���[�/�PyFȿ<7;^�ݢ8���c��ty���b��o�#/��a     ��U��$��i�4s���~�˕幎�w`����^=6�̼��*���ߘKV�     ��Ue0��f�[Z9
YC���=���~}zF�r<�#V�]����/ZKV�     P_��)�y%��      �	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�@�1cF��G?�ٳgGGG���m��b�رq�)��.��     �L��-X� Ə˖-��3o��fL�>=~���	'�g�qFz�    �*�j��O?ݥX�~k׮��~�r���q��Wf��g�     �D0�����-�̙3�2�䦛n�Q�FU��G�B!     �`5�S��T��~�����[�[�n]<���c���q�i�Ÿq�b���    P��qMMMq������_�%�%�=O�y�Nm��[o��7�\�P��c���:9��c���!     �`u�w��q���w��E��C=<�@��������b1�z�ʱ��Gkkke��=��3     �`	*G�/|����^��N�4iR�Y�f�ϖc˄	*ǁX	'cƌ�^�z    @��R0imm=��2&˲cK��y>��~� jV9z��K.�${���O3f��Գ��R>n���=zt�u�Y1|��     �5[&W^yeaڴig�y~y�eG��Z�� �CKKK�y晕�Y'�'O�U�Vm���˗�}��W9ޛur��'Gsss     Ԃ��SO=��iӦ�Rz{�8�xo�ɟ�ٟţ�>?�p���K�z��Y'��'�tRe��C=4     �ه������y�_�9�d���g����_��I�#�<+V���+W�\?����/�8�9�     �FŐQ�F5���ܖe��]��\q��Y'�?�x%���⋝z�7��M����y|��ߏ�;.     �͆�$kii��X|�^�zEkkk�={v%����?�e˖m��<�+�M    �} ��7�/K/_�-(�������3×544    @5ZLƎ{D��;���͋|0~�����o����
�B�s�9    P�*���+�,�����ށMhoo�)S�T��z��g+�K��C������     ըH~��_}&˲�>s�έ�$)�Q��;�t�ٖ��=zt�u�Y1|��     �f�`���eP���V�MRޠ��瞫l��Y�e�;��q�	'DϞ=    �4�;v����$m֬Y���W��Z�ti��0`@�3&�<��2dH     ԚƆ��1]�/ȁ��r������J(�:uj��}o6I9�|�ӟ�ҟ%    P��<?6�����kq�����ɓcժU]zv�Сq�i�Ÿq���    P����,��],�	&Ĝ9s�X,n�����W��^�z�����~z�1"     �My�w@[�bE\x�1o޼n����&9��c�]v	    �z՘e���6eʔn�%�0r�'V�&9��     ��@�ʳI�8�8�S�w��    ��j�ȑ#cРA[5�d��w����ʲ[���    R%�@�+/�u�wtz�������L�c�=6�1     �oJ�0 ��o     [G0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&�-\�0�y�X�x�V=?p��9rd���'     ��`l�����K.��˗o�8C��;�#���     �F06�n��XR��oƝw��^zi     T�ج9s�t�X3g�    �j$� ���y��U,    �	&     @���ƍ�]v�f������_    �Z � ]֣G��u�]7{Oc�?^    ���o4    ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	ԉU�VŒ%Kb�=��,�    ��L��u�]q�7ƺu�b�}��뮻.�     t�`5�׿�u�p���y��Y�fŵ�^7�|s     �9�	Ը�^zi},y��	&t��k׮��ܜ9s�����s,    �Z!�@�kkk���]�˴i�*    @�L     ��	&P㚛��V��w    �"�@�;�â��1��ۣ�s�1    P��qÆ��|�;q����;�ըW�^q�y�Ÿq�    �	&PN:�ʱ|����<�M�>}���!     ��`u���%     �:�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O062��X�hQ�}Ϟ=c�������     �W�	��ڵk�+��������5�\#F�    �z$� ��y�Œ�ķ����4i��&    @]L��^|���V^�k�ܹ1lذ     �7�	�^[[�6]    �U�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     P�����+ؾ�\0    �jU��#�`{+&      �	     �<�     H�`     $O0�khhئ�     �J0�>|xL�:u�ך��c�С    P�`�/~�`2cƌ��ݻw\y����     �H0��u�]c	1}��X�hQ�\Ϟ=�������    @�L��ѣG�1"     R"�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @��y�ǓO>��̜93֬Yө��o߾��~��ȑ#c�����а~�_����#��+����N���wjܦ���s�=㤓N���??z��     �J0�:���W]uU%ll�r�={v����[o�5����e�]���b���[5f[[[̚5+n���ʸ?��c��    P��7�t�Vǒ͝;7.���ѣG,_��[�,�x��+��n�B�     �F0��p�¸뮻�u��r^�]ҫ�^~��xꩧbԨQ    Pm�qS�N���";��O?-�     UI0�W�a��,����|��/���k��/������k���?���f�1eʔ��ۂ    �	&P���cC�`r�%�ti���;����M^;�s��_�z444tz�9s�lL6�]    ��`T�w�yq��V6}�]w�5.��.�    �Z#� ������C�F�=    ��	&�z奼6T(    ��	&     @�      y�	 Uo���Wf��>�>�ڶ�X���y   v�<L ��mKz�)����b��پ�-֬�{  �'���У���Y� �OG���I�Ʀ����y   v�����<`us�9��Ӿ��j���}��  `�$     �`      �      &�z�{o��n�^�    ��	&�zGydL�<��:�     �w�	�^kkk̝;7��(�1v��8���    ��	&�zY��W��ո��+?
�     H�`lD(    R#�      �L������s��[�l{�G��    T�j�'?��J Y�x��s��zj�l\pA<���f͚�����q�y�    @5L�ƕg���?�c�v�m�p��J@9��sw�׊�Ç�]w��&M������    �j$�@:th\}��Qm��k���    P�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     ժP�B����v��	     T�����M�;�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @��˖-���;�~��8��c���Q/^�<�H���ǉ'��
    �j$�@�[�zu\x�������>�gώ/}�K;�{-Z�(>���Ƃ*?�~��q�wİa�    ��&P�L��>����;.�(
�B�,�/�Œ�+VT���W_     �F0�7���έZ���LW�~�bg�;wn��    T�j\��Q+j�    iL     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L��eY������3�Z�j�s    P��q}�����'�|2�>����,Y/���F�w�}�     �F�	Ը�~���<����ҥK�s��\���s�}�Y�f�UW]��&���    �	&P�>��QG�>��Η���[��.�(N;��$ּy����o����g��ѱ�����hmm    �j$�@��W��?��&�-�?~\s�5q�]wU����?����l�TB�<�֭����=��hii	    �j$�@8蠃����v\}��zϜ9s���f|���}-?��m��e˖ń	�{�5k�l��}�K_
    �j%�@�8��Sc���q�7nr��{^}�ո�����D%�>�K��r����\9�﷤<�����F�=    �Z	&PG.���1bD\w�u���/o��g�y�����'��Ǐ���o���,��'Vf��7�ߒ���8��+q�W�^    P��3���{�L�2%n�馘9s��[,cҤI��c��g>�8��bȐ!�����C=����.���766Vf��7�8p`     ����ȑ#��c��ɓ'�-��o��և�[ެ�'?�Ie?����/�@���G[[�?�P(�)��R٫d��    P��c�1f̘8�����[o�u��D�<�3fT��ʲ�f��Tb    @-L �e��<��J<)�")�CR^jk[q�q饗�     �L0������=�β^����3�	��.� !���� fť�d-��(-�h圥�ǶDT��Cת�T��9�Ğ��p"��B�.nB�T@��p5W��o߽KN���f������{��;1����<����>���Ї>T�k�ܹ�v��m���������#�    �V �@�����s���:����?���)9ꨣ꟫�    Z�`�c�=��/�s�=7n���뮻b�����K/E___�=:&O�\�d���1eʔ     hE�	�Ǐ��|�#�     G�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0��v�����Q�FE�R	    �V'� �lٲX�pa,^�8{�X�~}�x-���q��������P    ��$�@�-Z�^{m,]�t���j<�������7&M�g�yf�v�i1lذ     h�	d��&ɕW^��w�6}���~����r�Yg�駟.�     -��(�WSJ��Z(��7�<����g�����1w���'�	    ���SJ.��hIEQ�w����w��ܩ�^�r�p    ��ڐ\O�`-�6�ȭ��W_}u<��#�LWWW�|����އ���W��U���7�1�\w�uq�9�Dwww���    h�!��O)@K��Q�p���%˗/�gj�����SN9e�7Dj�M����ƽ�����Y�bE\z��9Nj��9s�p    4�Z0�=�tf M��&ȗ�����;t�ĉ�2lT*�8餓�ˢE�⪫�z���k��K.�����/})�8B�    [{[[ۂj�ڟRj�i�b��g��>��[^[%�3t�q�W_~�����������׆�:��bΜ9��W     U{oo����*�O�)�_�>.�����%���?������~���__~��_���<��������_\�4�vX     4��Z��!�@Ӻ�k��~��{�w=�����P(��	'�P_js���Ƀ>��������.����!�     M=�̟?��������Tjo�\��[=7a�%��v�N%�{�{�S_���ַ���x�裏��V���    �h^?y�g���mJiT Mc�ҥ�z��-�|��q�W��ѣ�{9���o�\~����I6W�K0    �?����?:s��O����4�|�ɭ?���5�lTr볟�l�r�-�r��M��&�    hD��$,X���f͚�R�@S�ɵ5x`�Z4�=�`�f͚     hD������ݽ���o�hJ�rΒ�ho��?/QE     4����?�WgΜ�XJ�;�{ M窫��h�|��     h�otb��?>�S�loo�FJ�_��M��lm�u     ����N�t�M,Wg̘1�J���)�Y�     ��p�7��\�5{��O�[�nZJ�r�Т(&�ۣv��5��     `�P0�h޼y����ז]�����r�_     `lS0��ĉ#���zhժU�aÆ     h�	���s�FWWא=���D,Y�$     ��`     dO0�&W�T���`��p`C9D    ��L�����[�s�=cԨQ1���o���8    Јhr'�pBL�6-n���~ggg\t�E1�>�������>�l}̘1q��    @#L��Ն���׾�/�U�VőG���P[��^{ŏ~�����[�Z��{���7n\     4"�Z@mn�c�=6MWWW|��    �F'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {������{��{�1v��lo��j56�Uc�Kk�����g^.��     h����J��=���IcG�����W�?��Z��x�O/     ��2�EQM)��g��>��	1���bܨ����G�}|}y왗�ǋ�Ǌ�     м2���������=����W��gʞ]��ǂ�=�<��z     h>L���˕Je��{��w�ON?�Mv�J%E��o��cG��_?U�     �NC�����v�����5�c��������-���â	     4��&EQ<���9bX{|�}��X��a����G���x      ͣ!���G��ҥK�/7��{��ĸ�4כ���I�Њ⑕/     �2�̙3������r�C;�~O�~�1R��>vJ|e���     M�!��k�N
&3��7�^��G0!�z�      _���������.O)ۑ�L�0:�?*۴C&
&     �$6���'?yn֬Y?+7Oۑ����
���Ǝ��^X     @ck�`RS�T�Q���'����wL     �	4t0�������r����|�n�b���*�'t�_W     ��:��T��RJw�K۶~vϮ�1����-     �����d���̚5�r����Q�;b(��    ��i�`R�aÆ�>�������am�J��C�|     ``�"�,\�pMww��)7�ˈ�~.UR�����     ��4E0��?��===�U��)�a     ��4M0�����yOO���j�{)%�      ;ES����������V���R      ;��IM�M�3f���v}���      �MLjn����Ϟ=��u��}��=/�T	     ��д��f޼y��էzzz�)�����     ���:�l��ۻ�\����sR�Z��r�T��     ��d��������rʄ���٣�w|��?2      �DK��n��g�����u���m�|�}X���h�{վ�����e[����(�6v���Α��3     �-Lv��c9!*����bՒ��+/��*���7\����E���	     �4�������[��s��1qڙ����ņ�V     �:�׌�x�ƒ�R{G�ylO���E�?     �� ��f�w3���G���o{g�~��      Z�`RJ�J��_?|�~�	     ���T6""�_�6|d      �C0�نX�]�     M0     �'�      �L     ��	&     @���T��X�z�����cĈ�:::֗�@&:��    ��`���(b͚5[���l�`2u�ԗ�Շ �}��    v�     Ȟ`     dO0     �'�      �L6�R�O𾹎��      Z�`��J��ƍ      �	     �=�     Ȟ`     dO0     �'����r     ��	&��+���u     ���T���+/��ac����{*     ��!����G��SO}���7��5O�>     ��!�����7FL:(F�3�/*�Xu�Ϣ��      Z�`�QQ�3��1��=����69ݿ~M���X��      Z�`�:��LjQ�ewǈIFǨ�Q��^x:�>�HT�^	     ��&[�꟟��z.  xs�   h	�	  ۭ��-=�   �f'� ��*������_�����L��t������_�{�h����˗   �`@�K�����fAqw,�ߋM�����ѿ��tt�]@(8�#�  � L �����bI���_.��D���o���Ԙ    l� �L��%����q��������k.
    L0�&��և�:�ܜ)Fmv���ܨ��dP#   ��L �I���Œ�Qn�P.]���O�=�^񩔢    �)� �X�w���(��rw�f�ϋ%1��-�]�V��   �7����-R1���aP ���Q��X�J�S��Ǧ'��ƨh/��Yij�    lUK�"�u����SZ 0�1���8)����G��MOƿ.(�,n��iZ�    �������K��{~�x. `������]1-��r�m���Y1:���M����u   �&Z:�D%-��g2�� �tl,+�ɑ�r��ӧFG�/�ķ���_.w�#��    hQ-L��q��]يib�� Y:&���r�M��dL/�Nߦ����/K�45�   ������I�aI��'G�0 `�c��bI�\n�~��7�1Q�_�[�   @j�`RI麢(=�E<>��/��� �������Ҙո��}�N�后sIf*��Qm;#  Z��#>y�:�j������Y�����˃A���d������| R���6�#��K �ڼ#Ž1=6���D*�m��_$���W��y �V�x�%��(��ɱS>��#�����$͙S}�G�]Z��/�E�����oۄ� �����ruj�$��\���E_��L���   ТZ>��L9�?\>�+�>EL��L꙳6 �����P�z(    �B��64ֲ������W[��KVĵ����    @�"��t�E\>�YEQܒ"���(����vç     h*���f�G�]zZ��?FJ�w潋��E��'�3g}      M%�`R��s�c�.}Oq}��Νs�����#/8h��     @��.��L��7�>���~��ξ��R|�<4l;o�hJ�?N����     д�&5�|�sk�Յ�\w���T��*���m���jW�����S�;��      �Z��d�?���,W,���??~��'Eqr��H�ۋH��s���K�,E������>���     h���^{S��-     @F      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`    �PQ�SJ��x* ����}�
Y�    IEND�B`�PK
     t$v[e���  �  /   images/6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png�PNG

   IHDR   d   0   ��ߵ   	pHYs  \F  \F�CA  �IDATx��{LGǿ��w��AN+Py\0!���hB������jL�6��h������Ķ�i�O����i+MK�6��FKm5)6& ����X�x���3{�	��=�N:������w�7��E'dnݺ5��9���T߾@�I��ڕ������D����	�\���`pA.H��I0��\�����O�&p.� 3�`,(Z'��Duz �v����%HFk0��G�s
49�&�6O�����LJ{f�낈4w�C٠iڛ�o��nĈ�	������W
����,���������x^^.T5�����;&Ռ6�",H�&����$�y��f
rV�oP<��b�D���^�Iϫ��?5��������)�#G��X��.UB�%�~�+�S/�Xh´��R�>��Ȳ��E���"�H%Z潷D7b���3#��P�A�[��}�w���L��R�$�:��ϜGEަ�����9^Mo�#�{ox��*!�Z��l�BOk��p���\HNIa"%@GD�#���6�(P����@��59�꼼�:1�K7�����Y|
oF�&�-��]��J�G��Oh�մxz)#b��>�������������ے	�]��wpbd����F�����?H,����?zoch܁��Q�>c)I�.��(��μ�}u[�}�����T�yj%�C{?/^��f������L�#�ʩ�YF�DBK|p�"��斖���������b�	�Z$����|jkk������!�.$k7L&�����ގ��.444$`o��#"A�ks:����@__233��א��$���鍺�n�#|�7pZ)�Q/kԙ(gϞEii)o�ç�Z5�����!����v���.N�|@�����a�?::�'N�b������N�yͅ�Ҩi����>W�~�F+U"�!�E#++K_�ĺ��,����	�j��(�`Â���F�c������E�����t�jCX&���\��{Y��.56��F}��K?����7�����ڵk��ƍ�	=�ߩ������l�cǐ����%|>+z���^��� V�^=o��:L���~ϡ�$����Ass�>u��ۋ]�v�� �}�-��(ӒN�4Ҭ�X�V466"99Y�h�b��ˢ�,X�������dJ���|}{��ˉ� .��gKs�?U�C�]B�c��]��hL�px�^4�N�<�Ʌ��e;��G�r���C}�1�F��hLVp�Ejmm��-������%w��(/\�����@]k,"�)�:+�Nё�i��#Q/��s�9,'`x�^C�|��:�C3)=g��&-�[6c̻�4j*-a"C� �9�/f�
Ց�Y!��<f�@_�D��2�&���^J��!�����P���]�� D�P4U?��<9QN�p�(nTVV"xߊY/�_��!l)�p\��['��̾�7������7m�2`0!�P�{&G3�(²W[��]m�)�#}l��wLL�®_���To=MK�iĘ�����>�����9BުU�<)�twq�`|�7�4o�k�9�:��a�FR��:�F�.�}k��oDF�3�L}�N�I��Ĥ��Yw#��N�q��V�V��T"� K�9��$\���`pA.HdL���{��X��aT��Z�    IEND�B`�PK
     t$v[�;� � /   images/31959ea2-aec5-42cb-a646-ec7cb3b6e41e.png�PNG

   IHDR  �  J   yp66   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���|ս����ٕd�w\ c���!���)��dUK)���8��I��.K�!=7�RoB
$�$�$�1�m���Μ��Jbp��ڝ����~��n�hV����j�9��r��Z                 ��                 "��;                 (�賄R2&Q(q�-�!�t:�}�>{�Sv��P��*G�&K\�}x�><�f/&�d|�o3��){�k���X���=�C�ً�>��{]���
e�db�J̜3D���n��2�o|��=هg�9���9�9͑�q�s�>4;͜�ҜcMH�8{�{�^�      �@G�@��pdΨYW?i{Qm_ʾ��=����]�B��0'/����d�g��Ϸ�$��z(��$c��/L����}���u������ε��{�����d�����dR�N�����5���WC�w���:���xE��J(�NH������ÐTN����w��*���q�o���C�!eo/�s��|M~�������Y�đ�{���      �`(�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�"G)5h��+-c���y�24��8D\�Jaޠ��}{�C<ߓ�];�m��eS�VY�k�lص���               �<�qe���2�p�y&#�˰�!�}��D�Nz�6�iOw��w�m�m�n�&ٰs��7S^J�>�,�cFM��#�ȴ�e���2iȸ��|�������^��[��3_��                ��s�r��i2�<��8\��$��N�.�e����X/�������*�nY-�6� ��A�Pp? ;��3CN��2m�ݮ؞)�k�/��8GN������7<'��{R�X�T��                ��vsg��.���%'�;N�y�$��֧�>'��8o�����-��c۫�����ן�'7>�*�@���mΚx��;���lK�a�8dl���i�u�U�^�߿����lj�*                �{5���'�O>]N�x��+�)u�ާ����xǌ+���G_��<�ʟ�ϯ�U:ҝ���.��)�g���.����dJ��c�뱣��~�q������/=$��s�`               �Ɩǯ�v�\pę�(�H��'�L>��a����������S����]�����UG]l�2z�(h���cft?�|�����G��R�n_'               @.���ە��v��r��i2ٲ�EG�����������ꇤ=�!q˂��!c�W�%Sϕ��������G]"WyQ��
���gݫ�               �dP���3{�Q����#%WL:N�|��t����~#?|��dkG��M�
�v����F.�v��ʑ\dWu?s���[p��߾�}�               ` K�Iy˔s����!#
�I�*L��g^ݽ2�/V�N���cUt�E�}H^��x����#/���o�۱���O_�A�㫏���-ym�z               � �ESΖ�f�SF!q����ێ�T.�z^w��������亜n{;Jɕ�/�[f]'C�
%�Κt��6���s��������:               ������Sn��GM���(��Nx�\>�����䑵�K.�ق��ᓤ���ʌæ�{��ws�\t�Y������<*               @���g�6y�1Wu/z��c��J�Ok���Ǿ*wm�\�swW9r��7�|���+؛�-Ç�)���I���l��)               @T�8v�T�q��<J�fgL<I�s��|��~/�&�
�c��3�ɱ������!�Fϐ�|U���c               ��.n}ñ��l�p�#ؿ���� �w�4<���Z�:g
�~���~�JNk-��n����'�F̐���'���               �lW8Z>x�B9r�A�l۶M�7)��	�r�Kߑg6=/�`��]��-����g^-�[n��e�֭�����H��ˤv՗es�V               �儱3�γ����a�ޱ�v��}_�oi����<:�i��s?��n@��j��q^��8�XAＱ���۞��G�O���噭/
               �io;�R�s�lq�#���}`�����.��#e�	�K�߿$��e������_$�G!����{t�w��㮑_��<��a               2���W�m'�K�{v��իW�Un��y��Y �yB����=�3�K�Yp_8F�\T���s�r{�t*%>UFN.�y�g               �'G))>�6�|����������HˇfΗ��(�;���Wp�2|�|�J5h��wz[n�����L�!G^'_z�{               􇤛��3�ʹ�O�ށVnߗ��N�<�����嵝d P��F-��B%
���r���*�}G�S���w               8�|���r��������o�j��H��_��;��@1`
��G!w�WJ����޳�2Nn�~�|��               D�I��YH�����r�u�wJ񔛥��/ˆ��2�������.�!y���9�r����&�uG\&����	               ��r����%轠+���-��y�|v�
ّ�)Q����A#���P��֟����wR��<~����?	               �[�N�YΜx���u��7J��;��#���rIy)��H�%��W������������e�ϖu��dՖ               8�wͼZ�>�bA�����o��H��Yw�g����_�?E�ஔ��3�ɴ�z'S���TJn��v��Ε��k�                �cWm�u�u������(�+�}�|���KTE��~��k�Ad��ޣsW�Tw�|��#|�               �3a�XYt�q�#�[n�}`��3��9��L�3'�,����DQ$�'�?^n:����V����{���/���                �.�Mʇ�-���`A�d��ޣ��K�w����e�ؾE�&r�a�Ce�wp�F/e�ܾg���9y�q����               �q��7����c��/��BwG7[v�퐊��'K�R+��|��/"Wp/;�}2�`����(��8�ä��ۤ����t�                ��?^�>�bAﴵ�u���Yn������3�ڶ��{��\�$R�˦�/gN<Ippa��Ǎ'�'ﾪf��7J���(               ���y���9���-�ە�}?�+�w�ۏ9F�ɤ�g�u���&k�^���L�ݮ�~���\T��֥Sϓ��I_��                ��8i��(&8�(�ۭ�����o�?��uv���D����[dH^����Tn��6O�U*~�1��R              ��9i�rɔs�r{��M����H~���(��8v��3�T���Yn?~�L�4i���p���+�O�H               /�rd��7v/���Z���-ǿC�ǟ��k��-�c�ܓoXT��=���V��K����6               ���#/�)�'	,��vkH^��<����W%l�ܯ�~� �^n��ܤ�:�R��J              @<&ˍǿ]p`Q.���b��r�s��W��&a
���t��c���@(�����3�{�~&/m{E               ���1�r�W(ؿ�Pn�\��ͳ�����Y�j�����"�!ط�Tn�3�o8��5               2���>�2���r{�s'�&�F.������Vp�s��ΙW
�m���{�A=u�dVq              �q�s�J�m���-���>�m�?4IXB+�_2�\�?L�f��n�A}�˥�O�
               rS��'WL�P�o����I'˄!c��%��m	��3.��@.���舳�kO~O6��"               �=�O�@��
�l ��-G9�^7?�U	C(�S�/��N�-���rŴ�kO~_               �[�b�o=�-�7����L9G����ȮT�d[(�+����J�����/�o<�C�tv9              �Y'��)���-W��VA"_.<�,����l�z�}D�09}�ɵr�5�`��6�yd�              ��q��{�������M�(����ȋ�Qp��s�u\�n�Xn���Qp              �!����I��%��֔ᓻ/o{E�)���'�!�-����i�guOb�R�              ��ϖۓN�+ȑ����~Fn�����#��~��J�I9s�I��               |�O>]�[��ۭ�?C����J6e��~��h+���L:��;              @�,���+�G��?d�L>9���g��~��Ywq*�['�I̮��R              ���ı�J��j�8��Rn�qڄY�Yp�(���)q�r���s���g               �]ǯ�n�2�x��3?����Vp?a�LqW�*�����;��;              � w��$��Xn��}��y��ueeY+�7�h��8�ۭ�fP              `�5h��+-q�r��pr��i�����?ɒccZr�{��:z�TI�����              ���������\n�qܘ�s��n[��G.qC�}�����#��U�^               <3�&qD�}������J���a�K�qB�}oS�N�              `���Ů�*�Ȍ3"Sn���8"k��J�}���'���l�x��O�	Q?1�Y;:�պ;����w����cG�����*�|��:"ٛAs���������i'�����&{E����o�vl�7G�g�҉�{�o{e�pI���ӥ��傴�ou�L�����s���~c���<B���gs�/��9j��_�����k~l�����3�|�zIIӖ%K�8��ma�G�����k\QS�"���ʹ_)�O�?�~�߳O'҇����9���3��y9v�c�3	G�/�����9g��_(��c�w҉#�#��7�;׸�����sV����9�N������>�%�k��$��g��ϙ�d�!r���+�z�����MM�#\ϝlN�f���y{����%��9�|�����#)���W����1��1�j�v��_�{��ҫ<�{e��k}���1�~a��ϻ��1�W�y��$��Lߗ�xW�y����'��z�G����J�ɚ7f��m���gp�c���~�����z�'����m��ǖh�}�Ùh_���c�U�X{��_�9�ń��k�gz�7�~cc��e���=��q     �@���ܾ�����y���kg������ãW�ΤիWSn�#�M��|��JK�Vnk�����of���g>l��x�<�f�!����<QN��z��R�>ٓ}�JHKqY���7��~e}ٹ�/e���&yG�'&�Z��-*�W�����~������ޓRsu#����^iՔ����?n_��{KMŹ"^���f��;Ot�hiNh������}��f�����GYkm��f����os�􉯥K�n6���%���׿yC�O��7̣����,����;���E�jy���'��o������3͋��ߣ��Z.�����'M�~˞���>�h�.9Ü[�h�n%��3�(]Z�	I4�T��}_����U�-{��b��md�wfܧ��{�K*�����^R��YSO�3�o�Ge��S�)�Ŀ�E�}d�7sν�X�X\�����~���yT���s�Z�E�n�S��W��d�6����}�^l�����u��﫞�-��U�����#{{L��W�,+9Y�Z���!����^�_L(�aAE�co�������Q����$ǌ{3��%��3�uڜ�|�|Ұ����}��%K������y��~qku��%U�ym;G)����|��+f����������R�����ue'(_���=     @�,.��J\Pn߷ÇM��6>'���7('+qaWn߲eK���r�5q�8�|_��u���=o<�R�K4>h>}�uY��}GꔨK��a�Ӻ9���ȼ��6�u����?d>}�����ڷ��e�����Z�$���5��Ջ>���d��L�����rWYY�� _a���ߛ�o�/���U�(�R�ھ���|h΢�A������͇�W,-����k�/�[��|����s*�e_T��G��͵�0?�3�\#8(�z�S��*�������|�yu���ܳ��)ǩ6�9oTw��))��_T�.��XP��'��ֺ�O��T��﵂�ړ�WL�wί�?���Դ���J/3�_'8(��/�uG'�_TU�Z��Q���7��f�'͑{�R�z�A�d��ʝs���f�����|���s��������7�￿x��W�l�'�����O���VZn�'�>��A�_����d�)�����7	z�d����Tͯh|%��+�� �MK~�u�3�ko�'���������5A������ue��|�Y��=�^1����$*���#��E����R���}��y]k�g�     ���S�r��M:6w
�cGKPn߿��$�͓N�K�}�����ŕ�쏯7��Ѯ|YKu�|�|[t�쓧�u�d_R�����zE��Ϙ��V����n ���ٻ*�����!�[YcW����|�־;@�Oi�w�\������C�������*����Q��d�ߔp��K*�~�_o����͇k̜s��s�͸,�'�}�w�]\U����zEu/�o3��=fα�
�������PT����zs��^4�m�-���9�d��X�E)uCɢ�_��כ_^��|x��sn4s�
���>���-���.�h����z�U�/��l�)��EV�����)%7/j�i|�=űw�9�]��}�QN|���#���:7����?�ޞ����ʾ.������d��mJ��������z�+�lQ��֚ү�"6��}�E�9Z�S\����z{��yym�ה��D��狿��έ&�����sq�--ե_�J��e�`��9�vW�ۊ5|�?����z{Aԭ͵�_�Z�!�����(y��������d[K]�״/_1�~�      `���ǟO(������g��~��:������fr{u���QJ�����z��,��km^V���*Qc{I����P���5Z��@�W֯\Q[����?5s@|n��Kf�?����~�~AE�=-�JՎ�q�K'{)-�	7����Ζ����M�_h�.~�S��s��Ō�'�$y���`+(��s�Ҳ��1ߑ_8J&�b��SII�e~U�go��W�ז?�k�Wd�`/f�?-I������~"<�����J7���f��,�KZ��\�wIQe�ի��9�h�+{����;�9\����g璹�u�V�>���k�/}�Ow��G�b���ʽxOA�_����KK��v��^M�������d�����{ EU��k�-?��f�5]�3߿�J򒠫���E�o�+;������ڣ{1ٯ�K�K�5���_{aE�m����V�т��}��d¹d��w�jAeÏ��U��8���s�������Z.�S��b���Wԗ���Č{u�`/f�YS���s*��=���?i�Yt����3      ���bs�(�ܸ�)��U�����&���9l�
�x������|^Q�L����KK��\y��￘��`�����%c��ۻ7ז��k�AGe�=L��|�{+�ޙ�}�ۻ߳��ܔ�qOٷG���yXz����@CƲ��o�+;����s(����c�C/����n��>,nx��f�پN?�(E�t�.�{�w�,�i��>V�=u��K�N%��N�0��_=ǽ���.c�ۻִ֖�c��&�)�n&������ej��5+���N��	��|����w����fj��)&�sR��e�1�~U��n&.�a��Z��lOR��p�/i�W�	�9���p{�����J���鿤E?�'Թ%e5����1�k���o)=�����D:}μ���p�Ǟ��3�����XA7{1S��3��nC��a��|����d�7�X{�����F��s�/_��}�F��K�K��o�R����_JJ��9�h���Pj�Ҫ��nʌ{�%      x�Q�r�f���{gԠ��|5�����}�p��7,���co��Q�9䪹���X���-b,�-�R���U(1���g=׽�4���E�溲+���@�����Ġ���,���S��⊚�+<�l��}@�.�P(�������1Z��^�3�Ќ������2Yn�aߐ�3�<l�}n���3߿\��2�bY�
�=漿qMK}����4�g��L�����zKEY]Ƴ�+5/���\ĳُ��3s�+�t��������{�-�_�bi���L������~� ׽䎊̕�{���YV|y��<�����DZ���I�L��{̯�Y״��
�ҏ(%��KVZ��]?E�+X��ٯ�/��K�G�K�9�^��K��g<�9u��|�]	y���͸W�z��/��]���f�Z[~��͸��m;�oL:��6�L���|��.�B��#\�mWn�7xrq&��=�W�׵)_�9g`�	�f�orU���2Wn�aϥ��y��z��d     �Y.��)��ް�쌃�܇�p��r{�ˏ}���W~G�N�#e�+�h�.�����Ę�ug�J^;��&ㅻE��k�)�c>��Ę�>�:�f�p�cޢڿ7W��%�I����z�U�/������֖�1'�ߔ�]ǽn^e�w=��-ե��q��*����]��*���]U����V�����K�kM/��X����֚�[�K�I̳�w�k��٘��]{!eK]٭�`s��>���"�9�f�p��^��ZW6���&yGb���{�V�ϯ�|髇]ٷu��^���^{	I\�����l�Ӯ��R[>[��W1��O:�z{�K��i/�[^]z�(�+3߻S6�<���^��>��|�ՍZ��={W�;m��g��寚�7�����^BT��u�un�SY�&[���[su���1�k5p���oJkGԍ�b�l���W�q��`��     ؇�y���)�����q��?JN�\D���
���<g�ܪ�U������o�Ԕ��<�wK\��rny��_��ᾖ���E�l�+W/.*ox&ۻ-���fKM����&�+��_��t�w;���[�5e_3���Hl�������?j�.�����.1�E�UB�Eu��c��g?Gb�Q�����g{��5����|�=O�J˒yu�e{���b�QR$1�|�DQUã������_�q�l�}�Ĕ���.�j�C��;���׭ե��xS!1���OQe�ﳽ�u�i�.�5ϠRb����+*oz(��]X������j��Ĕ��υ��ym����ҥJ�$�<�KK5>�����n�.��(�!�)_�E����~�*��RSv���?$�ҾԔT6�2��5�)i�)����      ��r�J����egd���troa�����X@0]�r㶱+�ڿRN��m�U��L�N?�i������y�Ŏ�x��ͫ��K{�6n�<�����?��w8�b�}J{ύ���1���~�NqR�)Q�w�]�޸ulMX�O8�S���>v��1���[�-k�:���$�7(�r�vN���{k���χ��N��p�f�&1c�1_�m���ڿ����]7�9g�Č�s^�m�gB�2�7��d�)1c�s����a����/iO�b���3)�_ߩ�C˾ӑ��k�3��H̤����/�TX�w�?�.�y��~�Č�~�;��Dh�O�O�i�͜猗�I��4�k��_���d{^�{�����֛��,��낮OIG�}fΙ(1��N�G�ڿ_��iݑ���9�M     �~�t^�@(���q���{�h���%(�c�<Q^�d����[j�Zͧ�3���P���[[��m�~��LR���{{kk��-�WI�$���ٳ�酵{k���Ҧ8��h���̸O���9u̸���v�P�G�̾�Ζ��5e�q\�._�w�/jJ������M&��}hE��$����K�t���y��m6�W��H��)��af_RҴ����^�Z�2,y���w|�#���l3�ۋz�Gb&�%�����EE][��U}C��$,f��D������no�.��(}�Č+���~WX�/-m��\]�YQ�Tb���S����;�ڿݷyme�j�G������3��?�i�Č#Χ���k�6�֚��1���     �n������q��w���~2>�ʕ\A�������K{kK5ݿ ��'|�:�e�S%1a��d�ð���D��+$V���6n������Z�g/.p$&L�6n�ݰ����5鄲�&{�������H%��dZ}�L9�sRz)�oٰu�}a?�n����}�����6�Cy�z�3���d��u� ̜��J}-��᧺$/��Ul^����}�ֱ_�y�^��wS�)����0��4|ח�~R��$�ɏ��Y������_�yt*��@���*{�۝A�{�~��A-�������|�;���y��~k"�>�;d�ZwNj�yt�h�k�o�}�Ą/���ӡ�	��.�Z)�O���df�wu9N��o���)t��'�w'     ؗ\�Sn?t�b�./�k�e�������W����C[<�j�U)��a�T5��RS���>_b�U*�WU��ZS�;�D.��p��s��E�j��R[�[3
.��0��+�����7�i�.��(y�ą�/��r~�����[k��E_%1�D}1���{̯�Y�RS�3��[%&|G})
�/_o�����m�w�+EE-�����޽��c��<�wHL�s����z{������O�)1��|#���{�U�͸��yF�%.�ܷ8��{�U�͸����&�	��o���x��{KM�w̧0'��s�vw3�|ی��$&|�7
����ZS�-s��Ą�����y�y����^@~�Ą��TT4���<���k��s      v1�(����|%(�����q�(����z��t��%"����Hl
�	ID&{s�c��O�]Id�7��.��H8nt�W�d�bSpO*�{��JIl
�	':�w�9*>�����1����>6����w����ͱ�;�d�U|
�	��cSpwŉ̜�'���]?B�^9�k�cSpϋԜ��M�=�ߖ����*6��R��瘱)���V�����=��;     �����o۶M^x����.|�ea���S��L������TD���o_�e�Z? JI�[�����q��}��#q���y���JD(qВwW9{;�׷���D���|�M��Ӓ>l�a��P��sܸ����yX"���:&�/�����W�xj`��-m�����KD8�����cܛ��A�ID��{ �#�E<8�;E�N"��L����{s:�����H��\7�ދ�����ɾ��H��1�-��32٧�͸�Ǹ�̑�7IG�:�׵�҉�dߕп������~22٧���)����       �#����)���l�ۭ��Б
�nفQn�_�NA���_�dɒ�4k�I�d2�b��D��_�=���9�(H~�#�#٧|�r����Oq}�{��M����0sNd.u�n�ob�B�7�<�2{ɒ.�]�zV���JIη`R�[[��)2']�n�܄�RJT�Rۏ�֯-���y�3t��緬�i�}��.�ו�쒈x�m�Gm��
$�u����w���iuK]�.��`�qf�o�XT�&1���k��K�+��J�K�����~�DD���.�)msD��K��e�%"JK_o�)�b�sFJ�K����;[6JD/_�\S�Y����ֺm���s*�6�Ԕ��3Fr����ŕ��$"��6�c�zs�+9.���%UկID��4m1��u�X;^      bnW�]"����=��q�����ȼ��'���_[�A�i��DHii����J��Cڗ�%B����w6ה�S1xc�W:R�/^������u�2Qr�9)}A"�;���\S���,9�7�R!EE-��������̸�T��"���җE�Q��|��W�c�Kf�#9NG,{{AgKM��]<Nr��s"��R��k��~��8��_��Qʞ��"9Ό��$bQϙ�I��ܸW��?Sr\Z���ؿ1�-9��D�6�^�|�݌��e��cƽ���c��_��qE=�Er��      �c ��)���lu�3^po��.����N�=��r7I�(���{9�Ɛ�T�����s��!W�Ȭr�OZl�9_pW���>��JI�W��s��Z%$*2�����},���I8�J��|�-f���A(-�r�A���D/{3�cq�U����)&����q-�ϩ��(~�1�s"��V��s�������72AG���M�*     � �:V�r{fl��N/<����v�|O\Ǖ�`��Ք�3d[�������R=�*��g�S�s����iN�:��'r٫��{�U�D��>��}FsΑp$z�^$.s�D.{��	J��}��>��?��Q�>&�^3߇&���Q�N)�c��E�4���`^]i����x���)��d     p`�Ђה�3'[:d���k_6�o�q��%�l�}���/��r��~W�1Fvi�����bQ�Q���s�04��Ik�ܸWJ���hO�ȍ{c�Ā/~�O3�8��/ћ�ͤ34��}FN�S��:��gL���q���cp��EG/{3��p����c���7���O�{n"�츏C��
%b̸��uϥ#���	�"zߧ}N��      �~�&(�gV���/�[�wn�|�=�r�ĉe	�뺼Ԁ�z��D�Js�R-�jl�/�i=Q"�f�Z#�bpm���7�k=.v(Q��ޜ6����žM�!QJ������tVS������*��eoD�9e�8��1�}�G�r�J���9�J�{R1H_��e���X��H�h�9�Q��͸�����74���|���ބ��^     �0�E�)�g^�.t�J�}�΍r�D��̳c@k�8�;W���{��LV	$1��s�D��e'��Dn�LPN��_YW6��%����;%��Jƫt<VwD����/=Lyr�Ā��K�ܻ�rDJ��\F��	Ǚ&R[[>Li����K޾�u�J���~���~���Ʉr�J�|�swv�H]T�)	QS$B�����m2���x�{I�s��`W�hL��-Y��Um��1(S�ʙ�웛$�]M��M�J�d��<|� �<"���o������}���nYk^k�~�f�OL�������$�8Pj������ʝ`��#-нHJ����     ��@��r{vdkd�ྦ�5�*����W�����SK:�D[t���z�D@�u��]J�{O10�<���X<���i�D�뺁�������>_�q�w/]tgK$��|_���
�l����K�w�=��c�T�m�p=�� �єs�	�s�S�({1�����yZ�9'�<�*gd�҅��/���WZ��9�0眀�����[k�'ϯ�{E" O���>�԰�e�S���_�H�&{���{:��T��.!jHk]ٴ����%:�;Or�@���~�\��ԗ�XP��D��c�iJ�k��&�8��9�R�+�Kf�4>-�eĆS�(��ۅ;���;��[��'��D�jO�lf�>�m5b?��9�G���M��	�m<�|�7��I#7�d��>�Kt��߮{�}��[�fbM��ɮ�D��Wǜ����v����Ao�w�����n{}�����$&�X7Kk���ۅ9�-�d���W��=7��E"`em��J��}�.��{     �Ly}�z��R��F��M�={^ޖ�JJV
�/o�D��M(�g��[#ѱB?�X Q�T�I]d>��D�R�R���N?�7��1b�O���ͧߕ��\dѽ�0]A�Oڌ�D��ߖТ.�]���sTwa���}��_�U�˦��������U��W����3��c�!@\�}���e� 3�/�]g�%�C���o��/J��.�K��Hb��9AJw��zv��#Q��˂����c/�
���k;�WH�cm�o�+��Q��w��.�������#Qp7�%�|n�і�ƌ�\�}$
��X渷c��;I��k"D'�}$
��;�ڿ��y'O�|M�(_�6w�X��s��q���d�m��(�����.@o����B���>w�f���>m����S��>��s��č      ��}eM�Z9rd�n6L�=��S��=;���_�`��r{v���\�O���O"Pp���ղ�]A��p(oJu��ه^p��w޺V�;�����ƽ��>􂻽�����Y0�3���!��̸�]"Pp���j��Anff�7ս�Z�W�:��������xk�}�7�����5¾0t�=�>���۸�*��f�ˮ�����{wHD
�̛�~��G��g��@K��9'w�w�(����ص{ΉD���k��^�^Y5P�^w�M��f�X�u��d�𧱔t�9�7٨#�Ue�EMA
���v�V"����h�	;{ߗ<7������5;�V]!go�7��O�s�e	6� �xe��͸/�{�=�^"!ظ��XkK�}^��n�{���D���s      2奭�D��N�=�^n{5kYg�ྵ�M6��,���(�ܞ}�m����O���~s$���;CIq߶biըy��e����L��m�ø ����$,��ءӁV�2?���חVVְIB�u�kD�~������c���AN߳Oj��{j��̩�� !�8b�[E��A���7�m�]�dp�����MM�/_/!�4r�UZԤ ������|t���N߳7s�%+��&�-��*�֚�+̜�U��޲s�07������MKN*^�<�[謨/�Di�d۝~������y;3�/h�-�<��.�+|[��]��d۝!k{�?"@�y�s����)��^�-�.�Pi5#ȶ;B�sl�AJwy�{nӲʩ�U�/I��kJ�W��	�m������d��g�XZrԼō�K�̼w���� ����3�p~/�i-��3�5�����ӕ/'�6
�9��c�{Js]�̢��g$D��JOU"'�6
�0��c͸?yym�q+Ꞓ�,+9ټD<5ȶ;#p���>�I����bּE���߽��g�6�q�赕9�?�������M��,-��ٳ�l���e~�#���+�83�d�P�^к��X��� ۆ�=     @�<�e�\:�<����������ܭ�7=/>S�F�=����$wm��^�Lp
����T���2�~TB��� �٢��C´9�!�C����t<�~��]�٨;{/����'9}��U���}���%L��P����9��S´Ɍ��y}?)t̹N������"-*���f�9�q�)�.��Wf�wx�s�HB����e�wa��*a8J�T±c�\�䫻��9�&�i���Rp7�Z'���8["!�N�c�&/�q?"X������]$!r3�N:a���s�[���l������t���<����!�
}ܛc� ً6�����|v�����]*`��һ$Lv܏q�y;{��tڷ�io�9~��~s:��Vc}_ӷ;{ϳٿGB��|P�瘛�v+���t�f��H��]Aߧ����;d���oiV�tg��E�)s΄ K�RJ�Kޡ��(W]��I��|�c�C�;p��q�yN���!g     �)�6� Q���F�=Oo���[Y+�?c���[p��{qr�-�MH{SN)��������lKM���l�	i��%�,�hS����D/6�7��}km���IE�K��L�)�K�6r�����Ma�,k����� �n�]��V�����u�ZԴ��!��e���]g>\d�:��;�h[W��{��̩j����fyM�Ufƾ0ȶv%�г7��Լၶu�*2�/+����+̜si�m�u���a�s�t	��#������V�m�.�܌�˃l�ar����X;=oD�mq殬^�tne�*	AKm�e���A��wG
{eS[~:2�&�;���>֊�v�|s�{U�m�\�S��������ۺ���Z]�4��e����� ����N�6ۂ}��@ۺʹeym��a�,����<ߗ�lk���}k��>ض&��[��|nAU�����3D����=�e[��!{qn\Q[��yu�Il�Z��A��F���O���d�y��#�֚��|��Vj�~D�*��w���9��e�6���IG]�\]zVQe�%�nf����޽XD��;     �M�h[+;�vʐ�`���`���?�<��<�){8d�������9�r{���>�~	2l�!��犓�ru���Zɲ���:��.�(�;%l�L���A/���r��|z�dٽ�*Gt�Tu��ׅ�����`�cm���u��r��Ւe������&�_��¸����sDJu5�O���^:�&����>e~����i7GT�]���ĥ�w ��*V~�C=�syн������9tg�{L��d;����!��Ơ��q/�Tʷ���lg����Y��7�qH�(�S�+�,Yr�yd��83���1�v]$�1�?�}���1��F��Xk�o�o�C�~��{���#�D���Ι=��Y�2��{o/HmS-���9ag�z�вO��J��Y�ξ��<����+ʮ7s���?�9��9"�h;�iY�*�f/��b�z�}��f/ᆿ�ʦ�wL���&�ӳ��}K��mQ[U��V�������P��Ju�^����lgo��I��o5�>`�v�	7�C����&�S��Z�ze��^���A��wl�B^,b�!f��fJ�K�,���e�u      d��}yj�sr�ēC�?���i{M�tl����Vp�Wml���ٻ���{���3��� aWA@�խ�֥�V����m{�׶�%,���mKo��V@	Xm���.X���"��Y	ٓ�d�s��9�P��d���9��w.�I���9gf~�y:dl�h�6��v�FA����7Q���5�gΘq��5�%�f,]�M}��_��h@r�.���j�+�6c΢[$Kt�K��0�8*�c�E{$�jc�}����5U��3�.Z$Yd�oU�LJ���a����U��^7wa�e�T�"EK���ѩ~~],��>���%5ճ�!��FɢDI���)�~����ŋ�g}Ke�ɢ¸�f5��K�4�{��B��wT���,���q��B�y1��*ھ�>��dS�h�!r\��^����g���U��d�.�V�����;���5��M�~�>��dQ��l��I�~�+���~��H������{��1�ɢbK~���SS�|7d����d_ �3'T��T}�=ɢ�����OO���\q��I3{㌉���B}�mɢ���ߨo��T?�5٫��z㿚sN�0�E__~S����i�����\ېf����D�����$��u�/Է|v��_����W󽾹ė��?%�W�[����E*���o��T?����      d��9)�Snϭ5�����Vp��4o�+��0�_�r{��v�ol@��+<�����O#�a,Z2V��/|L����Y�ؔ�pOrÛrz%󰩲����i,T���V�KT��0�c��6���[U�}jܗ�>���U3w\7��G%�̯�������1�ܐ}BeoƤԗƅ�%�_�`��kg/|D�`���?QԟH��.(a��!	�������7K�g�f΂�K,���c�T��9F����xX*��4����+����e?��-�>��1�0������/N�*�_�s�6u���dAMլ�q��t��F��=�����Ӛ���θ~�}�*�o"W�s7\���u����>���ߜ���Ϟ�N�_I�����\Уr��N��$�c�,�������!Y�淙�?#�c��\L���m��SܶC�|������ۮ�����K�f]��}e:�pÜ����u�t��|�U�}[����vɂ���3Ĳf�s7\�������)���Ըߢ��m���|��Ι��1�0�̸��B2�0��}���Ru������,P�k�QsNZ�n7����wm�X����*����7f-��J�����ϭ�VB�cA9�px�����5U�f�]t�d��9N�9�J�u��g     �I��\t�(������.v�Ղ���ײZp�ܞ{���?�!;�v滢�rR񘔏��o��9�1��ɠ��Y?T��w�9F����5����X���N���L˺qU�����)� ��K���1t�S�	�k��hW�KN)��1�e˗T��еs<)����{�+�o:��U�^�	�k:�j�9-���q����T����9�ZR]��M����.\��J��g�%���K��F�2�YZU��k�.zX2hi��o�'3��9�.�4ǃ�;"���a�S��d�j�T���$��VW^���Y:��œ�X�ǽ�眳��^��ճ?vݜH���ò~��1��s�Q�dߥ����,�0E��9'���%�t��+���î�]rv��[�,��iVl��.�R?�Ju]\��1"fBv������61���+1'ļM�����௒A�%_s������n��^]ߏ-M�d���,�Vu��w��E�J�TU~U���nP:���K�wɸ���7�Z�����R�߾l���i{�Y��Gݱ���i����R5�Ԝs�d���K�i�b��}\e_�죝i����K��9�Z:���Z�F�*{�;�i�\�N�}_��S�9wJ��-}�N���RqI�j�I��n�9bԨ1���|���g�������Я�[���      ���ǵ]�e�IY�z��s�/��m۲�5���{ ���_H>\����������!ԖV�]�����g%oPTW�..k�XrM���j�,�#j��^NN7{�(6E�+�eb�;;{ӬR������������mi�5;{�|tI��k3���~�%7�̾��6�?�[��s�i�g_������L��u�yE]m7��f�{���6�f"7ب�O����(4��gMu��s�"��F+�U5��v�d��}:wMgoY�?�̟5����,������Z�#���6���2����4��R��_^3���/X(�7o^���V(i���mV�>!���;�4J�ҟ����}Iլ믝�p�8�?��_�X�L�X��v�֫k�����'j��,��ׯ����0��������N�X�#�.ʾ-����o Vsν5�+�s��E7:����~���4�j��^:�vM���K�{=�W���8��^��,��=嫳d&�=�穯�I3���N����#���2G�_���r�5��&s���Q�?V�����if�����OّiC��Ss�]jΙ��_f"�#*�~�oN;����}HgTZǰ�7�?/V�7w�����ѓ�@�?�����朳-�a�P����{��ޒ;��Y&�?rt������K�`�m�t�7R���s.(��֟H}���O5U3�5u����٫��qk����ߴ�^�ۣ]��      �NwC�Qp���+�J,����j�=a&d՞u2}���:��ݡ1�lߥ��e�XoƤԗ�$n�`�O7WU^i�eάY�ڝ��W�>�ЫYr��{=�&n�W�u,{��T�W�c��3��đ?���_;�4���0�r�x\���H���v�?�������-j��Y_���Չ�f��ӌ�u�e��N�M�6�%�DT��Ei��^�[n�ye��?ө�o��sj��v�!r��[����Ӝs��%7/��y��,����:��-�}�)��V��q��sӜSHw""#��iG1��[tK��+������f'���7�<�
��:�v�x����舆X�t��+��Zps��E3f|}~�ߟ��O�D���x��[qϸ׫:w&�*����cg/R�εW���k�����;{G�غi��������ץ��5f^���k�2{�'��%+��x��s�����t����DH��S_ͺ���o/��ti����Y�ȓ��Us��ܓ�U�"'���cAi�����u?ð,�75�g^v���_���N|5ճ��j2���_���t��-Zb}�e��1�Xe_SU��s����n��k�č6��Lw�xn�:���1���U�?����^SU�e��_�`�4�l[�>�̉�iܷ��^�5� �`�yn�t⨖��t�������N|�XS�>;�˝8���oS�7�9��BG��ɄQ�����v*�[VN1Ͷ5�]����4�����x@&��u��ڹoބ�-��y��kf/��������ڷ�2��;q�.�      ����W�s�~T�R���A��=^hX����Ղ��l݊��)���s���^au]�5�U��
�����>�����fqlɌK�R9�m��99Q���e��J�5m����C��ٷ���W���̂�.���WV�o�L�8K�gOR߳Ěa8�}c��~��-L��pKګ~%���d�L\U3�O�Ŋ���i�wӼN]9:��.Z�҉[��ש���_N��|�5��/����X�������T�s��;�_P�]�J|�p,��]�r����^�ȡ�}��#	�_�����P��_��o��f���1c���um����z��j���Ɏ�/��2b��5U�~Z.]�j�57]�����T�z���Z���q�"�ʾ@|6�إ�\����[4g΂�T��h�̉�q���u�l5�8�lZg�K�n���v�x�\�!�۾t�쟇|�0��Ο;AԸ�K|�a9�����7S���}�^��|�#�S��c��]�9?���Bu}ߝ�qt���������8�}�˲�����ee﷌+bnS��_&
������T�s�-׍�G����Wט��e8@�����55�\Q>Ցc�|�+�~k�ҪY��&�gμ�3���V={\²n0M����7n�F�D_c^Y>͑c����L#���s~�(LT��}͍׎5
�n��u���I�N�]*{}����Q�_�P�>øT]�o]2��}fA�Wo�)�g.�Sh���0�p${}��Έ���5�|���}��q�E�9�����T�����zˈ}S�H�N�=*�Qwe��#
�q�X~�x�@�7��oJ5�[��і?v}"a}K�9e�.��ܓ�|���-5Օ7J4vS�v��M_|n"a~�ˑ�{ͨ�k     �P���*[;v�	c�y��(��GW�Gֵl����z����-���"G���)���i��T�K���J�I�-�(����1B��n2��T���a���ؼꓟ������o��G��,�\�0?jXVa��(�ɋ�Fq�W��U�G8�����2���8����+�����G��|��kj�-�"ŗb}��c�gﾝ V��O�"g���[7��~�������3ꈦW'{#T8]�j����ٻoܯ
6˻Ըw.{c������Ú���0��{:G��7o�!����K��5�|���bI�g����v6�2��f�8�����ͻ�:ǯx�����+�G/Qy6���V�"'�~�ϑE���o����H)�9��^��*��TUީ栻;Ƽ|8�/��O]�}ֲ�P��h�z�g�y��Zj��ˎ�Ù�M����4�d��;���p�/�G.6��Y�[*{�ذ�K����e����jܗ���^�#K-��y�i}_go�uws׸��.��o�RI�{����V�T�;:�rܷ��Ï�aN�{1���?3C�߯�_�ƽ�n�8�ҌK��[��������^�ءo��s,�u��I������L�.�4���e_]=�x�i^dg�>%�����]�'�/�9�B��2Jԟp�/����^Ŀ��s􋟜7/z���٫�/��l�2?���8���
5��^^������!+Ig�~����W��2���u��Y��5u�����R'眗ո7]6�_W��B5���B�PV,����?�-5������F��}��w޼����Uޟ���)}��3�V����w�J��?��7չ�5�����Y9����Ǵ]`����|J��eN^�l�hp�K��i~�ߙq?��T�7,�_�5m��p���x�!�g�5�˜�s^Q�kj��F���*�tw'KR��"���7��T����sX�����'�gT��v<{5����     Ȥ'v=���;�vwy��%I�	ɶ����{��E{k'Qnw�����/�?d_0�ߐ>�t�����o��e��3�7��]\U��O�MbX�b�g�	�\��Ԅ$N��9>����d�K�+��m�#-h��"�.Z;I�8RE8ǧ{&o�?��O6�|��^�K���%b��o(М�^o��=�����q�.��7���"��e��w��uZ�2O���#��g�W��������=��+u�ܫo�Q�R�ϚX�ڧ�C|��l�?{�gM5M�T��!V�w�94d�eM_�������o2��>�9��5TSU�Be�YM���%���d��p�X�s���m�w�jM�䍰��}X��ա�r�C;�$d�5�����^��>���MÚ��7$v��Rd�z��eK$�3*����l��;�{A�}���u*��&V���g�T�n<T�jNh�8~G",�#)-x�QQ+!���ʅÝ�1%)�������.2}�:'�}��8�.ψ��|ߩ��v߸���q���^g�k�V�(�x~�*���h�U��^�w�U�SU�'G{Dg_���#�!��q�o������ˢ_�|�)/����/�o�^E=E����|�e����t��.�>n�*�&�ġ�#��٫k̯vT��ո_�������峷�Hf�桓Deo����3�1��^�w�K��7�Ow8{���Ɛ�b~Eg�=�}�#{1���<����3�H@=\n��[��P��e��^���G��Qm������v�yD2�Ni=Ϸo�pg��+)�]��F�_W����ڑ��5U�W�Vd����T�U�u��M1�տ����'v*{S���ǽ�z�K�����ڵ#i �/��t��}z�[�Iv��WO�o��B�����N��d�>���_,�Cg�>����:{�����ۯ��0{     �Lz�����OHY�sk�Pnw��΅�ܵ'w� �:�CR���L����ѝ�/w˩��8���[��.�]j?��w����^����[�o�to���^���ac3���]��b�.��ӯٗ}�%��w�ʚIzܟV2ֱ6��`�[�5��~���ܜ}��'����E�KTڗ$�����F���^�4|zi�(�\b?T�����h��@��V�Mz�o��S�{_f�H�}����^ddx�?��ӝѫ�䝥�[����2�������qq�+�}�?{�F�,���\��l�
{�Opleٷ(�]�Ҿh���]3�l���sm��d}V&��W�6.T�_������2��������W�5�Y�&8���[�����/�}�k�d�����sܺ�l2�Q��^�{ѫ�5����L���n�~u�Y�VsNE���oT�){k��3��n���F�ֳո]��&�d��P?�e�/��H���X�hu�Ee?1'��W��~��\����V{����a9�J�X]�4{}}����sj��7,     %�DL��{Y>�K9�v�ym�&i4��k����g�_�˦]���(���̫�6����s��r��+O���>�6�-n��6�[�1U�ͦp�+W�Oҫ2�7l�^y�6��e�۳�m��a�[Ը�q�
�I!Ke���p~{�\��m.�a5�u	��#��|�3�e��V�����o�;$��Rc^�;n����F�_�;���f�ޞ��*P'���w��7�|�?�S+u�䛆X@6G�;�u��@����$����Gܷ�xR| �O�c�Q�}���?�)�u��=���ro�����Ը�tŉ�ot��\������Q���ޅr]h��UBLy�g�|n��bd�ή,ӻ�qq�      ��ϭO�U�^"~#��(������k�����d���ŗƠ���N��x\L����Yj�W�>��L�E��/�ݚp�����y�}�Lȓ�]�vk�Z�t5�*,�|a��u�v����(��.�Bg�D�����~�L.ʯq��ƽ.G�qt��:�G{j��6���|?N���|�m��v#*��8��G���B���s�g��iţ$_��{`��i�3Ը?�(���䡞��ݥ&�H�lU��+$_�EΞ]��~k>f/�\���wF��Be�w�x�g�kwgJ�7zn�tȉţ%_��	�t}��FO}��I�c$_��iQs����>�c_㟪�3���au�5]>�     2�%�.+��{'���1(��Sm�nY�wSξ~�
�z��U{��yG����Snw����W�
�У_�_޽M�2�4)2��t#������~�iR�ˏ��r3&n�߰�{�v���Ì��R�ߐ�1�?���ߖW��U�zq;��r;��e�/?�ץ�n/d����{��s��R�'�^�;aq;��r��5�K�??���u�G��_�k��O��JG���k���ϵ�}E�Wٷ'B��w�k�)�^�}����G�sm�/?�}Ӷ^U�T�^��0�_,��逇�W��������{=��=�.˛��m��XP����]j�.��${��]�G�ׯY0\F�H>x.� ���      e�mzH�s�Y)-xM�ݽ�����\���f̲��˹G�1�AM�ݽ�����/�"3tIꡞ�ёǋ׭�k�-���3�괳�)u�xݫ}{�C�B���!�y��W^��췫�O�|�kU�����z�$�P���R����S��O�A�z�Yj��k�����Rً���n�u^�ތ�7|z�I깣x�^��55�x������L>d����z(�>�}�v�L�ɞ�^����u�Bg������*{����"��j�Y�"d���:����~��<�}،�7���g��ξI�"��Ԝ����͵�.Y�#^����~��~E�;�^�䥯￨��t��ε�h����(      C�^���=��%�����^�={�ݫs�=��^��hp��s�s(����`�<���Ц�#
���eG�W�v�S��]y1X*�-;J��Ve�do�x�./�ط[.(�$^U��=�}�<�����������^ӟ}��~�x��}`�x�./<l��ý�}c�׾1�kvF��^����UzeA�J���k�g�y���)�U{����޸ץ��T��{:��}#���볧�5���Sū�J�zp�7����Zy��i�Uz�����%��j�D���NWy8{�j��u�k������ǈW��w��d���9���x�&V/��GT��p�m���m�K���q`�|����^����m��      �{��rޑg�B*���mن�bZfN���ܵ?o���wԙR�{�o�r��ݹ��0�+X/����;����o���{�$$��s��6H��л�wm�����{wK�Q �N�����s�g�^e?���w���ߧ朸��wC��m��P���qߚy:����j�/��<8�u�/�[$��9������w3��m�ޮ���~E_�ʾH�]�q���K��j�^�Re?\]c�ǃ7�v��~���o��{7�v��޻ٯ���{/��DD���n�kt��BO�Īw:��9ӫٷH���`�������^�wxѯ�σ7��٫������/�K<xk���=�\��_j�b)�+GL�	�q��s�<�=     @&����Ws�������mK�{E�\�y����U���	���W���nz@���U4}�y�g�~9�d�x�.�.����7�5;��N)4|rJ�X�
;��͞}#:���Z)��i�^�|��p	 I����֧�N���߈�j	 ��@�}��i�ƉW��q߱���?��b���njꈇ՜�ٳ���z�չ�@��R���}��g��˞�I�ϧ�� ^�/�?���/�z'{]��Ke�|�R�S���e���=�{=��T��j�y��n(�V��9�׌��=o�@���e=*������g�Bp���tS��\�{�g�b���^��I����9z�{�K�=��^�Q�ۗ������P��x�&}�կ�x={     �L�k�r�`�9RZ8���vwӫ�ߺ���|$�w�[��Sϗ���������Ty�K4��K��l�����zt��T����;z[\�-t ��
����*��D�e ��_�d�);��v�MF��.���ҩ�{/�!�'�W��z�T��?�iy��}����|�޾�o�t'X�I�9��sm�d��.�x!{}��z�G���?�e_�{&���v�����{j�qD���D�Ξs.>UsG͜�7Pޝ%ߤ'�vy�����z���e�S�w��6p�vO�M��mP�g\./?���_*{}c����j�Y֕?�뛚�1{%w�g�iپ�      ��;�#���\}�'��)���ӵ/���:qW�C��]���{���G�������pɀ����~C:�������s���m�p����M���To�̨\:�h��Qe�`�N��)�Bg�,\:|�k��n��q���2�e.��"��`���Y��鐚�/q��Ռ�F�U��i��DL�(�"~Ý�o	w�sN���.)�Wz�;\Q>յ�o�t�����2�>����Ӥ���}>gTٿ��Ng߫�s���w眳]e��g��w�:��}���#W�c��F;�]�5��yp���t�z��j�4{ue7�钿��g�z��������]�<�;�[��kR�G�#�qm����{�ּX�`��q��?���w���]��C{%h���.ξ^��������&>     �Lypۓr���c+����)��_O�W�x�o��(�k/�^-+�ʻ�:s��Qnw���Y�q� ��J�i�u�GG/�������Lo���m�Z��$�c=d������\�}�2�x>g�j�q_A�Y��o����#�,[�k���Q��h��������yY]Xy��ϚP���q��_6�����5�}����m�wZ�G�T�z���:^����[��_�ʞh�|���m}���	�cj�_P*n�w2z�ow^g�!�&Mq��}Sz���ܙ���:���������\����������8�u��'q��/$�l�7F7�k�,.n��5�$O��ۻ�     ��tGc����]�����/f@����Yf����5wm��erʸ㥼��r���f��;������ �u��W�>�d\η�+�<ڳKZ!�wv��*��U��s��.}��[�}������?cظ�o��[e��P�^�9Ӈ-�tA���^y�g�ɾ����q�+���5�c���.��q��g�������N���������'�/���&;�]���|�/���rV�Dd�;�}����xH�ؾA�7|��=순g���GԹv�P�>џ���'�9�r�SV����g�9�j���c�\�����s�����ט�C$�?v�q�����g��[��X��=џ��e��Rwd���s�C#��U��${��#�;��u�]G<,�w�쏒w���]�t���4�zf��ND��΍r���V�>�;e���#�Z��v      _m�n�ۖG�'�r�G��_hX%n⪂{G�K��'������nJ�6o�p�s��!��-re�4�������<���VJ�����)��ZU�SebaYֿ���WP^?��ξE�?b�L,�~�}v����7���9G~���~���տt�Ϩ����ո��^�{5�Q��qog�~�����D̄]|Hf��U�����_*���Z�T�Q+!�v����9��<�߃���W�A���{je]_�}�=*�^�����{�vE���?�8�N��E9�*���eM�y�e�D�־������9�Z��nYz�?�ƽ^M_�99�^���{w˫}{��󇊘e���U�m��ڣ�Fd�{��Zzܿ��<䲷����~�T�R42�߃���`��
5�����_cN��9�^�{z�Yi��C-���9G��Ss0����)���qo��)����2�xTֿ���:�`�$Ԍ     ���˦����)��r�	'� ��H���n����6���ҸV��N.�Y������{�����H�^e���;�*䂲��R����}M����~cv�ҫ���c�L+i�|�����ӫ*�f���.��B��
޷ul ��+�޶oΙ��ҩ����^y%�d�!=T�գ�j��tw��>e�d�z����J���ǎ�d�z�?���|?-�d����v�t���;:���{ʎ��+2�5��4�`:Գ�;���A���W��v��F�U�f�S�`0T�����D�9�W��s�f���s�]�e�_S��������fEp�}C�P�wN�k�9��G����k�LRٟ�����/���k�      H]�2eѺ?ˌI��H$����\��r��1�ϩj�m�uߎ���	.�p���Y����(�N(�߾�DbC�M%�Oߔ�-�i?�Dg''��b�߱��WS��Wk#��j;���]���w�����2��N���P���/X�/;�w�+�!��%��s�ij�9�d���]
%��n�-���Ͼ���Ԓqr���[�k�9Ge�F��^��b���o.8]���՜S�s6�ژ:ת�~��q��>�ξ\N����12��q_��}De&����un�o���}����ƺ�k�-*��o�z���45ߟ��wp��;�F{�v��Ͽ�/Sُ�H�uр���0��/����kg_�sn�K�}���:G��C���Jf�w�:}��~��٫��W-'�7ۗ�=�S��Ώ�{��㾝����^�x��������-�5��Md�&�����%��~w<`�B�o��Wgo���k��"ǎ��~��~�     8�!�G����KN����K�r{a�s���;�������F�,�����ۗI�OK$��;7(���*�z��;�$�S�7���Q�V�)i�t����/��<=��]8��]n�c��C�E	�xLe?�ξ?�T���k#ݲK�O�o����RُJ/{=�ձj�g��CK�9�v��Q�eS�G��p蒊~<��׹OKc���Q٥�}��~{Te� �CѻH���F��}���3R�C��:y�ݮƽ�Y���.��xo�=�u�S
Gʄ�Ҵ�ߡƽ��ppz	�x�Ge_L�ٔ���@�L).�i��쟁.�:{}�M^�w�ל8�=��z�r,����u��=��C�;x�Ǔj���g���o'��o��9����ƬSϯ����s�!�<�A�}�3٫���s��D�V��f5���S��}����'��}���^�!�Cӻ�<�u&{+n?����_�t��!��S���g?%y}og?<���\��|=�������iu�=������7��y��w��s�~-S��.�     Ș'v� '�4MFE�2�u(��k����[���5[�Ηdzٹ�s�r��ݷ�!y�q� ��W��Z��1%2�?LF�K�P�s��/%�5U�}Ԍ�o��'��Q.M��>�����~��~�!����t����镦���b)R��f�����񰴙d�����6����C�75:��j�oӸ��u���b_�����+�%��Vyw�Bd����.�m�o���u���"÷/���}�v�j�w���bojt�����-ُ�w��.��1��؛"��O��w�טd�*����D?��-٫y�H�>S��=�ߜ}����������)���T�9��|�k`�)T��9��P?�bÿ_���=�_�!;
�9P��u����}���ϵd�{7�h����e�r�P�(��=�G��٧(���#`F�M�Ogo�Vfg� :{��X���[r��u����>5��J����>�����U���O��#�e�1�}�     d�-o,��8C$��.0���k4ˍ�,��_q+�ܵ�Vɸ�+䔂c?6���{�a�ܽ�d�~�)��.�����ϝ���W=Ev���UO��l#��!��!�ܱ�Xi٥uv���gqج���U�����M�#��>w�czuw�@v��^��     �*n&d��?��~I�h��cSn��h����u�{��.�k�\ƾ�S2��p옔�oc�V�Zu�X˚               ��bA�����I3��J��/�������q;�ܵ�;�}A����>������ �|�f�%�               ���+��}L>1�J1��J��/n���/�"[�w�x��W��v�|넯HQԟ�q(�^c�Y~��|�oE                ��ԳC,|V>Xq�X���1(�^�2�+�Ț���(�k�
�w[o���Z�����)�^CO�����KW�G               �t�n�(~���*.�J��O����K�Ƶ�%�)�kq3!7�q�T�Y/;�ϣ�>x;:�d�s7I���              ����K_",w����+�Sn�H"*�z�Y롕ۓ<Up��J���)_<��2E&�ez��탧�oV�H(               �I��JO�W���Q1��C�����'�+�xa�li�!^乂{ҟv�C>|�t9��$I$<�)�ޓ�^�[��YfB               �L���;�9�~^$r���)�^s�U~�|�4�ū<[p��Z�Nh��7]�}�7�;��7����*l{J               �L��W[�ʜ?/���7�;�탷j�:�^u��A�2Oܵ�{�Im`��>���ۿG�}p��:�+j���               dK,��m�M>2�29��D����)a�r����M�i��u�/�k-}���ʌ�?-�V/'N��ke��?J0�'               @.,�}R�]+�����)��~��q��(�k13.7�)g�?I����6Jpp�N�e����xT,�                �6wl�y��j���c.�0�r�:Y��v	D��O�����e��y|�|�����.d`���zY����Y'               �[D1�Ys�<_�R*���U>Q�f�X�������]���B�yWp�z�A�e����q��8�32q�8�H(�e��C۟�b�v               �Ӧ�mr�?�O��a��_&���=�.�?߰R��ڽ��|��?������}�|�ԏȰ���`~������IW83               �G$�;��M����|�{'�#CՎ�:�mݽ��u�仼.�k	3!l{J^hxU>y���i�;8�6o�?o��=�               �i�m�߾\#���.�?�*���/����W�i�2��wg�[j��%��|������;����Z6�=�)�۶               �u��l�o?�K9����'}X�=U�Us�U���ay��%I�b{R�6����]��'{U���>��;�KyQ��}W���rߖ�ek�N               �ͪ=�ۏ��'<n��稳�g�vt�Ƀ۞���_r���!WpO�
��+�����������.���xs���`�<��y��iu	               ��6�m�cK+���-W�>��h�P<,�կ�g�V���n�ܓ���p��2�(�p�䂣ϕ�e���Ѡ�h\#ϫ���u��z;               0Դ�u�߶<"��xL�9��`�9r�QgJi�0q���5M�兆WeU�:	�#�~C�྿��F����y�?�؊)r������i�ض�1�,k�7������e�$̄                IX��nZo?
��YNw��>s�r������3�-k�6Ț���^�����A�謳������Ic�����ı��1���"aF������I��m������Z��               ��b�ؾ"�6�t��<�r�z�0�X�<�)�e�JmZ�4��;�.���;�,��}���e��쇦Ws?b��:r�L1Q&����ecd��2��\���q��/NO�W�C����&{{ۤQ���F���                ��־vy�^?^�����ˤ�2yđrd�_:��W����./.~�w���z �@�W��=Ң��7�f?t��g����QpO����1�l?��_hl��{����g-a%$�H�LHo4h                �fB�������aRRPd���0M	������X�=C(�g��Ҡ#�%                �I��5��5���;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;r+!��L               rϪ��� g(�#�
��b>�-               �=��
IL�	�+�                �@�                �
ܑ[�!>�X                ���++-��.<C               �{��m�^��+�                �@�                �
ܑSQ#&�w�               �^�Ę �D�93���&EEE�H$�               ������5�I ^��b"�
Z-?~��5J,˒��:�F�              ��+--�I�&����H��G�>r��;r�x�)S����v�0{%w
�               �QRR��c�h�4�4Y=>��;r��;rB�ۧv��ܮ��a	�              ���������b��W�I(�#7(�#�t�}Z�89j��������,K               ��x\���e���RXXh��.�-��nJ��:
�Ȫ}�����              �@��u�s����q�DZ��;���;��r;              �;Qr�[PpGVPn              p7J�p
��8��               �@��F�E�              �[(�#�(�#c(�              x%w�
wd�v               o��\���Qn              ��ܑm��(��               ���;���;S��r;              @>:d����1� N��G�����               ��%��z%wJ�pw��r;              ��@��F�i��              0�PrG&QpG�(�              M�ܑ)ܑ��               C%wdw�v               h���4
���               �%w8��;�v               %w8��;�v               
%w8��;��v               J�Hw�v               %w���;�r;               Rq����bH�tSr�AQp�Qn              @:Tr;v�H�Pr�AQpb
�G�����#+Fʔ�S���ΎzI������              ��C��[Z:�@�޴�������MҺ�u�?�(�ةł����PH�����KLYR��;,�>�r;               q��{�1"�`\F��.k[��M]W�)Z(��?$'�r;               �u��{AA�����(��?ttt����4����r;               Җ,��7N���7-�h������,               ��tɽ��I����                p
�                 W��                p
�                 W��                p
�                 W��                p
�                 W��                p
�                 W��                p
��)�eٿ             �C��|b��+ o���X4��H$v�              �.���~)**�� �N���%�P($}}}��             �t7/�����+����III�]~���D"(�             �A����z�`P�n��w���a������               ;tѽ��G�Ѩ�����;����{�m�L<�V�)ɧ �=�������0��cw�ؽً�Fw'�c�:-���v�,D~��G)S�K�P�*ԯ��Ñ���իWQUU          �w{{u]ǳgϢ,� �G�G���Jq{Z        ��I-_j�>��3����pD�&�v         �Cj�R����� �C�Gr}}��"         �|��󸺺���� O�G�4M��         �I��l6��h�a	��^�~]�         ����=}�4���Á�u�_�         �Wj���1�L�v{{         @�R�wyy�����Lo        �� p�����K��         �ߪ��F�����          NG]�w8 �;���         pZR�>�N8�;P�u         �����"         �E��%p           w           � p           w8QEQ�t:��h��         ���i���:��y�6pZ�pb.//��ӧ��ѣ(�2         �_j�6^�~?��C\]]p�p"��������-         �ii��'O����&����ț�N��g��ŋQE          �I�e��ķ�~�}�] ��C���~         ����~���d��/_�'�;d,Mn�        ��|���QUU�z�*���!S��8�?         �~�x�"�����}�4�8�;�&���2(         �~��/uz_�u y���F�A����ɓ'         ܍Ǐ�x<���?������;��E.-�.i         w'uz�=�W�^}r����;h2��b�u��o6�         p���zw8,�qp@)nO]UU���b         w/��������GE���Z�[        �����Lx�K������h�����u         �����ڲ,c:�pXw8�t����y�̺	�         ��>��]\\���������2noo�i����?�_~�e          w'�z2���8<�;�ӧO�/���n�X�|>wi         �#��Kۇ<y�$���Ñ���?~�ѳ�������         ���|���Oq{j�����Gt~~m�����/�.�/��)�         ��������G��l6�x�pd���QE�w]����ӟ�ԟ�Bx         `w��<���럽/u|)n����	�!1�L�~�'�������?�W_}�0         ����m���Y�7��ɓ'}���2���?����~ss��4����w��]<�<�={֟%         �����>^�|�S��z�4�6m�<ȇ�2��%N�Ybik��_L���?���_|џ)         ��׿�5����X,��ib�l6�[��,ȋ�2�����~Kܫ��o�%Q��c�}�]���m<��;{        ��.�M�eSw��������O���Ǐc2����/ߡ����~l1M�p�         ��;;;�7��          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,܁�k�6���ٖ�        ��*���i+���I�ܩ�����        ��Z�)xO�h4�wJ��U:�i�����-         �k��,mUU�4�]���;��UԾ
�        ���m�V��x<�{!p��PR�^׵�        �K=Y
�Ӗ���bw�m܁���=�         ������bѿ�B��d ����3�R؞6         Xg՜	݁M܁OZ��M���        �&���&��G��}u�         ��j�j��G�Q |�����m������5���m�>W����_         ܙiE���Ho���F���KS���eه���]w�gR؞Β۷��muS/P���ٻ          #)z�)|Ũ��{Y�/FOX��y���~+
#Q�7�@/,���=��~�6]N���I���O�        `��o�RM�Fl�|��~�z
�ǣ�>z�G����~�4w`E�D�4���}��iB{�T�m         �)DO/�KS��帏�ǣ�r��4���i���� <pij{
�w�um,�y�mݿ        �=�uo��VQe�˳��w������c:<p���@�����2��m���ET�"b���         ��4�jnc��&��8�L�,�����Ե��������������51��Ѵu         ��nQ-�q9��d��D�U�"�]&��I��.q{:+nQ��S�        �CR�޴U\ϫ����}�i�WK��t:��#p�$]�e��.N��:��M)         "MtO��l2��x��ǧ��$wxX��@�uUUm�q)h�]�D��q���y]�]�        ��+R(vǟ����:��$f�󍦹�&���}4p�	��H�۷�ۛ��*�z�����(�����;V;��        ��ū?%c�/w�VJĚ����&f���7KXW���?�;�s)nO�h�D:�mQϣZn{Q��R̞��U�>�<         �ܪ�z/�J�{�o�����q[]Ť����l�4��k[,b6�m48=w��V�&�ny𰸎�mv���)l_qX        pZ�����_}�^D���W�mߩͦ����<�ө��1�;�Sm�n�/n��u���x5��         �U���/��b��MW��m�ˍ&����~��=���ۡ��ϯ���u[XE�         �X1ꢟ���V�YM\߾���E�F�a�u� �������	�C�q�b˸��v        �mՏ�3Y��?����z>���F.�r����p�4M�/�C�M�}ܾ��xs��rˉ�         �+}S��Զ觬o4s��6�ܫ�Z~�b���i��=��HK�]���mu��'Jq{
ۋ         ��+�(�/]�E侸���e�e9�CR��-
A�w�G�B=TץK�\��&�pE�<vܐ�7go���������M�        ؏7]�f�y��u\�_��S��N�� ��;�u]�܇H��⪏�Kg��S�O+ O�Ĵm����C������         �e�"�k��������A��S;���X���d�R���n����fq{Qv'�~���ti��Mi��         �������������p�N�{���7a� �jMS��"N"n�x���/I        �q��m�T�$E��"����oj�&�I �M�'.���4͠}�f��׷��<Dd��QS���         d.��D���<F�Q�����>���<	�ᄥE>��6t�yu����<��>l�S�nZ;        ���4@�������A����t����	K����{��w];�W��3#l        xx���y�f����m�oe�3�S%p��.�2h�����o�ۋ�gv���Yn�h�G         ��TU��$F�Ѡ}Mq��%p������onq{:�U�/���        ������������M�'*�a6Ģ�G�*�!��+n��~        �4v5�}S��t	���u=hz{�gQ���b���+����V��         �H�[Q����������	�)��r	〡�p�Ң;D��>T�ɕX�&Mn/��        ��aHܞ�>Mg?;;[���N��NL:�,m��x�v�e�~�����~        ��Y,1�L�F�)p:ȇ�N����}���֗w�C�^�5"         ��M����rY8%�c����|�~E���#�],��V�        �0�Lq��i�'�m��̳u�z���������j���         ���!�z���V�e �A�'���a�5ՠ��>��E'n        `UU�ΞBx�;��;���Ȯ�vm4��>�m/������v         ���ƦI�Ś.MpN��N��v���G��)n?��x         r6$\O�����O�������Nľ�8�:���$         �qCc�4�}]���o4�?�;���i���u�r^�_��r���к���G        ���ں!���p:�p"�Lp��z؝#n_@tq;         ��"��x�v��d@��p���o�0��8������        ��	��!�&��'p�04poځ��[~Y݀�         6UUUL�ӵ��o42�r'p���[�O�okzz{��2         `SC����>���O�'`��f����L���r9         ��.Z_i�&��Og����8.�;��!g��]��������o6         �CC�u��4�!s�K��3�̲�-�]z1�        ���n�$��uv��	�!sC��n�{��\��        �ݬ�ۓ���'A���g6���        ��!܇Ngr_�q	�!sC�~��jM~3L�          ��&+p��	܁�3�        �C��� p�{aؙg��5˃��         ���p}�w�x!�i;t�=Dwވ�        ؟�q�	�p?��!I�]������         ��2P�wȟ��L&��M          �����4.�         ����^tm�C�         ����~�          ;��і          ��{љ�         �������          ��ؙ�         �}���          �]	܁�u          ;��3�         �=�;��w          �B����v          �D��X��         �>܁�t�v          �D��/܋          �]	܁��         ��܁���;          � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p8q��(&�I@Ҷm,�����Lz�@R�u��3�N�(��$��I?s>%=^��V��yt]��}ʲ�����$=^��f��x�o�4MUU��/��I?s I����Yg6��9&vl��noo����>���>���>���>���>6��>���>�1��> ��h�ĥ_Z��{V���+=f���d�_x��:�J��!1�5�w�5j�/�<nxא_x9&�}C~�3~��J:�Y����Yû�����}�1��ر��|��|��|�c�7��>�6���}lc����c'�2��> ��h          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�����:���&�o�h�qܴ��(�2          ��ڮ�y����]�g��=/o�QM�F��M����Yn�G��7���g�f1�j���}D�          ܙ����U������On�+��3.�;�v��ݳ�g�?����4q�u          �o��Z��?�ў���V��B;���o�X������DQ          쬝D\�KՋ2�C�|T�����v������4w          ��\D\�۸�����I�e?��(��F�         �Vڋ"^��(�i�'	�Y+� ��_�x�ߛ(�          ���I���3���A�$��.���l          ����Q4�����2��8���         ������E0����\�cg^��q         ��2��ˀM��Hw^���2��W�         �q���hg����;������          >j�����9�;k��<��          ���q�o�)�;[�>/b��          x_�������J�Y�&          �}�3�;�����2          ����lK��V�i          �uS�َ���tc?t          ��n��;�ѷ          {&p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p     �?{w�"�u�a���O�-am��I���&��%[aG�q ��5��U��	e2]U��u]�0�Z�N�u�     � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "��r�ݮ�i*h殅�fS}�4�8κ����ƜuӮ�n�7�9eݰF��}���7w-�=q�u�0�i�1�(�͹�X7�iΞؼ�}�}�1go�xF��ކ5�<��=ɺa)�>�-y�i�Ǎ�{b r	��r�˜/�,վ��B�R��`��rúa){ְ�a������a){ְnXÞ�5�mXʼ�5�mX�ކ5�� ��E�          @�;           �           D�          A�          @�;           �           D�������c�s�m���v�kk��h�a��rrrR]�4�^��9wi륭���nk��;���a_[/m�rttt��f��ƞ�}s�6���i��9��ކ7m6���X7�3�c�>�0�c�9�>s�����yk̝��˄�-׾�y�΍�/�� �P�m�8g(tvvVp��o��<�Q�kϨ9��uþ9/�ڞ�vn�{͜�M��x�žC�i�y<��7�^c��9�y���Xü�5����mx�yk�����y_���������\w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�         x'L�T@6�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D���T           ?*�;�t;�;          �놪I��
��tW          �ꮦ���`)�;��,          �UkM��	�Y��c         �m��M���	�,'pg���O          �9֚����Ŏ����m          ����t��;ŝe�,v��_�          p��'c���Q�w�/�u��j,          ���WS]~4�x�w���Ƚ�C��         �Cƪ��N��S�;�	ܙ�����          s�<��Q��Q_0���Y�S]|1          ,�ޟ���~W�{Nr�0�;��S���Xݮ          `�n[�-����5��ܹ���;�����=          �ѿ����z�Y�$w�$p�:�f��/'�         �k���χz�I_�G}�m����r�{��k��         ���U��i�͇S������i��'�;��������������         ��D;���ۡv�:��_^�/k,�3#p'uWSuߏ�}��ý����?�����׏k#n         �'֍UO�������r��骞�xZ�Ϫ~qR�}M�Nx���1'����ɫ��o\�����w��m�ق� �:���;�N:��{�﹀��ۘڻR������X�xF2ǉE������(�N ������/�z          pW���Gq�?�"�>뿖i��?Nc�O��C�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @� n�\�|>H]��o�XD۶)G��Xû�<��>~oxאu���zn3t-�az����UU�!�#��d��]C�)�7�o����x���؆���Ɛ��6�Ϲ��|������}�x8|w��'�N�ٔ'��t:�D>Q���M������Me̓lb6�l�Ŧ�۰������k��|�pN�6<��6<� ���          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"ܡp]׭ߩ�,�         x��JD��C�v���ʺ��        ����~�C�,��]NpwB         @��v"x(���.          �O���m��        �͘����
7x�ͭ��/����Z        ����!p��]t몎�[�;Z\M\ߡj��        ��u=h?!<�O���7�ƚ���}�~5=�V         �u�ږ�i�A��C��P�\Ls�����g���J�]�Ϸ0         Ґ(}�>C��wK�`P�^���ƬWy\W�        p7�Lp7���@^5ֶ��4�,���z�λ^;=         nǐ��&��a����*u�u��!|ty��Nr����l        `�2\������� �j���X.�ػ~��V         ��u]7(Jo�f��Lp�� p�0tQ5�X.���t����j��t�,         vb����h}��2���DF�m{�t�Q=�鐃u�Hw�K�ww         �l�w���p��@��.p���r��֔��n��^�?۰�y        ��t]7h�z�uC�����Á����q����Ի�j����'��q        `F�a)�)�@�p �����k��u��k��v��p         p�!S��x<t�����H^A�\^?����h�Q,�����?9m}��{sy�E�         ܪ��>$\7���H.����4㵁{�)�Y���´�򭫻��+�         �]C���l���/H]���f]w����h��ED�~�z���G��.:�;         �([�!��W�p8�p`rA^,�Og���b6�X�_�UQe��)���?����         p&�ɠp}H�E�fh�>O�Oq��~߷���Q1�         v-��܇����ÁɗKɭm��^]���I�3r_���	        P�M��j��_�}���F1����7�|9[?�=�b�j��5�lMq        `������x<tL���0	�� ��*�ք��˰��b6�X��Cu��E�y�nyy���o         \o����>d����p��p��
��S��y��r�A�7��w4x�w�N�         �\��1Id�P��5t�{����b~�����ݛm]z�i#�;*�        x�����W�u��I�,�0�����kF1Z�c�\?��j�{u��wQ� r��m�5�        �����;���p����Ex�\F۶k����b�.�����Oz_��!�q�L�        ��r{�C��e�Á��1�N��WWuON����*`�[FT;X�/�:�Q��/         ]�uQUÇ��?�:�	�����6�I��4u��Q����]���FT7�^����n��	        �=�M�>t"�h4�:�	���+Ά�)�e���>��˓����a��˟q�'7=         �h��=����󸦷�� p�{`�0��â���q\t�h�v�t]t�W]T7���?1�\k&p        ��rj{No*cx�~���D.�9�}H�^Wu�L���,�"������i�[��q����         �w]�m4�=��'''�oW׵���p�L&�����o�G�q>=��ׇj����D�[b�����8s��        �m�������������;�#��z6�ڿ��~���٫~:�`]ݛ��W��檦�̋�I�         ��6S��jr{Ndj<ou_@��p�4Mӿ��b������Q\��7���f�nyyR��[�ԣ<L��        �^�iܞ�P�o�?p�p�ݶm�1jFqR]E���ۼ�]E��o�W�(Tu��]A        p�Va��q����F��s��?��រL&1�N���!r����Q������{�t���I�         ���I�ۄ�)C���7�}p?	������(...6�M'��o"��vw�&t����ݫ|����nV��c�        ثm��w5M'''��������2	��[]�6��Or�_���qL���n���۩���3]t�U����d�F,���        p�ޟ־ٶe��)q;�w���
�4��6����8�j��<;��qy��!��yE����{;��r~0n��w�:         ؏�C�����X9�}նmr��x,n�@�@���n�F�f���q1{�v�����}���&x���/ߏr�{o��        �c�F���㻎�G�Qou܌�7���$p�b������d������Q,���.^G׶��Cv����&ku��y�yk�;        ���c"z�G���os�l��ZC�����k�NrO9ͽi�l~������Uy^R��-���-         7�q���эn/n��E�LF�y%�t:�h�{�.ߎ�'1Mb6��b�y(U�^u���        �d��۷�or;<\wx�VNrﶘ�^WMON.o{��t���s�;        @��M�m۰=e�~�c �K�T� ��q��<���VǨ����>]��v]��>�>t���s"        p2Dω��G�Q,������䞁{��ݖS�W�������"�<�[��?^�*t�"��Ƚ��        �[�!znM���xٳ��X����	ANt�N�[G�k�o�8�c�e��2ڮ��n�<����7�{����M�n�;        �Meg�ֳ9���<n���@��r����Q?�='���x�o�f�o)�������{w��������[��Jw���t�0�        `�l�V�S�}n��]�G�����x+O�%^2F��f;����f�Nt~��d�|����O�/?����w�F�U��v�e�;        �pd����6��|�����4��䞡�m�OS5        ���K���� F�|P�@����|>��b         ��U�~����&p�ʓ��2r��         ��F}�0��,O2r�        p��Ҟ���������V��r�|�        @]�o�v�m܁��	��$$��g�޶m         �pdԾ��LknJ���j�{�uoC���s         �WQ{���$pv*OT2t_y7xϏW         �a����p[���z?xO����	���"x        �ە}Wn�k�>^}}�����ػ�I���          x��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�ဴm]���      `�� �CTU�s8 w(T����<f�Y�-�          6���h4�������I��ɰ����q~~nR;         ��j�ln��5M'''���;P�;d:�Ư��*l        �[�\.�իW�0�'O����Q e�C�ʰ\(�0         `?r �˗/�I�?6�
 p�;�q��/��=         �/�f���GE]���;ܡ��+���b         ��ɖ/���?��$w�Cw�C���         
�M�˗/�I�����9??��l         @9�������4����X.�qvv         @y��;::��i�/�;܁W�^E�u         �'�l��={�~	�a��EL��          ʕ��r�4��L�{vqq         @���{��Q �#p�=3�         ���O�{�/U�         P�U��4M �!p�=���         �l��?w�#��        �h�`��G]�         p8��_w�#�         ���          �"�          (��          �"��@UU��$��q4M�         Y�u�\.c�X�t:�?�����i|��G��ѣ>l         ��m�x��U�|�2���8w8�����g���;         p�����ӧ�v~~ϟ?���� �&p�����UU         ��.���3�����駟(��
�׿���         �����>������?P&�;죏>�        �e��X,�ŋ�G���F�駟         �[9����,����}s�;�?wأM��ۛ�	         `���;���.���a�rA��ӧO         �O�<��.��k�3��K�{4���E�K�         ���N/{�/^\����K�{4��w||         ��:::Z������;�Q^�5�Lb6�]���I�         ����[��l���Q���^�w�!         ܾu����q �%p�=�����,ڶ��>��"         ��5��?���i����~	�a��j����x�����n�         v�^���d�w`��p2p������_�5>���          nO�zf4��;�w�#O�<����O�7��b:�zi         �%����������S����ᎌ��>r���_ϟ?����*         ������������w�n��;�/_Ҷm�����{����s�         v�իW���l�����;w�c�=��������}����wX��         ��M���������O��ۡ w(@�����/�\.�~=����7��_��        ��^�~�~�m��4MϞ=�;>���K�B�����O�����V��3x�����>��?�8��
         `�l�~���������y�㝞���6�!p�����ѣ~Z{^%vqq�v������ŋ����R         X�_~��1��i�yNj?::�[���(��
�f��e�>����������O?�kn����Y         ��Ξ��b��̞���_o�&�<y�ɤ�(��
�i��f�         �7��ٳg�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;PUU|���1��~����          ��z��i|��'q~~ϟ?x���?8==�Ǐ�������"          ��gϞ��������d/^�����%p���i�mu]�������         �ڻq{���X,�i��w	��'M�'���~��ˋ_�~:�8b1_ƿ����ꫯ�F�_~�e����          �~ܞa�7�|�����w-봞��u����"p`��g��?�����������[�V��E�          �gq{b�忖q�sz{?�۲�W������Y_>X��         ���q����9�;$r         `�v�%p�Z"w          6!n�&�%r         `q;7%pg�;          ���w[E���|_~���         ����]������Y��         ���[w6&r          =}�T��N	�ي�         �a˸��������������         �����r)ng'�܈�         �a�s��ܘ�         �a�P���?�vvB��N��         �7q;� pgg2r���E���#�/��������         ��#ng_������c=���E�UU���.r         8,�v�I�����W?��         �Љ��7�;�B�     ��o����*����m��%!��}a�����!�x	ۉ}�'�=�N&��so<���8��x��1ccC �`��KX$��RkCKkW/����c�Iݒ��T���s��U:oש���{~   7q;� p��tE[ra��         �8��)�;�*���P��         �(��)$�;�N�         P�������         ����4��7"w         �t��w�J�         �.�v�D�N�)r߼ys477          �oРA�vRE�NA�v�^WW�ܓ#�H�         �C���������I"���"�7ǘ1c���2<          �ǁ������[�l�}������j���ͱ~�����l6          ȏ�{��"�����쌶�ʀB�SP��1xpM          Px���P(w
�_g��<yr          Px�:WE���P�           ���          �T�SP---�x��          ����y���"p��:::b��}         @�e�C
I�          @*�          H�;�Y�	          
/;�2���Tgu&:&؆          ��          ���          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�          H��q1`X�0"F����cp߁1�Or�DUeU����{������f�@[c�?t0�6Ʈ�=��iWlol���ۑ�          �w������o��'��뀓&�oU�w�����ƶ�8��[�@���ݼ/��hl���I̱�wS&��1GŬSc�Ic��1qh]�?�iO��l{l޿-6����n�����=s?          �M��1%��49&��IC�ň'��u���{7����c�����aM�m�t����{��9qƨ�1g���g`��YUQ����	���Y[�=V�^�m[�-�u{7Fggg           �oe��;rF�9zn�6jV�8:7����7$��g^�˶Ɲ����`ےx}��hnk	ޝ��mN82�7?.�;+��AuEU�1-w|b�swu����xv�˱b���vf          �]��~q֘��q�s�y�����=�6��|Qtd;bю����W�-�`kc��x�
�u��h��q��b�I�"풻:��zI��ռ7���\<������          PN���� �+'_�=3�TVG�UVT�������xy�xt�ӹ	�_�y�>v����i��E��ݭQ���7��@\?��XtxS����b������          P��U��K'��zi�.FUUqnݙ�cG���'㑵OGc[S����g�������)Q���R�<��G���o�V=Onx!:��         @	�wPn��US����D�Y3<n9���q�����+�]�{�ܔU�>aH]|d�����Q���n��⣳�����y<��Y�;          E�u��f�%q�̫c@u�(U��n��q������Ǐ��K�i��,���㓧���͋L&�"����y7�5S/��-�'^߱<          ��TVT����ξ6����������&_�N��Mto�h�RWҁ{���a�5�W�.W�����}_�ݺ0�XxOlol          H�3FωϜ��;ht��~U}���|0��tA�����7���d�9���y7��f~��ǜ����,{0~����          H�dR�ͧ�^n�9o�0<�ù���(�񵻢�iw���ܓ;>}�G��IF&�	�*�d���~nݼ��Kߍ-�          �Źugƭg~"�����O��_5=�XxO<���(5%�O6!�x�gc̠Q��%�����Sܷ����G��4w          
(�|˩�ǵS/��U����O���ķ�0���RQ2��u�.�O�zCTVTG��fc���1�sRL?������Es{K          @��<&���[c��A�444D�=1�⟷<KVE)(�����*n�ws\:�{��}ժU��ؘ��r_g�������ڽ          ���1�ǟ��1���=Iܾq����쌦���%C��=k�bWԁ��~��K|>&t����.�����c~/�\<���          �ޔ�d��7n�����t�Ν;sq�okmm���s?������F�*��}T͈��}!�t�{��]��ĥΊ�)���          ������y���~'�dr��M���ϒV���o���[�k+���e�>i����Yn�;�s����7-3.�x���W�          p"���y���)#gݗ�����G}\gcG��S?�XwW�l�Ŧ��9�����\��tOw��.���Q�:$�l����ߙ�          �W� ������S��K���7v���-m�I7�w7���E1)��}�ɧƟ��ǹ�$�{z���A-���>_[�}�;          �%��������2lB�}ݝ��v����o�o��$�4m�bQ4���#gƟ�wkTWͯ\p��w�i�:��$w          8UU�X��3=���vm����?��-��E-�|�_��9q{������C���������{          z�"S_8���Q���;���o����N�X���ES{K�]���k�/ο-�U���D��]F��7N�:�]��          �����?�����x'��]gk6�8���_�'�;;"�R��S_���1���{z#nOtvvƜ�ɱe������          ���s>�N�,�5���2-���Y��ۗ}/�,��{E&����ƘA���魸�KGGG\;�}QpKl9�=          �\8�����k��;ѓ�߮�P�������FZ�6p�����s����KsSs�6���E߈C�          o7qH]���[����;;;{m��ܳ�'�i#f���#�R��[wf|p�A��+n�Ҳ�)>7����;          ~[��~�������ݓ���K[[[�0��X�ch�O��܇��ͻ%2�Lpt��ۻn���?/���|          @�?:�8y�Ƞ{�����>�k�6�?�������3/Q}O�*p��T�����ԧ&8�B�퉓O>9>3�c�d���Ѹ+          �ܱg��~'螮���6`���>yz\s�xx��&�
ܯ�rI�:rfpt���Ǎ#G�yW͟�����nOݝ          ���~������������ӧGeee|��b��e����H�����Ms?]Z�����q�������          ��g|<��	�.q{���:7��/~��"ۙ�4HM�~�OD��~���)n��So�W�X{[�          ���1���u�KK��e���q��㑵OE�"p?{��q�����1nO$w�$�����         ��RUQ�:�#�ѥ-n�r����^����߮��{nC�zCpdi�ۻ\6���]k��          ��w�_c��,�q{b`������~�V������ĘA������=Q���O�zC��S�          �ap�Aq�k�#Ks������/�<[l�B*h�ޯ�o\?���{+����)#gƩ��E;V          �/i��W��[1��ʊ��؜����)
������.�!}ﮘ��.7��p,z��          J۰~C��S.�[���]ί�?��ذwsJ��dz��_��b��3�O��G͎�ۗ          ���f�?�V�	�]��퉊LE�8�����R������Ǡ>5�;k���Cӯ�         ���U���I���.玝�kjc[��(���I��˂w*��=q��91i�X�wS          Pz��zI.r睊9nOTd2q������P��}��s���R��R�ۻ$oZ�|�         @iI諧\�S���].�x^���Es{K�[A�+&]�U)��Ɲ�[���lj          z���ƈ'oU*q{"������uOG��=p�h�?���7
��?>jkkO�y�M}�����u�          ���IoUȸ}ڴi'4n�r���#p�x¹��%�M��w�d�yw         �2����?��7
�WU�N>u؄�0dl���������qgo*�=1s���0<v6�
          �߹��Ee�"xS���]�7����5�1i踠���D&�������          ���u�7�zܞ����ђ"����7ΆN�C��圱��         J��>51�vfPq{b̠Q1~�ظk�K^�y�O�rWNq{b��7����          �8����L��r�ۻ�9zni�������S���[ܞH��N93���j          P�捞����ę'���z4o����R;#*+*�\�c��%�[G�         Pܒ&���cܞ�=bj����֎�����g9s��(W��'f��          �Q5#��C�\�kܞ������&Ʋ���Y/�d�)Q��=nO����ā��_          �߬�;캜��.�k��V�^���U��F���L&ӇO�W�X          ��'M�r$nӌ<��yy�u�O�>��QN��o5aH��         �HM:.ʍ��7�����Y'qs9)d�>nܸ��퉉C�          �'����!c�����jĀ�b`��8���}t�����92�h��;         @1�X�T�r!nw���e�{}��<�Q5�(����m��=�ܽ����         8>c��r!no�֖R�><J�����U���}žC�         ��1�Z�����FՌ��:y�
������3j��;         @��P�-pB�~t%�Wf*r��K������          ����v*n�|���~5��L&J���g�          �Rn@��ݗ�}���{��(E���ܷt��          J�����=���ׯʀ��Qj��Ǧ��         @��g@�q{���i�������R"n?v��         @q��(��H��Ǧ*���ׯNUeq� �F�~|J�f         �rPJ����%7:d2�^�v��gJcj����UW���;          堲�4z`q��I���Le�w���:�~�::;�؉�O��l��         �r�-�X�~bd;���F�����I�~�e{�n          N��"r,n?1�a�%��eۢX��O�֎��          媽����O��<u�~Ś�Z���O���C         @qi.�x׮]��(_��ׯځփQl��c�         �r��Ё(6I�^__/n?����������fq{���R|on          ��@k����!n��H�ޞm�ƶ���i'n�]�	�         ��ޖ�Q,��g_����fh�wq{��Ѵ+          (.;������;�N^�⎦��8�.�J���:���yO          P\�aȱ����h��>�˕�v0?��������ol�<�a          p��l�4��G�nt���ܸk���=6��          �7n��l{TW�/�����}��N^�h}��LO2n?~|���F9��         ���llڷ5&i"nϟ����yo^��S�%��7NE&i nϿ4��          @���ߒ��]ܞ_�8�:/W���-8O:.
M�^�v�          �Ӫ]��	�F���oŮ�y[+oWwyÚ�����hhڝ;          (N�w��4���Rܯ�zI���p��         ��ٸok4�5ǀ����텑\����m��]��;W�\&��|�֢�+         �����ҝ��1�d}q{�������zy��{[�����b��O���[�}i          P�^۶� �����^ݶ8����j'�s>wq{�mط9�v          �-	��M�^x�~��z�_ܲ ��yu^�����[_          ���Ɔ���C�򲞸���6Ɗ]k�f^�����c[��]ӻ�==���r          P���j^�B��5551}������|�;�y]3�<��^��.nO�-�E��-         @ix�����9��5����\�]�=pz�K��������/          �c[��X�{}L;iR��_ܞ���ƒ�+�n��d���]�b���'����t�����          J˯�?�+���=]_�ld��Z$��']��	�������bw��          ��<�����i��U�N�9��钼�v]����Û������<�s�����k�          JOs{K�z�q��KN�������ű�qgA�.H�~��5~����Ȭk��<��tڰos��}Y          P�X�h���Q���y���t��G�vA��ë�~U���>��/nO��W>��7          �g{cC��eA�[w�1�CܞNk��ǒ�+�~��}��ǯ�?�zi����=�v4�g7�          ���V�<~g��9�)�����w��]�`�{��?��']}+�t������D{�=          (mɤ.�E�=!nO��״�
��i��\�d|p���z��=ݶ�Om>�X�  xIDAT|1          (?^�/q��Ӣ"ӽh\ܞn?Z�@�_��+h���w��㒉���>��8q{�ݹ��xC         �?�m�'6<�O�ਏ��ۢ���7��(|�~��1�^�@�љ7��c���hǊ�׭�          �凋��͋����1���ӦM�E2��{iP��=�躧��S��Խ�����ב��.�;          (?�폟,{(>uڍ���������_��A*���l|�;�]��Q���������+~�o          �Ӄ��ǟS�Mx����鷧e_�h�����wo���<�M�<����8l=�=�]�p          P����_��q�e�)*+*s?��|�hlk��HM���k��1o�)1��V�^���l�7��l{          P�6��?]���Ȭk��E��/�K[D��*poi?���Oq뤏�=n�d21a>|x�=?Y�P,oX          ����c��IѾ�%�k'q�ԩS����д;����H�T{����U11F�u�q�Ɖ�{`�uqﲇ          �d;����_�rK�4�/r7��g:�N�������%���^}���?����|$A2�}ĈA��;�?���?�66          ������P��qՠs������3���~�觱�au�Q*�������ߏ�8����ګk��{&{����KwDCӞ          �w�¶���a3bdǐ^]�+n�����-�տ��Je��hlm���>qud{�΍L&�Ǐ������/          8�﮸'�jέ���;S���=�a�������H�V��+�������<��_Dq{�=���xh��          G�љ������M��hoi;��������_��z4��D��:pO<����礘[=儜���c�|���          �][��ό�>���O�9��=���_~���iw�]����6�*M��	���\���[�cy��߉l�?�          �t�t���Ѷ���#wq{ϵv��y��~�(E�'~����m��cxǐc��&�����W��f�eO�3          ������Ϫ��4:�;�����k�h��<��X�sU��	��Z}w��bLg�#uq{�-kX_~����P          ��X�kytd;���+z���{���%��ߎ�ۖF1)��=q���⦉��䊱�z�����mK�>���G          ���xϪhjo���\m݋���=��e|����{��]���kÃq�؋���#�������u���W~���          �i큍����I���ܫ��{n{cC��O-�8�#�QQoy2v���(�Z�9e�������{�?�,{0�5          �-��k�/��tDӻ���܆}��o����ݼ7�U�v��Z�3o���Co��q�Ɖ�{���9��ʝ���W          z[c[s|eٷ�Of"���D6���]��s�l���֫?�涖(fE�'�l�//�V|~�'�Sun�x2����6螵{��o_�N�~          ũ#����θj�Eq��3�P�!q{�e����W?����DkG[|u�w��)&\�#�����'���7t��k          ���Ƨc������c�xq{wm9�-��ߎ�}��T�D���k/�X_<�31e؄�5�5�7^�3���j          @���[_z�����ک�F&�	�ۓ�/Ʒ_�+��[���T��H�B��%��zI�4��ѯ�o�V/o}=���G�д;           -ڲ�q����_����u�N�jO˾��w������xp�������y7ǩ#g���XxO���          ��Zְ:�����Gf_�qUTW�d��#���xd�S����;�ښ�T��+����n��FΊϜ��7�<��h�h�W?�-�y�}          �)��~ג��uO�'�~8�7���d2Q��Xw�~Olػ9J]I�]^߱<��ؗ�I������G9��v�c��{�?���          �&�`��_�G�=7��P̩��bݞ�q���孋�\�E��h�h���<�Z�L\=�����+cX�!Q�ڳ��T�Kqc���          �nY����'�����}]I��k���\��uatvvF9)���ˡ�ָգ���_�E�ώߝvEL26J����ܝ)�y"v7�          (5�v��S�M�͸*έ����(vIȾ`�Ҹ壇���(We�wI&�?����1���r�E���D���Ql�;4�����/EK��          �R�fO}��߉���eϏ+&_�kj���i�Olx>[�l�qpG����[���Ww.�/�{F\P7?N5;*+*#�6���mz%�����         @��۲?~��񳕏ĬS㼺yq~��\��V[��-�ͯƢ�ˢ�3�I��[�ښ��������i�fǼ�O�3F�)�o˶ǒ+�mK��m�c��          �)ۙ��;W�;�8f�g��g>&����~�o�ۖ�ko,����=�����=hm�MGO�L&u�F���5bZL6!����7yC��X�wS�ص6V4��ջ��"w          �Ȳ����aM�k�����3GL��çƌ�c���zKs[K����v�{��ص&7i���wC���i����u��~VUQ㇌��A'Ǩ�1�fx��?,��rx���}F���w=_����s/����bG��r`[����          ��K�_��uQ��2���?�.F�Z��&xh���8�����;Ε���s=pr����Z��M;c㾭��iW�q����%	�n���q$Օ�ѷ�O��lG4��          PX���掣��[;ZmA�����Û��F         ����/�;           � p           �           ���          �T�          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�9���Nw#�    IEND�B`�PK
     t$v[�Ƚׇ  �  /   images/ce527fa2-4558-4370-a5e7-21077342728a.png�PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK
     t$v[�c��f  �f  /   images/cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     t$v[��EM  M  /   images/48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     t$v[������  ��  /   images/27b84e47-6648-4cee-a869-6ff1a6fc12fe.png�PNG

   IHDR  �  R   ���P   	pHYs  H_  H_#�
{   tEXtSoftware www.inkscape.org��<    IDATx���yx�y&�������7 ���)�(j�6[�6Ӣe��H^�ǎ3��s�L�sg�vnf�8�d2I�+�"�Z���H�i9�lI�H�%�;A�@��ݵtm�	��H�]]������1��h6��s��	�낈������*K�t DDDDDDD���������*0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
�* Q#۴i�"BD��� !˲� "�PHq'!B�q��(������+��A� 
������EQ4]�5EQ�[��0B�P�u]˶����ի�`��DDD�a�u+Q�{���'��8�u�	��LEq��M��6	���I���}���q_B�u�!A�Ar]w����s�(�'A�w���U��+4Q�c�NDDt�>�l�$Im��L���s�;�q�ɂ L0ܕf�w]��(�']�=��c��p�u�c��{o��aU/&�DD��^z饴asA�#�\�ug�$� f �W8�zS p�Q�u��`�$I��ٷjժ�ʆGDDT9LЉ���;�P�� �ug� s����o�� ����_�}���$��������Z��#""
t""�===r*����"�q���b �H��w�u�] zEQ��7�n���������LЉ��&���SLӼV�� ���{� 3���Ƙ��� �%I�[�(�u�]w��t`DDD�b�NDDU��g��-I�
 #��r �*U�S� ��- oٶ���{�=P須��.�	:U�g�y&)��2�qV�p���X鸨.d]�}�+� l�e��;�c��A�`�NDD�$����\׽�uݕ n� �XḨ18 v��_����=��Ӌ��扈��t""3===R*�Zp.!��� ��t\D�v]�uA^�	&�jŊf��""�������y�搦i�����V �J�ET�! �.�ˎ�\(�loo�+�'&�DD�^xa��8w���������<� �o~8������.i�uݟxQ�W�Z���Q�`�NDDey�Z��8��\׽K�Y���.�yz��j������b	�H�߀���u_��?���{3����jt""*�s�=w� �X�z R�C
̥�l~~^���H�mA~�8�&Q���'>���Qma�NDD���'�L&?�� ����1�e�s����:?iYy������
��)�����o�+U7&�DDtQ�<�̤p8|ή��	@�pHe9?I�X�.��^�	|A����
�����OW: ""�>LЉ�h���??M�ϸ�� �����$��M�����M�m � �m�O�^��x�""�������=��s3 �/B;���L��d���8���n��O~�{*Ut"����x��8�AX��J�s%�O���EW�FWڷ�h�v��ի�T:""[LЉ�ĳ�>�,��\��� w��W���=?���O֫=ia��8?�B�<�ND���ձ͛7't]��u�� ��tL��q��Ye7]��7 �P��ﾻP逈�(LЉ���7���ꫯ��eY_N$נʪ����8?��ڌ$�U��\�}R�G��_���_����C���V0A'"�O?��"�0�a��b��&M�(���+�T�ޟ�WSҞ��2�㼒L&���{��Y�x���|LЉ�j��͛�gΜ�=�0~�0���OO�ӈ���m$)��՛jXaw]}}}p]�  ���D"��?���~����FDDea�NDT��zꩻu]��b�x�i���U.�2Ə?&11!�FT�d]�4d2�|_�$'��
��졇�ɘEDDec�NDT#6mڤ
����/��9�J߿'N��P���p�oY�g	х��N�`�e�L4̈́��d2��U�V��	:Q�{�'�/����i�9�S��d2�d2�K,#��@#��ju�q���]�$�	�ÿ�D"��C��k0DD�+&�DDUh��͡����d���>���jI�0i�$��u��|~&�\�\���H$rZ��oO�8�oo��v��`���WLЉ���/�В�f�i���bԯyǏY����3)'
�H�����ӧaY����p،D"�&�����'?y���DD(&�DDU����V۶��0�,����j<G:���g4��(ue�X,�̙3�]_�$W��-�X�wx���|����<a�NDT9��?���}�0���^H�����$�+�D���D�R	���TU�ڑH�t$���z�; ��@DTLЉ��XOO�,�_��[��'����͈�bLʉj��V�]�ũS�/�(�rA��E�����@/FDD`�ND4FzzzҎ���akMӼ��>E�dѨo�ډh���n��ڡPȌF�=�ƍ��w�ygv�.LD����lӦMS��w���i��X^[�e(�Y���LD��,�B����uC���F�L&���O~��^����0A'"
ȳ�>�$���O]�o�m{̲�P(�X,�h4�J4U/�u��:4M�i�cv�s��H$�~�}���5&�DD>{���o�u�_�X2Vﱂ �&��pxL�ID�gY4M��끟M!���.I���v��_��E��t""�<��S+
��w�X6Vﭲ,#�!�p;Qs�b���٪���{B�Я����E�����'��V���u}�X���k��x<�P(��������k�6&�έ���(������ Qc�ND�ѦM�������i���Z*�"EA,��r"�P���0
ض��έ����֭{3��!&�DD%z������k�v�X��r;��0���b1���#g�����O��o~A"�:����
=��S3UU��a�8�h�,��h�7nc'"�ضMӠ�j����%�[EY{�����bDDu�	:чx��'���C]�?t�4Q���"���8t]����oEэD"?7n�g���@/FDT㘠]���?��r��4틖eIA^+
AQD�Qnc'�1�.��"��<,�
�Z�PȎ�b��d�˫V�2�Q�b�NDt7n�C]���4�h��	�B�+�DD�4RP.�6m�p��(��=��C_�Q"��0A'":Ϗ~��v]���0��A^G�e��qȲ�e��Jf�&TU���^'�b��noo�a�""�!LЉ� ����0M�S��yA�/F�Q(��p8�5���`�6
�t]��ܹBr�#�Ⱥ|��و��1A'����3�L)
ݚ���(��Qͱ,k��{PA��(�(���}��w*�U9&�DԐ��o�.��B���	,k�F�H&�L̉��9��B� M�[Q�$ɎF�������׿�u'��U1&�D�p���?S,�[,���F4E<gs"�;c�����\$�͵k�n�DDU�	:5�'�xb�aOh��,������hW6"��9��iZ ���H$��������r"�*������͛C�O���B�𥠶���5*۶�����.I��(ʏ�����?���t"�k���_6�ۦi*A��s"���N���p!��փ>��@.@DT��Q]���iYֳ�a,
b~Y��H$�bND�>�e!�ˡX,�>���� ���>����*�	:����������Alg�$	��@QY�'"��a ����m��E�Q�׮]�;�ONDTALЉ�n����T,��u}��s���x<�X,A�����.��]ב���8�wM�ey �L>t���o�}r"�
`�ND5���WޱcG����	�=-�#�31'"��q��
UU}o�&E��$I�joo��<�a�ND5����aM���4͘�s�b1$	�b �߉|%IA��8��T��u]��y������pX���_|��7�>9�a�ND5���'mY�&M�n��},
!�N#
�:/�刢�H$Y�!�2"���0dY�$I�B��=8�m��², @�X�eY0M�i�~mt]�i�c��$\!9A��~�8��Gyd��ɉ�� t"�96l��i~۶m��yEQD"�@,��b<ѨH$�X,EQ��FU�#�m��u�a@Ӵ��Ț�qE�c���}��B�b4�Ok׮�G_'&"
t"�O>��B��c�0��s�s+.�����N�iǗH$�J���!IR��*�뺣�z�P@.�C>���15.�qP(����v477߹jժ~�''"
 t"�	7n�u]׿c�����,#�J�\�D�)����	�t�d���˵j8��|>���a�r9�J�KP��%I2E��5k�����	:U��}�{�X,�cUUo�s^I��L&�D���L8M���tþ�\�E.�C&����
�B�C���:r�����A@4}�����U�V�l:U-&�DT���5�|���eE��S��q(�¶i�I4EKKZZZ�L&�:��4��d088�L&���T����|��yeY�B���֯_�����	:U�-[�������w_�p8�T*���T�X,�q��aܸq�����ض���A`hh��$�eaxx��.����lٲ{-Z��~z"�21A'�����u�a�۲��_s
��D"EQ����$I?~<&N��d2Y�p�eYD?��l�á�ir����1dY�F������ܷI������������M�qǷ=ÑH�d�E����d2�	&`	�� ]���ߏӧO�0�J�C5�u]C�u����D"y���6)Q��Q�����2��aL�kN�4�RH��I�&���Ѩo%�
���L&���>U:�A��e�x8�uݺu�|����&�DTQ===_QU�X�����h4�d2��O�P�h�&M¤I�X��
躎�'O�ԩS<�N�D�tI��X,�;k׮���MJDT"&�DT�7o�<y�9M����}(
!�J!�2կT*�)S�����Uث�i����C__�������Eöm_��,�\Uջ����GDc�	:�����kt]�I�Xl�kNEQXȋ>T*����ӑJ�*
]�q��ׇ�Ǐ3Q�Kr]�B�B��9eY�B_�~��&%"�LЉhLmܸ�
�?wǗ��("�J!��1թt:�����O�]ׅa�u}�u]�i��,���gY\�E(� ���("
!�@��~)��X,V��A��ɓ'q��	&�tI~�����(��k���/]&�D4&}��h8~I��[��3�"���աj]1w�|~tկP( ��C�4_�H]�H$2��'	$�I$	Ȳ<�\�mۣ���P��M�D"ۛ��n^�z��]t"
\GG��e�d��/{йjN&�bƌ7n\�C��PU�l�l��þ�s�H��t:���&���hYhY�9�S�N����4��@6����
���d����g��2!�%0A'�@uww�����կ-�H�t����$I´i�0y��n�VU���`ݬ���ojjBKKZZZ*��k��C�!��T,�^�� ����7]E'�}uݺu��eB"��`�NDA;;;��4�S~�ό$�kN#&M������T�wgΜA?}K��(�hjj¸q�0~�x$���144��BӴ�\����i����S�P(���v���	:����k�eY�4c���a455U}!+�EQ0gΜ1��oY���q��i�9s�}��b1���b�ĉc~��q?~Ǐ�}�m�F�X�e>Y�O���׭[wԗ	���a�ND����y@U�n˲|Yƌ��[���&�"���0eʔ1;��8p��q0�EQ0i�$�����ϰ�iؿ?�����TF�A��y_�$�L&�k|���|���LЉ�G������:�Sv�$IR�T�U���N�1g�D��1�^.�É'�����
\#I�Ә:u*Z[[�����S�p���9�O��� P��׭[�{>�FD�������#�ş��Bm�rt5T���"�"fΜ�������8�h�����^#�$	���hkk�#	�b{��E6��ZT[����0��e�h4�KY�?����'xDT&�DT���������4Ͳ�Y	��x<�x<�GhTgE��y�}�E?~ǎk�bo���Ԅ�ӧc�ĉ�Q8u�<�#	������P��3�$�����!4"jPLЉȳ���{u]Ҷ�ϛK��t:]�
�T�A��)S���h�@UUq��A���1�C��`���:uj����B{���]�j�i��f��ly�$ɌF��[��YB#����<����sM��o?ΛG"�R)Vi��Ø?~��UUŁ�����*y#�2f͚�iӦ�^���C����3]E7�������ChD�`��Q�:::�4�3�����t9�T
���lWE�PM��YX=dY����1cƌ����~�߿�;%����.b��s�ׯ�קЈ�A0A'�+����G��u}i�s�J;]��ɓ1s��@�&�E�۷'N�`b^Ţ�(�Ν����@^���w�a�� ˲044�˖�h4�N:�^�z�j�� �+����HOO�t]׷�Ų��ɲ�T*�*���$aΜ9?~��s;��Ç�СCl�UC��$�ϟ���f��m��������sSms�l֗���pxP���֭;T~dDTчڸq㝚�=kYV��݊��I{%�=�H.��(��}��I�۷���5lҤI�7o^ Gb�9�cǎ�>/�6�uQ(P(ʞ+
c�ؽk֬yɇЈ��1A'������MUU��8NY�AA@*�B4�+4�#�x.�����6f���Q1k�,̜9����gΜ�޽{y�>�0d�ٲ_�(��D�?���ۧЈ�1A'�K����UU�\�<�$���	�Pȏ���455a����ypǎþ}�|9GJ�%�Lb�H�Ӿ�;<<�w�}�i�:/�>۶��d�~?����u����O�Q�a�ND��������;[���Q.�͢���|޷9������6̝;�ׇ;��a���<A�.��,�({�H$���~�����&�Dt���+���0�%���ǑH$���Ќ30u�T��s��C��M��(��%K����n�&v��Ue�m��|>�˹�H$�}����}��_g�J"���F=��M�Ph�aegM�t����fϞ���V���4;w���АosR�3g���ٳ}ۭcYv�ލ\.��|T_t]G6�-{�H$r<�H,������ED ���9�ڨm/�M��#�"�����
�� �;w.&L��ۜǎÞ={x֜�N��d��:ض�ݻwcxxؗ��������!8�S�<�px8
-����0&�D����|>�s˲"��#I����ߜ.JE̛7�ƍ�e>۶��ۋ��>_�� I/^�I�&�2��8سg}���m��e��K]�$#�����u�B#�����uww߭����e�Ub=� �N�Z��(��?>���}�OUUl۶͗s�T�f͚�9s����8�}�]d2"�z��f�.,(I��(�k֬��>�ED5�	:Q��������+�ǹ�(H$L��A��y�0~�x_�����Ν;�^�����܌����,�=��8����vw�(�uQ(�~h(����~cݺu��ShDTc��5����?�4�o�y�d�X��Ȩ�̛7Ϸ3�{��šC�|��C4�5�\�d2Y�\#�*X8�.EӴ����*��׭[�w>�ED5�	:Q�����B����!���|Y���5s�LL�2��yFV/O�<�CT�h$I�ҥK}yPd�6v����tI�b�l���q�  �s�ڵe}VQ�a�N�`�������o���J�t%��s^,�}�v�P����`ڴie�e�&v��	M�|���eY*����(��~��_��/    IDAT�),"�LЉHgg�UU�l9s�R;]���V̞=��yTU�֭[��of̘������yt]��o��4}����8�#I߰~���>���v0A'j���O���@9s��a455A˪)Gu���,(�h`>��֭[a�O��5y�d,^�ؗ��Ν;��M��u]d2���(������W�U1&�D����9M�V�3ۨѕPK�.-{����0�n���I
̄	p��W���qpp��.x?E��.��l�c��O~��;|
�������\WW�K�&��hMMML��dY��N�3��l�����ߏ�۷�����҂3f�գ����v<�4��=��/|
���WЉꗰaÆWu]_Y�$�x�D¯��N����K�"��5��� �m��-�4f���q�ז����~�:uʧ��^����; D���y�}
���WЉꓰaÆ7�MΓ�$�s�"s��);9�eE���Lo��Vٯ�Y�f���>T"�@2�,k]�oذa��B"�*�����=��[���(g�t:EQ����Xkkk���s��z뭲�y188�;v�u�\E̟?��'�C)�R��1]ׯ}�Ƕ�U	&�Du����U�0��3G:�F4�+$�c�D3g�,k�|>�-[���,�"򠿿o��vYIz$�UW]�z���(�j�򎎎7}��� t�:�aÆW4M+k[{SS�s�"�p���/�쮦i,GU�ԩSx�wʚ#�N���ͧ������k������U�"�
c�NT':::~����^�����D"?â:6o޼�^/�ib�֭(�>FET�cǎ�СCe�1m�4��i���D���T���������B"�
c�NT:;;�i�G��ió�t�&O�\�M��8رcTU�1*"�ݻ'O�,k�y���=���,�hnn.k%]UՏwtt���aQ�0A'�qO��z��� ����,��1EQ�����ۋ��A�""�_oo/���<��es���1"�g#Iz�G�����x�ǰ����հ���nM�>�u�(�hii�*]1Q1o޼�n"���_��$Q�����ۡi��9ZZZ��p@�#���������cXD4Ƙ�ը�����P(��:^�$��� 
�չ������������>FD�b���۷��#}���,�IW,
�����$�����Q��"�����uvv�wM�~��xI����I�|���]2�Ĕ)S<��4;w��1"���r9�޽��xI�0w�\#�z7� ��$]U�/tvv���a�a�NTc����HӴ��:^E&�T2A0{�l�E�F�±�9բ'N�رc�ǧR)L�8�ǈ������AWW�W}��� t�����EUU�庮��#�ڙ�S��N�Z�����^��m�0M�_�mW:�������1c�}PI�H�5M�����/�L�z�ODc�����B���m۞>�EQd+5�$�b���W�O�8�]�v�U��m�\�\�B��B�uh��4Q,/{6:C�eD"D"����_MMM�����(X�r�燜���ػw��QQ��,�L�s-Q�x<��5k�<�shD &�D5�G?����|�e۶=�
���p���ŋ�N�=��4���/���C���\.���d2�P( ���D���MMMH��|�w�N��E�y_n�6jL�i"��x~OEщ�bw�[�n����ߘ�U�'�|ra6��n۶�;�>��&/&L��y��y�.�|�M&#�`�&���p��i�>}�a�4^���, �pg�^tḀf���.ƍ���VL�2���4��,[���r]ױm۶�*�Sc*��f��_;�P��J��>��{|��|����=������b���2��9�CE,_��H���`���>GU�L�ĉ'p��q���_v5,*��,��E��f-)鸈椈X�×?r�@^sP�\d.���qj����6
��?�S�&O��ɓ'�����߷^ɲ��+Wz��8|�0�?�sT�������dr�<p��Ј�'LЉ�ԦM�����æi��2~� ϙ�Wmmmhkk�4vxxo��W	qv'A?�=�'N\��۸����$�laz��I�<��"����q䔅c�m>eúD}�T*�ٳg����E&�?~<�/_�i�m�غu+L��9*j�bCCC�������X,6���]�94"��U'1���`rN�"�2�N��i�����m��ܶm=z�h�oI�Na�0�ja\jl��K��qͼ�;l���a�Z�=dB=o�}xx۶mî]���ֆY�f!�L�i���̙3���Ckkk�c%IB[[8@dT�dYF:��||�4�	�(n0��Ȉ�\A'�B6l�w]�o�:>�N#��5�y��a	��>|{�4�G�4q��A�۷�b��&���!\�@��Y!�".���v\<ac�A[���.�W�Ǐ����R�(+O�e�t�M������۷CU� "�F`FY5>b��O~��;|��|����tuu�s�P�u���$�;QY��.]ꩭ��ix����m�طo������<��X�D���h��rY��m�L�����}V����X�hQî��S�=��`���>GD�DUU�r9��E�����{�� "�1A'�"���R(��?��D�x�稨�,X����[o��3g��Q�;|�0v��]�/����>zM��!$U�jy)���xeGo�5aZ�O	���ӧc��{��Css���;w���+���Q(<�O&��f͚��1$"*t�*����|>���8���c�R���aQ����X�l������ضm��U�L&�m۶!��^��i$�}C�f�-�V)9�ŋo�xmW��$	s������!���S��D+W����$��b׮]DE�dxx���(���(��]�v��a�LЉ���O>�pxxx�eY�
7F�Q�R)O7�D�[�p���@�q��k�5�yZ�4�{�����,�ޛ"X<�>���:x��:��3q��D<�5�\㹎A-Z�`��\E'?�0OcC���(ʲ���^��"�1A'��6�l�>j����oY�������V��y#�;s��n�z��%*��#�ui�p<j�O��!��p��̙3�x�b�B��4F�e�r�-���\E'�d2����R�p8
�f<�����"���'&Qu���59�BH��L��ӧO�4�X,����>GS}���ݻ�w����b���n�"k���#�l�l�����C��	�p����uq��A�����CSSS��T�XġC�0w�ܒǦ�i�R)��S���42�,���?�>�i&A�`���ITA\A'������k��/c%IBKKKC�����z��;���ѣ>GT]4M�믿�L潅�椈���0z�=�>x��O��=d"p��2n�:%*@7\<�_���^E,]��fͪ`��E7�|3b�X�c��������T>۶��d<wӈF��y䑏�]!&�D�aÆ��u�w���ƍ�$I~�Ej�ܹ�8qb��t]�+��ǩ�Ŗ��~�����\~���n�!Zz��������GO�hI��m����d����u��Ɵj�Pokkòe��z���ɓ�d�Oc�m��0u(X�e!��x~o����Y�n��{"*t�
����\.���ן���&D"���F�q�u�y:*�{�n;v,�������c�����a~4��4Nfn��[{��ɖ"Ngl����,�*I��k&��x��T�;��v���f�x�uێM�|��P�䱧N�������Q�X�`�O�����֬Y�!�`�N4ƞ~��E�Lf�m۞���ɤ�?�K�1c�N�Z�8M��ꫯ����Ν;�o߾ѯ�7I��U1L�;W����w��.fM��+"X8#TR�z��M���2F+�+���+W�mkH����`˖-0M���0��4�sm�P(dE�ѫ׮]��簈�2���������i'L��T-)�#�H�50Q�b�
�����������DUY��`�֭��?=��"�[�s��Wwxy����̜\ރ���Lt������w��a�t�Mhii�#�R�*��#G�zW
��\.���,�YMӦ|�+_���1R�����P�X|�kr�F����&L��)9�u'O� ��ro��&N�81���h�=V�����b��_�2a;.��'�c+d����c`��0��"��l9Յi�x�W�r�ʺ�>R�~���%�mmm������K2���8�u���b1�H$^���Ȉ�b��N4F���-
_�26�������wW_}��?{��šC����l��믿�S�N�~��"���<+=�x�����uO᐀�q����<��:�_O00|�h�(�X�r��"��L�z뭞���ݻ���DE��u]d2��'E������ߨ��b�������/
��y�y�$	��ͬ�N�S�\sM��l���/���n�r]o����}A >uK��~����*-p���Z�-���_Opr�l�P(��+Wb���_{,͜9���+y[�Q�i�&��W֬Y�/�FD�a�N����\.��KQ8Q���\�-��rf͚�ɓ'�<����سgO U��x뭷p�� g���o��֫�SB��҂��\���|/I���[����PU
�B��G>R�V�u�u��Z����mx:B!I��D�]�~�� B#�s��DQe���?������S��s
�(��V+]׭�V�w�M���7�_rn�.�|�����㻛
�,`��1��g�ȲȘ'� ��	�����|��Ѳ,���k�4m�c	�eY�j5�Pw��:H��t:�i�m�R�X|yӦMl%C &�D�b�詏P2�d�s
LKK���pgΜ�\��7���E��k���N/�xy����A�/i�G|iu�.�����<hIE�W�S�>w��0���ku�f���?���3�T="��碳�e����f#"��1A'
HGG�3c����h���)P^���S[���l۶m������č�Q.��x�u��0��w�&��%��Ʊhfi}̃֜���qD�Ac˖-��?�B%��F�u�'�*/�{^�u�����o����( 6l��0���26
!�L��(I�<��5gΜ	 ����:^���s�s����㱪J\��:x�������Kf����	|i����[hr�x��G]�����;�S��s~۾Rp�;�����1:�0�h�ƍw��	:��}��&۶�q��[}A�N�!�{�e����O��z��<��|� WsRį�RPˍ����|Q�7���^7-����%����o}̃�pF�V�����;�\�򮖝>}�S׃���פ@555y�<�m[�u�駞z�~�:U	V�"�Y8~M�uO����4��Q�no�R��ٳgt'@H��Uʘ���[��y}d�Z����=mc���gзlق;��q8����>L�6��q�p�T
�l6�Ȩ�I��T*�����ǚ��������GFԸ�LG�����u}���,
Gc!
y����d�8\&���(���E�6�6V�G�.�{�·{����y����mQ��瓸�h�&���wk>����ۓb�xA��Z�u���q�|���B���4mAWW�w|���1A'�Iww�ݪ�~���H$¢p4&���=mg���Ǝ�`˖-p �xV7-�+Օi���9|wSf�JBT����G?y�$>\�ʗ�fQ(J���@4D����b��j�������9$�����===i]ן�r�<{�IJT����Ǹ�[	��ﾋ|>�l{�5�v3:���*-��UZ�O�p�u�=<ٵk��b#򇗟#Y�=�n�"�Jy:f�8�`�S�>�(ϣ���]�|P,�ݲ����G�±�A<Uo�d25��r9�ݻw���|4�D���r��Wwxy�����U2f�6�G��E����6��"�~�m�X���a����Ә={v��ZZZF.)�N{jh�f,�np��A5�������ot]_�el*��T˥���$�IO�#}}}D3�v��1��}�����pD�v�Vi4�*�1�s �D��0�A��ѣ5��/��y������^� ���˺����琈t�2<���k��'^��b1D�Q�C"�$/7��뢿�?�h���ӧG�rX���W���ci��g�Ka�]1L��Vi~k�$����ܹsg�񇗟�x<�p�z*Q}�F��G�Ӟ�����BTaLЉ<ڲeKXU���;�BH&�A�EtI^Ο�r�����.z{{G���2M����;x��w7�����x爉;���k_H���bH'�{�X�č﵍#G*QyN�>]�A�J������rG�u��͛77�v"��ȣ�{�n2��g�0ϝ�X
�B�:�����Ǐ����Eܾ�:Z�.������q䔍q)��-������p�XD�]�G��/4 ��ݻ1m�4O��A6�E�X�,��A���`"/F�U�nIc��bs__ߓ >LtD��6?݈*�����B�੥ϝS%�R)O�j9Aw]�w����룈E*����U�e�m����Z�19��[��w�7��i5���.2�L��x�ƚ$I�w��������a�C"jLЉJ���Ӣ������F�<wN�M�i� ��q�СѾ�M	�,�\��Vi��[��_k�U��D�s�{����3Z��yY	�F��D�c5�X,��<��0�{/��BK a�5nq'*�i�?�,��$I�x��*��kopp�䭍��u]�߿��{n� T��+ê��v���"��{�U�u��*�O+���Y����ѣ�1cF���dpp�Ӹd2	�0|�����$LӄeY%��,+200�o �&2���t�lܸ�5M������f�;��E��6E/�p�ř3gF�F�"V,�
�g�l<�����Vi3��*�O�(����@:�L��4�S��x<@4D�'�鴧{M�Vtuu�q a�-&�DW���c�����2��Ω�����l6@4c������i��m!i���y�������b~I�����pM�H���T)�P��Q) �u��;::f�Q��c|�+�8�Om�.�;�x�'J�/�n�e!��M�TUE__��g�W.�����6~��@�!���;���#�"/JWoB���x�ͳۼ��ߏ���W8*o��,�M�VҘ��m�z�j��((�%��m[r�g j�L
��
:�����{�0J�`񺵘�O^�����M:4�����W��.�{��ߘ�w��Ԡ�O��׾��=7T�b|��e�{;"N�:U�g��`E�S�D"���iO-Ø����_���0A'�O?��"M�~��Xnm�j�%A��������ã_�r��U�GZ�}󱳭�l����R*.��g�W���c�*�7�B�m�<��6c"?��୪�����}��!�nq'��|�Ƕm��0+��%U� �V�ju{������	s����L/�x}w?�b ���59�O���!���غa��݇�V�>r��̙S�J�.������\�8��J9��iZI��M�|��NtYLЉ.����[����:.
qk;U�X,�@�H�Zs�����/���G��Z��u}�'qwL�,����.��,
�BMV8�f�%'���N��k�5�0�wvv�����PhD5�[܉.���g��i�e��v$D~�r3o�f�+#�b�8 ,�S^k���J��'��
��
�$`�����8q���x��AWЩ���]��?}�'X՝���Nt	�b�%/U��B!�hQu�r3_���#+� Д1u��$�X��_l+b�"䰀�������	>Ӯ&Kg���;&��;'�͛W�J��g-�@�$O�׉���H$J~;�#��<���DFTۘE]�ƍ���z�OwC�PMn����FKS�����޾xV���k�U���83d"�:�,@<W��q]�u��hJ��,C��/~?̟�P4]d2���p��]cMUU��[�h4:�0���E�a0M��q��]����g���PhD5�	:�����LUU�/J'������3/�
UU �����}��+K�\�}���*�    IDAT��q��Ƹ��O��M�媫�nZ.�4�W�T*�	��cV2v.9���e\��BUu����Ɣ�2&4�~,�CfM����뢿�S�L�tX%�m�����EQ&�TA@:����@ɭ9��7~��<����x@��$&�D�cY֏�lm���l�FU���Z<nY�h_i9̝z��7�v�m���0p&�`�x��a�U�����q\�?f��d̝�M)��J9l�q���(1J�SZ�������a̚Es�~����x���"U���gۭ��s�!TM$IB</y��m�R(z��`"#�MLЉ�������.)u\8fe]�:�(z��[�+��l�s6Q�:A�x���#��~���aթ�ViC9N�X�p	��Ӏk��UQ1c�8̘҄=���D��!V�_�D�w300P�H����&���ꃢ(�u�KU�������nݺ�Q�a�Nt��øm��.u�H%SVm�j������u=�h�5444���I�h�x����~�T���M�\N��G�O\5k<�s��:�%W%����%Zǉ���ٞ�e�\�N�0J�t�6�ou/U�X��͛7o����k�Ç( ��)F I��(�%�����!���e�M��ѕ�Z��dF~�}f�ƿ�]�k;M�p�|��;��`bsuWd?t�D(6�,�����r��\�h2�����	Ģ����0m����Ϯ�a�����4^�q���H��R�#������p0�Ֆ�C!#]]]7�~w��X�������z\���M�p��F���!�7v��iI��$�������iR�W-X�5dY��ŭص/Ӫ�2�6��l6[�H�a�N��뢅������)���j��� X������d2�h����&��V9��4��s������T<i#����(nZ"#*���Ἅ��ĵW/)��y��a��O��=g�|Q:�ki��v �b�@/[���0DQ���.T߼nuw]�b�G �Q��e�1����-�0&�:NQ�bPU�����,TZ.�=�m�.�����/$�k#5��;����m\��1�f,B��8����#Z[/A��!T���.�u}�ƍ�2���j
tjh�<��$]����q�$!�H�o�lq����`/��?����2BRm$�#�4q���c�xM�����	�����pޑ�ZL��)��5�����ֳ������??!���jtjh�B�i˲J�a�v�^�b�@$�:� ���RU�K�0��"�G0�urE�?wF+��S������t�4a����c,NJ�l��M�L�=@HD5�	:5����5M���q�h�[۩&��j~����i�����v씉��W���x�f�)��[���g��]��?��{x�y/��}���@	�`c��'���[����69��wڤ�i�&=mOJ��Mz���yzڜ��\��� L쐘�Nm'����K ik�ٳgf����X3ڳמ�����S;�5�I[��z׻.�~�7+�LЩ؅�aW�}���[6o�|�!��?�d�� ������pB6�#�p���q�q��ḋ�� ΍h�={��f���7�

 ����u��ILЩT%�IW��L�{�C�LЩ,=����fg:�L&]%=D*�K�>�,�"�ݴ$"�J jc��C߀��@"z��ΏU ܃N��m��0f>���_� $���L���Ν;�����:�ż��n����ON����Z8�C�������<�l���"�N�����e1�E<wU��f?�u��jB"*j�t��s���-�e9�\***��|����U��܄|X�;��1�qA�'���6t�'�N�[�C���큦i�2����CTԘ�SYټy�M�L�V�������%?��O.���-��Hɱ��h i�y��j�����K&7��$��B�f�w>��c�=��h1A����fr��g�S�����,���j�hʕ�A͗�k�rU?~���	:���>>�e	]׹�Ne�8��
`˖-��f���~�***،��F�$�NLNT�xLXQE,�,�)�&e�LЉ���i�<t]_�y��{QQ�ߓ��6m�2���v���p�g������BJKZlY����L��ߟ߿��JY,C(r4FJ�L&��>ꂨ@��SY��k�&��V:WY�xQ�(�}r�������@&�Q @�-D���������\:���Q��#���5*LЩ䵷�'���g��s󖗨����׍���d���Q��!�a  r�}I�5��M�k���M����M�'
!�:�����?��	�<&�T�,���i��2m!��W!-?�A��"-��_�RS������R��9��'}�ݜ�����;?��@4.�L:��2M3��QHDE�ObD<��c2���N�%	_��M6�����c���,��=b�\��0p~�@u���[ I_,��㑘n~߰ĝ�, �;��d�iooo� $����JZ6��l۶�W������ATl�<��q�qr����t ��sM���p�'��z6�L���nJgU�t*G�D����m��4��{QQ`�N%���)�ɬr:���������
���'-����4�k8��^e󛦄e����X0����G"����r�%��wBWǮe2��nݺƃ����?M�m��vs���.�����s)��ǣA�s�u]���Nc�VY��3~�wS���Q���b��H)�N���QHD�1A���e˖꺾��87MK��U��A��б��W����_(�����Ce�_�]��c���2~ܞ�i��c�\΃h�
�ͱk��/ݼy��C����J��@��s�z�F}��B�N�$�~l�5�D��?K� 	 ����<o^A津ěG�|��dU��<i�'/gq��D<r�O�p�RLJ�t*�p�H�lv�c��0�_��.2"5��N%����׳��\����`Gt%nV���`+�N�@��0r�,s�yt�~�2���`n�`�?H	8a��S���Q�l�{k�,��R���G$�-o�9�TJ\���lٲ�W=�H����L�P6���.�xܗ{o���0�c���!&3)����]E��#ؿ��t�7�`F����⮚0-���4�����:Fa��=�/|"�����gR�DUU��H�qS���s*5�@���)%t]�'�B"R�	:������d��:'c�v%*vnt�n󨩩���S=�݇ �X�(�}��������nK��7{��4��ݐ��kY|�;#xhWq�nK��?Z�떄��J�O�^�z�1A���p����J��g1]��l���x�2\2����f���x<��pT����
�|� ̘1G� ��6���	�]�����3K�^�||J���8ԍ�s��.ҕ�ᴍ����k�����B�cmͳo�v(ecpxl=��I��]U�"/�b1d2G����_�o�"*<&�T2}��?�f��N�!|�@G4�\RJ�/��Ѩ/�qGϚ���{7M,����A<�󟣥eM0G�����X\�`���r��[x�u���ABbUk�.���w.�;�}q�|�̙�|���wt*U�u�Q��0�7o����|�#��ahD��JF6��_N�$	hwzP��f����%�I���x�7b���$R�R����o_q����ą����'��f��mlD<q���Җ�L�lW?`[�?7�d��������2		�xm�[AU��?����"i�̙^��7+�n�c��`|�dtt�ѸL&�% LЩ$0A����#�|�0G�{�zN� ��8N��z�A]]R� ��i�dt  �Ί`�,`85�cG�gh!D" �e"����LacfUWϏ"(����]~�'�'rH��X�{VD�L-V)�7N\\A����*T�!X�N��D�L�=����aT?��#���G?�C#*&�T����1�dҗ�DNd2�K�M����Ǐ ��0��U�lx�n*�AT&/��6-����mK¡0�(���Ro�4�ԋ:��Y�Y���[��qi!�e��z,�����/�X��b��Hb�N�l|e���T��	 t�=&��{�7o��a�Z�j��jՂ�o�6�������#��,�4��H$c��.�H�
�0��g�W���X��c�ǰzq��/���.��766�)��rӵڲ,��� r*�#�N;]E�����[7n����y�	:�ޅ}G�p��ʅ�=�C�4GF� �����ݰ%����믹�>m�֨.���,��k �K�o�C�ᚖ�?~8q�,�ٳgO�~*TTT8�N�=����!�H$�C1�+ �����;�ږ-[��a�:q��ʉ��y!��ġL^I�s��9��Fll}6�/{?�e-�����$>��D^���6z���G"�K������3�ͳ��*�9n��z�c�=��DDT\A'_�d2_v:Ư���i"��!r��\UU���!���Ncc#����4q��������|](]v�l��������¨��o	�/\|�2{�l�VDq�蝹]E�d2_�mO�"* >��o����o������!)��QD��͊�nce� ����&����.��H��Na��n^Ɵ<P����{rnZ�������޿P��� 8n�E�g.W�6o޼ѣ��<�t�-�0�^J�h��S9Auu��1N�/&MMM8}�4���d�����{���xG�����x�����Qi�]E��&��aT�쯪�����NOW  )���D~�v=��~@�7Qy�	:���͛o�u���M�\�V����X,�P(��n�uuuH&�H�R�x�h��b��|�m��C�y9��A{ZG����׳�>�|��󊛗`��ò�w�����b1���:j\�����{�}�Ї��04"O0A'_2��8�ǹzNe�mIluu5�������X�p!^{�5 ���e����[�J�S��QiN��p�g,A�Bhjj*��p���t���==���#���DE��A'�y��ǯ�u}��1Bvn�������q~-������p��.#蝌�O�B�_~{O<��:���m	��G��nI�s xn������f|�w!�:}xx؃h��_,s�Ȓ�f�m۶m�G!y�+��;�L�N�����LT�FFFo����U�X������СC ����u�󄨜����W�xq���\=/�;�F�4KMR�{��+�.n�X�`��8򡦦�UEWЩ\i��x<�驔�t��|��Ȉ��ʶm�f�q��1\='r�`�H$|ݷ������{裝���*�Tt�x�G|�{#x~_���G��ħ��ʒs ����»ٹs�"�H(�e�jkk���rlGe-�H8~����m=���8"���N���d�ɲ,G���xܷe�D�r��yW�jjj��Օ�h
#c���8|�0 `��Y|��A�����=Y�q2�HH��ea�u�	���,�rh�h5!�,Y�8��q��s�����^t'��ei���=����(����%��ݻw���Nƌ��;]ב�f��·p�H�ɫ�'�M�z�x��EJ��	��%�olI�t��;�F�g�Q��n�Er O<�O��755�ڿ],�񸫪.�?'r��7��~t���\�$��7+�F���r9G��F�Q�='�`hh��������A�4G���H$�ŋc��� �Vѯ]*�q`��mG�U��vӵ�����	�/4�����G4=n_z�;w.ϑ�����N�{�r�p���w��3�l6�Y�c�zNt��А�1�@����`�+��Fl��S���	��,���<�+�@@�c����OT�=+�/97r[v�A�����=E�����u��ω.p�l��f���y�	:���͛��u�QK�p8<Q�JD���;]u/6��a�ҋ'3�d���V�ULG�9��u�}���8Z[[G4=�p����nv�JQ0D8쨠���>���yQ^1{!_�f�_s:��~�����J��߭���N�7,&hhh@WWlx�'i|��	�53͓����3%���k#hV؍}�N�Xxn��cՖ/_���������Wc�Nt�x<�pV����
�Vo""�������޾8��.v2&8~�JT'�P555�(��X�b������p��_���u�=F�J�l<�r��A`ek�������sFN�?ve`]�7g�̞=[qT�7k�,�cl�v�=���E"�A��ԏ��f�K:::������ahD�����i��p�r��s����y��kll�}��F�t�R��� ���^2/���z�Qi7-�QiN<��s���+V(�h�ܖ���,""�x<��t)%R���X�]TD����Tv���oG��������IDo��:���q�����ȶ����� `��*�����}�?G�Mի�sxa����U�V�DE��ٳ]��x���9��0�;������B%�_����D��?�,�QV��\=�7��@�Uyn1Z�r%"� ``���(?n��m�7��C)|�c#i�{o��O?Y���"��GОA���b�����Di;0V��m۾�\!����\.(��#�B"�&�T�L������|X���n�b�D�v�ډ��7N���/�����lN�g�e�����>*m�2Y�o�L#�{[R]]�e˖)�*?���PQQ�x�����%*7ne����!�&�T�6o�|�a�N�D�ђ(�%���訫2�����yV[[�k��f����_�Q�磧2cG�}�;#x�Y5�8*m*l����=7v�Z(��%��͙3��8��]Y ����*�0f?���xѴ�I-�4��9\�$D^���EKK��qMMM8t�P�R���CCC8}�4�}&�꤆EM���qp���^��QiS!%о;�C��V��X�vm�4������,o'��X,]ק|�����{���Ƚ�x5M%���=���:'cB�B��W!����>W�ϙ3���TV�Z��ڱB����8�U��l<�����)<�/��B���+��x�$� ��y�8p�za��娯�WQ~566������g�v�)�Î�����������%*&�T���iY���O��M].�ùs���%�;�aݺu���V�(:�me1��4����;��M�B��OV�cw�|s��T��Eϼ|q���E�0�|��_SS��q===y���t9}�,K�4�yѴ��oz*�a����y��s�����577��I	�p7�t��^&+�/[S8�W�������汣���ZcG�}���CE�t����|1���br���rI_�RPWW�T_�uG�;��h4������
t*:�=���aT;�惙�ܝ?�\��x<>Q^*b�n�喉}������}��e]zTڨ�{k�Ɋ���"���&%���:v���Ѧ�&�\���>��͛�j�ۗgD�J�x�&���x�'n�($"ט�S��f���pD޳m�u"�6�(f�D��r��牞���)8��c�ƏJ���ƎJ^8*�O����wcY��?�৯\\9ojj��իF半�
���8'�dy;��x���RJ�����7��'�4	"��Ν;#�����iN��4
aƌ^�ET���0֬Y�j��^r����e2���?G*� h���(޿��Q>���H���,��k �K�o��k"����:�{a���#g.��hii�ʕ+F�+V�jv700��zQ�tT�u��ů���>g��
WЩ�����p�Ɣ�.2�����.\�0����r���* �-������L��K��a[���+���~�E�� >��I|�É�Hλm�c{������+F坊�
ם�;;;�Q�p�,.�o߾�y�+��T@�b�槜\�i"��j����N���9WSS�����\E�F����[��K/��� ��~gz-<xW3+��~�k����r8!���!ܱ.�ڪ�y?��X�8=;�rL�	    IDATC�4,[��亵O������FFF�Q��F�H�R��đ��~�׽�����S�زeˢ���CN�'�����HD�޲e�\�,bϞ=DTl�ƾ}�p�ر��-����/|�sw�wY�ɞ,�8�C$$���>�&Z���߉aO<���/V���a\w�u%u��[UTT��np5�����sDD�%�Jattt��k��������w�	�"�:��S�0M�+lG�FWW��}ƌ%���=�-_�555x��WaYҺ�wv����0�5�hx,�x㤉]/�8�m�2�Ꮅ�wE�$��_��?�Q}�/�bUWW���/��m��纮cpp0����h4�(A�m�l�/ <�]TDS����a�\
��[�(��d\%O�/Ƌ/��R��jjjBUU^z饉����C�s���2Y�ݯ�=ga�� >v{��
A+�Jv c��������/|;!��҂e˖A+񿐚�W�E���d��3DT(�`�`�9�8����S�`�;���mppp��1���%�CTHuuuX�h������/��V�ea���8~��ے��uܹ.�kZB(�㼧��c9<�s#W�#�V�^�Y�f)��0�����]U��r9�ٳ�ѾY"zg�t�Q?!fΜ�+��{�S�E4%��*�|C��/8�^��pDy��ߏL&�jlkk+�=�{�@ ��˗��o|�	݃Nv[�������>��X
�~2}Ir>w�\|�(�� ]�D9}�4�s�<�F����R"����G�9�tR���=��d�\.7�z�h4:q��tVя;��G��9��e�&<��G�^�\%c�������KxN���]/x���ɏ�X+W�,��{qs��7�zq��s"o�?�lv���A3�G7n�hyѻ*�G�`0�)'�9���(MM?���\��͛7����W��&b�ҥhjj¾}���� He$:�S��W��uy�/��T���}�y9�W��.I�� -Z�E��E5�d,p]�u��&�D�F��t�4��m�7�����1A'�t]�]'׳���;RJ�>}��*z ��%K��+�xY񪬬�M7݄��^�߿CCC ���/f��KY�X���"hi�g�j����xn���g/m��i���p��W����d2���fWc��,zzz�c=0���/���0A'�X�NJutt����Fl۞r?�X,���J/�"*{˗/G2�t5���_Gwww�#�)%�����oNt{�lN] 7]��!ģſ��=h�ox�`��KWy��;w.�,Y�D"�(B�����P]]�j��Ç��ח稈h��𰣪.M��%K�$o����(���tR*�J}�Ir�����?�e˖��x�b ���9��'�@cc#��ۋcǎ]��l���g2x�:�7�t~K�1��xz�vX�{4��Gs�x{�u0DSSZ[[�617w�\��y*�B�#"�ɢѨ�ݶm��ٳ��u�"�2&褔m�8�> {]022���A̘1���p8�E����D����������(N�8��'O�0 c%�GΘ8r���3X:?���4nu}(%q��ġ�&��a(u�ʺd2���̛7�P�`��h4���V��O�8�sω<�ݜ��)0A'�X�N��ر����o���)?�&	�e�D�L4�ʕ+�i�Vw_y��Nb�6Μ9��gϢ����i�5#�9ug�P��*�I���>q7-�％�s6z-��p�����;?��a466�����˚R�j�*��ֺ;00���9""����Q�R�)_�Y���뮷�S"* ���2������`y;Q!麎��n466��5���^�X5.w��������0M������BOO�%G�+3�� �&�j�*���dL �A�`��@��I������1����X,�ٳg�������_Д���f�ɹm�8y�d�#"�w�F%�e�t:�Y _�.*�w���1�ל\�[���N�>���ZW[K"����j���kD�o�`pb��m�D__p���˖c�600lc` �wLo,CMMjkkQ__�*�w�L&]�r0������1""��@ �P(�/�a�	:)�wR�駟Ntvv�8YA���D,�2,"��3f`ɒ%���߿���y���ٶ�T*���!add�t����:/;#����������@uu5?W�4�֭CEE����W^��s�sS����Ry�m�M}Q�p9��8���9-ogs8"5]7��%K�����H��y��4i����JTVV�����_6�E6��a�f�0MRʉ����m�+F�P�H�h�Hy����:9�#G�09'R �8.s���� _�.*���okR²,G��C���W�ѻ8v����\��\�/��",+���(� ���,���a޼y�����`x�=��T�&餛{.��$�����B�s�ΈaW9�R"����S�\�O$��k�Q���q\{���r�i����9m4���<����D��
.�N��i����������=��ٳg��d��؍W�Lg���c�5�"��s�,iY�8{���(�w��
.������ٽ��8H)q�ȑi��_u�U����cTD�Z�t)���񽽽�cDD䆛��e�D��
���=���չr���x躎cǎ��iV�X����.ĬY�\��uǏ�cDD4.�ܯݴi�%*(~�Q�}�4MG]��~����������z|8ƪU�&:��ٳgc����K)q��Q6F$*"N}r�\pٲem�CtYLЩ�L������ �ۉ�бcǐ�f]�O$X�b4��������`�ҥӺ�ٳg144����(ܔ�g�Y�C����i��\��s��d�&><�3�kjj�ٝ�N<��ˣ��a�>}:�QQ���aG�[�u�G�]t*����kr�\���?'*^����>:����/�SDD��F�z��im���r8t�д^^�w�.�d���-[�,�(��a�N#����MӸG��ȝ={v������p��<ED�N8ƚ5k���PJ�C��0�<FFD�
� �p4�4��z��0A��1M�W�\��s"8r�2�̴�`�̟??O93�����i���ɓ�wN�.�D��Q(Do��
�駟N�1���{��H˲p��Aض=��������)OQMM(��ի�L:ځ�6����STD�%�	�a�O?�t£p�.��
"�J}ʲ,G�DLЉ�#�N�e��%K��ܜ����l|弢�bZ���Ç�y�E�81<<�)��!�t*�0~����P��/���� N�<9��,^����y����+97o��ƴ+H��p��9��r��e��bDa�J'�s�9�?uvv���{���?>-Z�����.�bݺu�.k�,o�������gM�4Wx
�%����x�kL�t�y���D�u��q�;wn��iii��%Kw�%��D"��k�N�[;p�c���h�"#�Br��iFb۶m,�"�1A'����FT>��T*5�{555aŊy���݌3�n�:�� _N�^D��P���t:��<
�ht�i�w8����D�7^��N��}���:�]�6/I����F�Z�
�`p��:u�T^�r�ZNWѥ�wy
�&��M�6i�i::ܘ	:Qi��r8p� t]���***�nݺi7���p�B,]�4/�GϜ9�3g��!*"R�i�����}W�)&��U�V}�4�)�	!�������䥉V$�ڵkQ__��Ȩ�A�X�,������p�ԩ�܋��s��=�y��[<
� t�����`0ȆPD%F�u�۷�\n��
X�b-Z��
��D"�u����NOO�?��{Qq���X��_<
� t�i���2����4麎����%I�:��Y��7tY�f����_�D"�������رcy���GL�|�G�`�Nڽ{w�0�9N��y�t:��_�l6/�����7܀����܏�O�4,^�˗/�[����N=zNN#!"�p������G��g���g���n�,k��c�NT�t]�޽{��������x��4 #�J&�X�n����vϳg��ĉy����-��4M��G�1A'�ض����C�����\.����ctt4o�lnn���_�.�eʋ���ӧq��ɼݏ����in��}£p����wr�����N?�ȿƓ�����s�
*_���X,�5k�䵂BJ��G�����y�?�=�LӼɣP����g�eY��������������/o�߃����&�@ss3n��F̘1#o��,o��&zzz�vO"*~.���硓G���'6o�|�������#۶q��ἯVVTT�����ŋ��,��CEE֭[����aؿ?Ν;��{�?8}5M3��c�q�<����	˲>���p8̒T�2v��i躎��Ty|����D^�Kj�A,X���-���x�7`F^�KD�0ި��g�a� �sr��<aY����,o'���>d�Y,^�8�5�x�V���� :�T*��{����;w.,X�����~9r�m���D�Nt۶��a8TƘ��'L�tt��ۉ �����k�᪫�Beee^�=s�L�p����ơC��Z�3f���ŋ�L&�~o)%N�:��g����D�?.��x
�9!�T��;v,���>:�����c�;MB`����={�'�7M�N��ɓ'a��'s�{UUUX�p!fΜ���s�<��S��ߤ������B̜9���{���W\A���5'��A&�Dt	)%�;������K7�����	�N�©S������*,X� �����1<<��"��y6���`pʿ��0�� ����Q�a�NygY��N���s"z'}}}H�R�ꪫ�H$�~�P(�����'O�ę3g��)P]]�x�b�=L�9sgΜ���rB������e}L�)Ϙ�S�Y�u���y]I&��޽{1w�\̝;ד��P(���V,X� ===8~�8FGG�>]$�@mm-����z���躎#G������(
!��L�z�4�y�)�A��joo����,˚�tmm-�t"����J���"�z:�����8u�=��܄B���-^���'N��eY��ED�fY��#9��L$��7���+�W�`��N�s!�s"���.����G}}�g�7����C&��ٳg��ىl6�ٜ����s����Y���S�r��ѣGq��9��"���iڔ�]�,Kh�v;������	t�+�0>��z�?'"�,�#G���[���X,���V,\����8{�,xn��b1444����X� sJ)��Ӄ�'Or՜��B�^��r�����	:�eY78����[���x�W��Ԅ9s�x~��Uu�4��ׇ��&�o�FQ__���zTWW���t:��G�bdd�`sQi	�Ît۶�y�!&�W�e-pr=t"�)%N�:���~,X� ����7����z?ʲ|"�@]]f͚U���d�m�̙3�����"��`�Yzd��B�B�2�&q�7;w�tuu�N�����y:��xW�B4�)%���'�����<�+cƌ��|�r���p��)� ���R���w�������ۦ~>�p��fdd�N'��`��9��xb<g�̙3��M(����BUU.\˲0<<�s������rt�n�������jTTT�	���8q�R���P����70�j˲D�- v{�&�7R�;�\ﴄ��h*��8s�zzz��ԄY�f){PSS������2�FFF022�T*���躮$��
���H&�H&����@UUUQ}^뺎�'Ob``@u(DT�B���&��e��	:�I���%߳,�Q�vp'"/�r9;v����;w.���W�!����1k֬��ݶm��id2�����:Ø�'�� "�"���(��("�b����R�w��:Ξ=���ޒ�6@D�#
9zqj����Ce�	:�eY��dӊ�.]�q���9sMMM���U�����i���Ķmd�YX�)%Lӄ��t��]R�
�
�|����9��gT˲y
�!fH��6m�ZZZj��)��P"*o������8}�4�̙�&����
w�11'"U�>���9� �+�6vq��ضm۪�����z��i����2$"�+
�B���GCC�����atuuapp��9)��������������_�0$*\A���d2�\��ωH�\.��gϢ������={6���ʒm����CWW���p��
��hY� L�iژ�S^H)opr=��Q��R���===H&��5kjkk�� ��4������{�^z""ծ��!
�&�{�A�B!��!R�b�DyaY�'�s���Q*�B*�'P[[�Y�f]�q9g�&�������3̉�h�7��4�r��ۮB�*�Jt�˲�\ϕ)"*f�eM��G�Q̜9���,�wɶm�?�����r"*z�p�gϞr3Q)�R�C�2�&qy���K&�3-˚	�V��4G ���9!D����?���$�@}}��Q�_4Emm-fΜ�d�]X����A�ܹs��-�JY)僲<��4��m۶b �R���7fTV
��;�m۶VM�V
!�]xS�r៙JSH!Lӄi���r�,�\�i���`0��3�����JD8FMM���Q]]��  �LCCC8w��������i���8N˲<�����'�'�l��_�뮻���O����m۶5��m۾]�+ �U�Tl���\��r"Q�'r剈J����Fee%���;~.��\.����chhCCC�:�+=�^�m���sy= ~&��`׆����1A�����< ��KJ٢:�b�/"�K	!�H$PYY���J$	D"�aM�m�H��H�RA*�B&�jF"*]NWХ����� ��R~���~Au0ņ	�O<�DS0�u)� \�:?a�ND��ƫ������?ŸҞ�f��d�N���d0::�t:�O"*+N�q���rRJ�p0��,�S�	�رc�z)�x���"�	N�]r�E�P�X�H�h�h�p�`p��:Y�y7�[���,Àa���d��:?������$�� ����m��.Ke��oڴI[�f� `��x��	:������4�@ B��������mO< J)/�bY?����s�{�]&���ƍ��/���M�6i�]w�R�/X�:�R�.""""*E���Rʿz���/}�lJ�&A߶m�*M����c)%,�!"""�R��(��i�o�_��EՁB�'�[�n��� � R�glGDDDD��i��g]�� ~��������?�:/�t��}����^u,��	:�*V�� ����Ձx�$����d,� WK��[E""""*ULЋ���������7�Tǒo%��?����G,UK9`�NDDDD��ICd&�u�G���^SH>M�u�ttt<~	&���l^&�DDDDT��>Ӵ,�BGG��$�Jb���=p����������"�2)����d>S
��>A߹sgĲ�����X�t""""*e<j��O���mܸ1�:���u�{{{{Ҷ��`r�Kx�����.�gd5����b���v�R�t�v��'��m���PK�bWK""""*u<V�w^�4����w��_���ڵ��ɹzlGDDDDDEf�mۻ�z��q�w	z{{{L��09'""""�"����4��=���O'T┯��� �ձ�s\A'""""���0��w��T�~J�E,�&��UBDDDDD���"WЋJ���ȿ���7	��;���T�A�Ç���������:���E��۷� �����X�"��NDDDD�g���i��m��s��U�n�~�����!�xLΉ�����ȹ��iwttԪ��{�.r�ܿ��:��ۉ����.���Ei.�����u��}��? p��8���������o߾�s�����݃�����  ߝ]W�д��߱m�Ǭ{VCn    IDAT�/�ٷ��M�\z�}��P���
�7�䜈������'�Nu�(��۷��n�q�;s���o�����\pzqB|hǎT�q9EW����B�R���Ł. �8�M!�))��< ���4-�iZ��r��*)�J k ���� """�rQf%�&����ٶ}PӴC�m�ڶ=u �RV!k�DJ��� ����d2y�m�ݦ�d�bL��'���B����?jkk{������s��J�4ߣi�}Rʏ ���DDDDD4N�m!���! �B���e��{���g'�ǎ;��R��c n�w�y�0�J}��U2YQ���ڵ�J�� �U��R �UӴo�_��P>o����F��	!>`u>��@ ��z����9y��R¶m�ɛ=B��M$[󽒼m۶Ś��������hж�/$<WT	zGG����8.cT�w�`�?��z=م=�!�����b�NDDDD����_ڰa�S^O�����B��� �^�����ھ�:�qE��wtt�P�:����4�3�ׯ?Y�yEGG� �@m��~W܃NDDDD�D��ؔ�d��q�Ƃ���1�_x���NAO&���q�ƌ�@��J��?��c�!!�ݰaC�� �m�6KӴ��]eoUbo�������*H���r����*�رcǯI)�@��8&B���Iu@���{�� �ϫ�c������9 �s�=={��� �?�,�����H�bY�t��?��ٳ^ur 6lx�u ^U�8)�^�I�+���۷�	!����۶}15
���q�� DU��t""""*'NK܋�5CJ���w����@��駟Nd���B�_Q H)��}��;U�Q+蚦�>�G2���bL����m+�6 �*�p��DDDDDDJ���wcr w�y種��P^� B�U� �
���պ Ĕt$���o��6Sq�j����B<	 �b~!4m��v���!�k>{�i�v�����*��ڳgO���k+���C�M�l���ΫB�
���
������s ����S |��rŝ�����`��A?$� �f͚\8�U /*%
�>�8�	: ե��molkkK+�Ñ���� ����c*�zNDDDD~�E���Ј�7���QM��Э2)���J��;w��Ya6���N�1�����E�����|���L&�g��pc���ݚ��&Ԟ\�����Z��M�m۾��WQ���������e͚5����B�룷�DDDDD�B�m��7n4T�օ��o*AB�G��jt)��N�c��/�.M�~��C �FuDDDDD��_�s�=GT1]B��	@�y�R����P�]�^J�E���%��|�i�qјBV�
!N$�ɯlBmذ��?Q5�B�"������j �X���***��h�۸qc��U��N|�_�����ȗ��_���t�q�KCC�w�'T�-����'���bn@a����T���/G�MU&��
���	7��"~�J&��VD>�Y�&u�BJy�������V4��U4�g.����B��&qDDDDDE㛥�z>NJ� Ê�V��*M�W(����lɱm�� �����S����� 6��[J�Lż��}��I5M+���ou�k㋪� """""�	!���:�:)y� �(����=@������џ+��`��;U�@DDDDT�
�-��BL�J2�|j��w��U0��=��b#�O7n�h)��`�?QQ�+DS9)�3�O�Ѕ���*�Z�S0��=
5���O�[0/(�=�DDDDD~Q��ц�����D5)�n�j�V>	�m��*��OѼs�H�C�� """""O���_��+��NŤ���ժ�TӴ�*�-4!DY�9������U�<�+����*&P�`N㗿��i��m�GT�@DDDDDޑR�r��	�t�$ S��5
�T����7��/}�V0o�	!Ϋ��������y�$�\��/4�)��R���� \�	��BϩP����I!�W�4�+�g�Pq�ZD��jt!DH��is*!�Uø��HDDDDTT�^��m�lNnB<��4���ʀ�]JY�n�R�X��T(�:�q\A'""""�?M��&��R&
=�m�F��ԕ����V(�S	!D�����Z"""""�)eRu�"��*�SY��+��rӦM���%�����\'""""��,T�8��.�pO�5M+�]JyN���5k��U0o�I)[U�@DDDDT�
�����	���ի�(x3)�@���5�S�m{��y(�?'QQ*�
zY<�U��IХ�}*�B\�b�BڳgO�U�� """""O-ٽ{wPu^�R.U1��_ż��d�R1��=*�-����(�.�DDDDD� %�t:���IT�R�WѼ'U̫$A�D"'T��������BJ�~�1��B�fd�vI?�_��nU0���Ee%	��w�9
�[��ՑH���]� """"*w:��������Pӭ����-�`^e%� �OŤ��}Bż��u�� 7���x:�'nٱc��AxŶ�M���y�&�{��ѝ;wF��`0�I ̆�����ʃ �q�Axa���Q Q1���t!�+���1M��V�/|���8������p���U�����BMy;���rUu	�eY?Q5��K�H����OhT��h�Q9�kYփ��ȧ��������SU+K���N �M�pdd�c��λݻwG�T���p]Y����XJ��X�A ����������A���Us!��k׮*U��S*���y���M߈�����8}.�3��4?_�	��s��J _Q5�BY�7�8AW�����d�\��y�s�΅ ��:�+aBODDDD�-!ğl߾}��8�˲�� hP5��Ed@q������!�J!~wǎ����v���,�� ��c!"""""�bB�����֎;��+Aحp~�	�������!hR��?�䓳�����ȗ�R�y���
:�E}�n�sO׶m�fI)  �0������ί6A�໊�e����)�;vlB��l8el*GDDDDTR�?ޱcǇT��D{{{LӴ�PX�~��ϯ>AB< �8���R�G�R���q���(��MJ�жm��P�T���b�����2�-t�4�Ǡ>�۰a�9 �� pO*���bO�;::n�|��%�DDDD�w>{�k�־m۶�Ur%�w��b��aձ �~�}��W�������O�R�����c�������<�Re,Y'""""��"xf��4���Z����O�R[<�: �P��\Q$�L�I ]����X,�LGGG��@&�q E���J|��������TD���ttt�>��y(ߺuk��� 6������ƧT ���  �o��y!�ߨ�c�A!�onذa�� :::���<J���������gF��ۀ���B~��f`dF�Im�H�\���B!�/$Q��KNn�/�&��bd��l�%�vX�06���w�I���VU�����xF�����~���9�Q=��������Yֈ��%?_�""b���\Qk-a�X   ��(Ͽ""A�TIlWض��s�=w<�"���?""���,�Ok���6m�����I]D�u�O�H�[�/�Zk}���������O���W������Tr�   ,-/M��k4�8p���$�n�5�\s����/��H�¹��V��κ���t�ED���ʿPJ]�u��VJ��a�<444��v���7k��ZD�N�ϊ��A   ��˞�����M�6ݘ�t��ׯ�V��?�������Rݸq�ǲ��)W����Z��%�MЎaRD�YD>=<<�`�7�����6��J��y�a�֖��
   8�.]�����'�|`�ڵ�$o����T��ok�? "+��w�&��i�s�Tօ4�*���8p௵�ͺ��E�F������7o�?�M.��2��Ed����Ț�JLW���   ,I)%�����Лi����ת��M�R��&W^y��J�sDd���Ar��z	�e�E̗��~�������D$�u�q�RD�+"wi����R��a�h�ka��Z��y���%J�3�֯�׊��i�1E�a�׵8   �qui}1U��R�Ga��0��� 8���1cR)�a8��^��:U)uf�/SJ�NDNϺ��RJݯ�~����\ֵ̗��."r�WnUJ})�:�4:   zE�:Ͼ���:?����)�6m���Ⱥ,�   `qQYh?���y�"9�""�i~H��^    �fV�U���Y�������{E䯲�    � ���_nܸ�Y���t�[n��oE�ڬ���E}�a�   :U�gY�}s뛷�r��g]ı�r�����կ>׶����G록,  �ân��ù��a�ذa�cYr,�����<���!"|�    �
��;��E: ���lڴ�F�Yׁ���  �Nųlg�Z�ŦM���u��]Ddxx��D䢬��3�<   h7��sgﭷ��7Y�\�ED�|����Z_�u!    z����J���ݻww�fX��e�ڵ��V�)�Z/n    ���J���T*ճ.$��
�""���s"r���,�Zz�w    ��=�Fc�T*�f]HT�ED���A�^)ugֵ    �^Qg���ʖR�N�4�<22�Dֵ�ё]D����HD^���nֵ`y��  �NC��(?�Z�ihh����c���ƍ'���E�@ֵ�"^�   ���w��"�����CY�
�_@��r��裏~FDޙu-��4�H�A�R%   @�È�y��Ŀ����oݺu~օ��+zӁާ��'q���W��  �nFC*�j"������("]l�*���8p`���R9#�Zz/X   �VJ)1��
�ZKv̑۝����M���u!I��5�ٸq�-�i�RD.ͺ�^�6�   Т�)�^�m�\�;���߿��"�"�:�Z�U�)�a�q   :B�:Ϻ�;�����7~.�B��u�����?c���暤�:   ��i��i�/��p.�������W)�>��zUֵt�(��Y�  �N�l�\�M)���7~/�Bڡg���7�`����W�����Y��-�   �Fl���_��������O[��
�M^x��W�j���ByY��t:^�   Ѝx��ĽJ�������^
�M=Л��?��d]O�b�   �3E�����n��֯�޽�g�"{:�Ϸ����Ȩ��S��	   ݆������|nxx������^x���W�r�a��Z�]DNʺ����   ݆&Tj��D���r��r�|1��8p���D���9"�9!�r'j@g�   򎀞�9���^D�߸q��ԱiX=�/��x��_�r��oj���5yj:��"R̶�l�>   ݄�ٜ��'O�~���n��7�|�O�/=!�\s�� քax�R�Ok�JE���`�)�����	�   Ȼ�����K�H��Zk�Ԥֺl�a�4�{��Y���H�UW]u���r��s   �,�k�:+�Z�;��p8��O#^�V)   @Kb<�ޙF�=t$"û��   HY!�#�a�A  @�"�#V��;�ax�rBw����4)
m�   �����b��ض-�e��8�<Vز���X���!1W]u�aY��8�}_|ߗz�.�FC|�?r��5k�n�   �*9t�г>��۶�q�#�ݶmQJ=144tb���AGb*���Fcu�ѐF�qܣԂ  �   W�:mHk-�z]�����)���vՆ�G@Gb��j�R�,�z���q�+   �i4˾Vk-Z�S,=�M���MQ����   ���%��a�wS*=����X�uE��	�   ț�Sؗ�4�+S*=���$}�0�e�:�qש   ��a��S�4��w�y0Œ�c�HL�T
,˚�2&�"    -QgxZ�5�{�n:NH��,�(�3�   y�yd�f�g_�x�H�al  ��u�9�!it$ʶ�/E�>�    ��;�_�R)�Qt$j˖-�6Ms��p��A�%   ���~��R�ts�%�Б4m��Q0�   Y��=�,�1Y�	F�rБ8˲n�r=   Y�q���S*=�����qm��Y�  ���8b��JA#�#q�m�SJ-����}   �$�ay����AG@G�l��eY�(c��  ��D}�m{�T*=�R9�at�²�_F���  ��D]ri��=)��G@G*LӼ!���C  @V�>��q}J���Б
˲.�r����5�T   ���?w'ҳ.�\t�b�֭-�Z�+�֚i�   h���7FFF"+,��,��(��  �n16��7�R :�cƷ�\�:t   �[�gP˲nH�������}!���F���  �6q�Y������Ԝw�y7��,�z�u�:   ��bt��m۶ݔR9 �Ҏ�<e@�VK�   �(Q�=m۾OD8z�!�#U�e}+��l  �v����7R*:Rf����\�:t   �C��ϕR�I�@D�H����M�mGZ��n�   H[�gN۶k�R閔�D���60M��(��  �����-˺3�R�#�H�m��\�Fq   H��:�3�aW�Tp�SJ}R)����0d�8   ���}�z���+�dpp�_S,	:ڠT*=hY�L�1Ls  @Zb�?�<��sM��:�¶�F���  ��T��H�[�u0�R�������r}�^�5   $.��j��^�R9�Q�h�0���)q�   I��9�i�ᩧ�zYJ� G!��-J�R�q�����:�   8��K)ǹg�ڵt��t��Rj����z��5  �c�s��eY_K��Y�h���7ǭ   +�F#��j��bI�Q�h�͛7�o��d�1Q��   �u	�mۇ���N��Y�h+۶o�r=��  �����u��R)���h+˲"Mb�;   ��_�0�1�r�E��V۶m��mۑ޺d�;   Zc��ڶm۾�R9���h;�q~�z:   Zc��S*XmgY���r�����~Z�   ��5	� ��ԧR*Xm����4�H��t�  W�gI۶}�0.I�`It�]�T
\׽#ʘJ��V9   �r1���V*���܁Б	�0>�� ��  ���Lo7��)��x�_�/�iF:�3�  U���e'�xb�f�:2�v�چ�wE�:t   D���8��֭c�&2A@Gfl���(׳�;   ��3�ݲ�ϤTp\tdFk�I˲"Msg�8   ,W�gG�4���~֟#3td�T*Ulێ4ͽZ���:��   �%�֑�H��{����*�:2�8οF�>Ci4i�  �.Q��%#M��q�9�r�e!�#Sk֬��eY����;   �'���~��K�`Y��Ժu�|�qn�2�V�1�   K�ZGn긮{�T*E�QH�3��Q�Ð#�   ��8�ٶ��)�,�۾}��lێ����  ��D}V�m��u���S*X6:�@;�sc��Z-�   �~AH�^�4�u�o�k(�9:r�0�����4�i�   X(j�\)%�B��T	�p����8SQ�T*���  @�����8��������"!�#7l۾,����s&:   ���둗Aڶ}IJ� �Бn�f��?t�  �uz�i��0��)�DF@Gnlذ�1۶�2�R�H�i�  ���s۶V*��L�$ 2:rŶ��u��   �����R9@,t��]w��)˲"-,���K�   t��τ�m���ϦT��{���u����}_|�O�"   �]�^��<h����w�f�$r����q�Q�D��  л�l����JZB@G�lٲ�f�u�2�Z��Y  @
�0�D��>2::���Jb#�#�l��T�����	  ��gs8�q�)�r��БKg�q��,ˊ��hnn.�3   :[���g�q���R9@K�%��H    IDATȥ�k�6��V�1AH�^O�$   �L�Z� "�q]���k�F:5h:r�P(�>��  `)q6�+
�B)@"�ȭ���;\�}8ʘz�.�o�  t;��#Ϟ,
���?I�$�et�Z�P���c�  t�8�s˲>�B)@b�ȵ;��ǉ�={�V��	   �#��ݶ���~��O�T�:rm��ݡ�_�2�#�   �[���
�v���T�:r�X,~�4�H���  Н�֑�4������T�:roxx���y7E�!]t  �.T��#/gt��y��xJ%�!��#x��!�\  @�\�t�RJ��HJ� �"��#�w�y?�<�(c|���5  �.�h4"?߹���m۾�RI@����m_uL�wX  �_q����)��B��:�ڳg�T�V�2h͚5b�fZ5  �� �C�E���]�V���::�.
��:hvv6�Z   �F1���9:eŊ�8�eL�Zߏ4   9���T*�Hcl��O9唏�T�
::����ˮ��:��  :W�����:�h��g�ʕ�7#�T�j���L   d/C�V��Ƙ����H�$ 5tt�s�=��B�pS�1Zk��   (�~B��������)������T(ޫ��4�R��E  � AD^{���B��JRE@GG��P(�e]t  ���٭P(�222rw
� �#��c����/N=Ô*  @R�v�]����JRG@G�:���z���(c�  t���9�:���ݵu���T�:::�m���0�}����E  ȱ0�=�PJ%mA@GG۶m�7
���Q��E  ȷ8��B�p����u)���u��g\�E  ȧ�͔b���S(h+::ޖ-[x��P�1t�  �\.�Y{~��͛�M�$�m��
���n�1�r�s�  r$�XM�uY{��@@GWغu��
��#Q��E  ȏ�k�غu�)��]����CQ�E�����  �q��O���{)��]c���_v�Ѩ�fff�(   ����c\�}x�֭_K� tt�q>��^�դ�h�T   ����X瞳�݆���r�|9��""���)T  ���,�8ν۶m�J
� �!���8���]�z�.�Z-��   ��F��9����M�$ 3tt�m۶�P(~u���l�]C  К8�����m۶ݐ|5@���J}}}��iFJ۾��E  h�j�y/ ������;���L�ѕ�?��;]��n�q333t�  �@kk�y�P�i��ͷ�P�9:������i�a�1aF>   �U*	� ��4�i��H�$ stt����G<ϻ2�8gp  `��0��s��۷o�7���\ ����X�❖eEZ�w�   ��\.G^VhYV`����Jr����6444�y޿DW.�#oX  ��k4��
�-�J�)��]O)�a�q"����  �c�3SѶ�O<�C)��
]�T*��~4�F�!�j5��   zR�V�z�y��8�n�:?���\Q)�^�gϞGk��IQ��!k֬�TZe  �C�E޹�u�Gw�����Jr�:z�mۿ5h��a   G+�ˑùRJ\�}OJ%�C@G�ؾ}�~��n�:�R���3�
   � be�R��Jr����bYֈi�a�1Zk6�  h���l�c��=�+�T�Kt��R�t_�P�8�z�Άq   1�}�*
{�l���Jr����s�I'��u�XǮ��"  ��i�ezz:�8۶��<����P�kt��u�����}(Άqsss)U  �}���"o'"R(>�v��F
%��1k�Y{�R�����֬Y#�i�Q  @��}_>y\�P��Ν;�H�$ �蠣gy�w�i��ߡ�3M  ����d�4Mm���:=kdd�b������0  ��*�������<ϻ|tt�G)�t:z�)����q�J�q333��Nk  �	a��l��xŶ�j__��J:=�Ϊx���8�q6:  ���md
�?fG^�46�$��q����8N%  t�z�.��
���ܹ�)�t:耈��9l�  ���LMMEg�.��P�q耈l߾��B����� ���
  �����ƚ��yާGFF�N�$��Ё�Y��۶'��+�˱v)  ��FC*�����8�����BI@G"�O+�JA�X�g������  �EZ�XSەR�yި��<��̳m۶����Q�A �r9��   �mvvV� �<���m�vm
%��,P�Tγ,�uS� @����27�d4˲��emI�$��Ё���̸���8c9  �
�u�m�R�����R��N����,a�޽�V*�WDW,e`` ��   rcff&V��P(�`�Ν��BI@ǣ�,A)��4�F�qsssR�E�!  �1j�Zܩ�b��!����@@�066v�X,~8�����X�  �]���������ᑑ��	�t��Ǳw���*��oD�8��Q  @f����Z�FW(nݹs��J�t�8<�{�eY��g���)  @^U��X��4�F�XJ�$��Ё�9\(�(����Yi4"/c  ȝ bOm�<��GFF�H�$��0�X����۶-�����J�,  ����x�<��;v�&����CX&۶�lYV�9]�FCfg9�  t���-˪�ȹ�Wt':�L�Ri�X,�#�X�^  ��^�K�\�<N)%��{ǎ)�t%:A�T�R�X�z���  :M�255k��y_ۗpI@W#��y晛]׍�Np+g�  daff&V��q�陙��)�t5:�ڵk���4��;,�j5�^  ann.֑j�ah˲�{����Q6@Dt �R��b��Oq����J��Xu  ��ie�[��>366vc�%=�cր�ݻ��J�̨�Ð5k�p�  ȝ0e||\� �<�u�v��uZ�U��:���mێ��P&''�7�  @�����
�e5����S(	�t�ccc�۶��8c�Y  ����ΕRR(޿e˖�S(�t�Eccc������3�\.s>:  ȅF�!333��
��o߾�3	��:� �479�s8�����X��   �A���m�����H5 t �R)(
����P֣ �,i�ejj*V��0��uݷp��:��R��㾾�?��3���2==�BU   �6;;+�F�|],?�}���.	�Y�$l߾}ߜ��{s��+V���.	  `Q�ZM&''c��<�;v�xk�%=�:�0˲��8�q���̈��I�  �,����m�۶=�pI@�#�	{z=��,ˊ����299)ay);  ��5����4���K�R=ᲀ�G@RP*�����w����]TY~  ��ʦpJ)�<R��)��<:���[������gl�^�})  �����J����y�W�o����K�46�ҥ.���{����q�i  HR�R�}r���ڵ�ԄK0t ]�q�Wٶ=g���t�w�  �k4�g虦Y[�z�o%\��@�J�Ҹ�yÈ5]err��� @K� ����X{������6<�Bi �!�mP*�n,�gls#vv  q4wl�����GGG��pY �t��.������[�uGV�Z%qv�  �kbb"��9�u�۵k���K�:�@�ܹs��8�����   �V���m�W��%\�c ���\�r�eY�8�+�����k  ]�\.K�R�5ֲ�����+J�R����F@����{�X,��4�X��ggg�V�%]  �"�ZMfggc�5#,�C###O$\�� �(�J7:���'''��h$Y  ��z]&''c�UJI�P��R�tc�eX6�2t�%�|�\.��8c�R�z�j�,+�  @��}_���[ٱ�;v�xg�eX&:��={��R��^g�i��z�j1&�  ���0���q	�x��]�=�k׮�&\�x�2677�Z�q�36�t   �ùmۏ��ͽ!� DDȁ+���ĉ���|��⌷m[9# ���Y�i�����V*��L�, �Ar����6#��ލFC���b�7  �Ik-SSS�����7΁| �9Q*�~\(�aF����q*  �3���J�Z�5�0���?�}��[.@Lt G����y��q��������L�U �<���������]�ݽm۶�,	@�X��о}�>;77����������/ɒ  @����f������ t ����{C�RyS��R,�,	  �@�Z������=ϻ~ǎoK�$ 	!������sW�V{I��X�B</���   �j��LNN��v�zy�%HkЁ�����t���i��jI�  2�j8w��N8�	� atЁ�ۿ�������F��J)Y�r����ti  �M���LNN�>Rղ�Y�qN;�pi Dȹ���C}}}��,+V+\k-�����G  ٪�j211;���Y+
��p�� [�n���o2Ï{���Ii4I�  RV��[��0��7l߾����:�!FGGz��v�Tg��Z���� �!�FK�ڕR��C۷o�9�� ���t����o���a��<�N:  ��h4Z��n��<�;v\�pi RD@:���襮��vܐ�����	B:  9��pJ))
�r¥H�@;v��l__ߟ(�b�o�t�� �/��y�Z�&""�b�����>�`Y ڄcրv饗��r����|��8	V  �H�s^,�vtt�O.@�Ё�o߾�W*��'� йZ�""}}}��@�eh3��nll�#��4��s� �N�^oiC8����!���:�%�����J���V�r�J)
I�  ��Z����tK�X,����ػ��
@V�@ٷo������K+��b��TI  `	�jU���Z���y��رc,�� d��t�K.����ryK+� � ��r�,���-ݣX,~ill��PI r�5�@�����wY+����i��  ,�R���s��΁�C@������Ba_+�H�}  p���Y���n��b�;v�ؚPI r�)�@ۻw�W*�w�r�ue�ʕ��J�,  z����T*���Q,�����#�� �t���ر���ϵr�Z���  �2��LNN��=����ntЁp���c�V�`+��e����� �\a���4�����9��-�� �O�@عs��z��Z����211!a&U  ]-Co9��ŏ΁�@@z�����y��׭�%�}_&''Y� �q(��V�I-�g``�/���� �� �S܁��/~�wggg���:r�6C֬Y#�eI��K `J�#K¦���\.G��a�X,������.�� ��A�^z�;���>�a���f�q���Zk�� 0��p�4>>.�ju��0C
�w����{���7:У.����J�� ��\?88(��=��t� x�b��СCR�׏{�0B�uK;v��J���?:�������Z�v]���[�r�����^��� �S)�����0�СC�����������[*���F� ���K/��׫��|�v{\D���eŊ˺! Ћ�X��AȓO>���0˲*��vll��4j�� 䢋.z�R�'�z}p��=ϓ�����-�)� �^q�)�Ki4r�С�~Vڶ=����[�ly8�t: ����k���Z�T�ue��ձ�T#� �]�p�T�VebbB���8�#��y��ɄKЁ� �����F�q��h�}�s���y�t @�j%�7��e�V������R��1 "B@����a���>8� �m����8���6l���$j�=� u��W��Z_�D��_�4����  �dɄs��:ܵaÆ/&R����� ]��o�W���uY�1�KjNL��  @&�Rb�f�?˪ڔ[���p`)V� ȯk��y�B�f=(+U��{���t @�Ib���ȴv�:��2-�]	��K�ApL�ڑ���.�|/�0� :F��V��}rE�t��-��� ���M��q��"X��Rt @�%�<��p�\�*�.�� �%%��/��O��X�>It%  HRR�\�ȏ���w��I��. ��t ��� s�#o�K���|�i�M  kI�7�Ő����@U�%�� Dv8 �JY�-�+��!  Z��̮Ym���i�s ��T ��ړ���ca��q  +I�&"�hX�+�ɸ.$P�^D@[U,��?Unִ|/B: �ݒ����`P�	N��f38 �@KBQ���2�y������N8�a�֚u� ��$�Qr����J�~ z@"�WɌ��[̇�����՜n��h�ַ ��$��%��O�'���� �)� �D����{P�(6 @�����.���$�'_ ��[4N���Չ܏�� �V%��D��O��r��T��
 a�� H\(Jn�O�_}��qTk�ɕR��bm:  �$��7Đ��'�}��D� ���p@&���-��2��-߯����fm: �L3�է�+��_ ��M� �S��jJ;rE��v�e�; �x���&��p�\�8�p ut��.C��?O3��:�11��i�� XL�o���f��rgxB"���!�h�{�U2�(�:�aY��-ߏ��  MI�5yjJ����8]s m�w muH䫍�O�dvyy����@oJ�X��v�9�v����1�`p�<���z�Qq$h��͝��@�H�k�C��,�d�v !�����
9��d���<ר$r��A �W�M�$gN=�=����h'�{@TLq��Ym����� �x��� ȇ�O�Pr{�F4N#��O� 2��'�/�	b$�Iz�#  ;���$_���^=(?��+���	����
 7��+}�)v�_͝ޓ�
	 h���"�R�g�2+l ?� rE��gRVE�j3����; t�4��u1eF�h����@.�Œ�6ΐ�������3� �/�#4���+�IUXk ���@nUĒ��ʯ���*�	1%L�͠�N� �?i�x�Ő���g��� �� rM��O���`�/�7%'s���0�Z� ��4�NyB����d��t :��0���?M�4'�5��b���J)�ZK&sO ���}1����=8A��� :@��"��`P~����_��rb�f�; �_Z�a>�;��2�� :@ǙѶ\�*/1&����b'�6]�i� �iu������w��5Й� :������P�_^g�J^�p7�9흠 �J��ˇ�~�^p�������]� :ZYl��?U^h����cR�Fb�f}: $#����S'~��?W�	W%~o h7:���`8 �Ջ�
�Iy�9!������t�: D��:s-"�W���D�j3��@� �F]L9�$��+�l�1T�D��Fr �|iv�ǵ+��'Oh/�{@�� ���(�7N����|2�#ٚ�� �: <[��<CnN�ۂ5rt�.D@ЕBQrgx�<����r�1���AP�g��ED��}�$�e8 ]�����hG��O��ey����T����f�����ڑ��I�P؟�� O� z�#a�|-|���8,��:$V�g��p4�ޓv0ohCn���	Lg�3� zF Jn��=�U�j�	y�1��#A@/H�,��������� z@ϙӖ��?O�6V�k��w{!��Ni�á+Ó屰�ڟ yF@г����ty�1%g��%�ۻ��A�3�t���y]rsx����tv =�Ⱥ  Ȗ�{�Ur{�:� �<C���; �RJ��4S�a���j�y0H8�������.w�v��A��� �*��ߚ��,b8 x
 �0�T֨țvs^� `qt XD��]A]�7x`�nYt� �#��1��i�o޿� KX��v����1�(� ������45�y���vu˛� �� �vM}a�;��3���" �G@���iC�ƕ    IDAT��DW@��.�� $�� -h��."myf�w �Ѯ7E� �$: ���P��ܭ�A}����1����-!�@� ���Cjs3�v=(ϟ��F@oi���xc ���Ws ű������5w}og`VJ�i�m��
 �����0� ��w��?[`Qt K�3��i�+�M�ܘu-�j~Po��l�{OX�����v���M��x���Og]��"�8��֟X�
�����4���{
:a�|�.y�����[�D�,�qғ�EG�i~X'����^����E0��u�K�,��ғ�ugjaW��do~0�"�g�b#����`����rӥ���)�@{5Cx��P�w�9"q�s ��DBHO����,�W�;����<�7Ƙƞ*�9�X� "k�t%�?����a��bk`ē�Pޜ���o�#���� ��֟X.x�Bzz�?Hg��j�,6�:�³ʳ��Y8��`�*�9����FHo�<u��w�Y�<c�2�,�*_(�qz�@�� ZBHo��u֭�.y^ް�[��9�D������fP��x�g�[�CX���.y��ny֯=�p 1�����ҳ5��</v�	��47w��Oyڧ���$�� 1���i��<���}���t����N������� �H@���0�8�<>�/�����C>���!�H@������>O�����tIk~--���uF(�-�9�������O������>�/RySȗ��|�t���s�p Ut �!��['ǴX�3��[l���@�w��A8��������a~@���˱Ԕ兛��;����Ra����	��p�-� RGH�<�֛qC{���^3��h���bo�t��3V��p�m� ڂ�޹��N�C�������:�b�������Ŗ�t��O#�h+:��!�w�n� .��3}�؎��^lZz7�.�=�M�'=�p��� ڊ��=[CۍAd��Ŧ�/��.�n�=:ͱ����/�������b�7t��A"�Ȅ�u z�E�O,����7T+��k�o̺�na(��@v<�u֏������Q��?�p�r�b���R�r��k���F8�:� 2A'��-�*vs�=	�C�bk���|9�-6n��~��4�n����8
�@�� 2CH�7�"� ��#�k�g�d�� S�����Hr��`��!��{�@.�d��'����U��Yׂ����w��%A	I9�C|��.W�Km$��:�\�3�����'���p� E�±,�:��o8����/�Ⱥ aw 9�JXͺ��b�j�glt�{�|O�FTT�� �� ��5z�B�P�}�{� ݆� �J��/�<�5�����q  z �3��q_�׋}�x����� �^G@ @��5e��C�bgLE  :  �%p�_߼�X]��Y����?�n  �G@  ��ظ�6�0�j�&� �.:  9G0 �7Y      �     �    � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     ���.  ��W2 umf] ��CR̺ �: �ȸ.ȸ.d]   zS�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     � rCk���:�B  ]2�� @�� rCi]m��R</ �a�g~m(5�]% p4:��0���/	�� ��	��Z��t�� �Q� �#��"� ��������W@{��y���~��Jt @hY��>�3, �B@�SA�����  H�
�7�uݶ�ɲ ��� 7���j"�@���Z��  ��U?�k-�Ⱥu�f3, �B@�+Z��_�bV�, ЅN1�ٴ]i}0�R �Y� �E�o5���o  �z�����Է�q) �@����V���6�Ǻ �e[��G-�҆A@�+t ��Ʒ�����͏_jr<-  /�fD=���ox�[�̮ x6:��1�/4�kִ� h�-/����֟Ϭ X@�Ap���"O��~�5�qE �Nw�9++�#�wbgY ,�� w�p*�}͏_c���� �I�ȫ��y�P_z�9�<�YA �:�\2��	EDVu�u��� �x~͜�5�l�C�>�e= �:�\z�9�ܥE����l��T�eI �TP���9��'������ۗ �!��-���PDfED<ț�'2� �i�d?)�3o��)��H�� �����o=,Z�U��X3�rk*˒  �%֌��:j���>�-oy �� ��� r��8� "�m~�f�	9ѨfX �<Ǩ�ۜ���`��>�z `9� rmݺu����"rHD�RZF�GdP�3� �W+TCF܇�zj�Q��@뱵k�6�5 �F@�{�54��6�w��g�T #�G�g ����0|�RxD�Ϭ;���x����eY ,@Gx�[�z�h�.��D_���}P��̱9 ��ڨ��YVZD~�����ϰ, X6��κ X��\w�G�ȑ5�5m�u��䞠?˲  ;Ü���c��Oj���[��o��
 �!��8߻����ZJD���~�X%��#�VV h7S���9$�iMȼ� �����_����U ��t�o_{�fC�/�ȑ��Th����}A_�� ��TsN��<1J��HYi���ׯ�RVu@\t �W_�1�/�R�1��E9�8A~zY� H��FU^c�����ߺ�T�מs�]Y� �"��h7�t���|L����X������+�ޠ_�	 �RZ�0g�׭)9Ř[�ہ��W���k����� �)� ��w���7�0>�D�^�{u1�>�O��PP�imgQ"  ��!��y�Q�ӭ�8.v�����9�����@�� ������o�a�QQꬥ.�jS&�-��#�{w�i]p���̮�e�nfVb�ه�EE���D�DHt$t�IJ�P�AD�lV��a��b��k�����<���;�����N�{��f������>:/�#ci�\�dZ��9�Ǯ���{<>v/���Y���m�<_���P�-pJ��)��7���y�����1�g��{ ��y�ʘ�Ͽ���o=�� l7���~��z��]��1���1ƛ��� ؔ�4�2������߷o���T!Ё��~�g����-O�E�<�p��g���4����p����;:�y"���Ӂ�<oi��C��GO�li��l�M�:��v�#���V�����//>w;nZ����{y��mu����5+�:o;nZ����}������=�o~�wz���ᤅͻv=8_rɷO�3��y>2��1��y����y��k���d�p�t ���7�c��O�C������ꚿ�x����|���������꒿�|��1�۶�����W����.9t��4��{��M�����ƭ.�}Ϟ�Mc|p�ٌ��=x���L �|�   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t  �Tv  IDAT �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �   +'�  z����e����c��s�����}s�}��~�ɛ�G7�Y>:�̍�rdZ{��ii�F3����W�i<m�}�<��{��,?���fn<�yi��8�v�F3��s���K�Yd����}�>��l8�c��M�x�g�G?�6�v�F3w������Z8�����޽�Ȏ���&N<��ȑ��KK��h��k���ع���y>�c{�F3k�ˏo�F �: Op�ַ�q�ׯ�暥���{���{���;~�ջ��+^��'�yt���O_p��g��E'���^����lf�O��c��Ⱦ����K��-��g\�}c��6����������<x�uw�����C��cܿ������c���W=��	��S�?q  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      VN� ���������_��/��q;�0M�c��������|�f}a��������}�&�4Mӹ�>r\/٤i��<Ƹc��y�׏�9 ���y�O�   ��O�   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �   �oO�=�     IEND�B`�PK
     t$v[�����  �  /   images/50196d33-890c-4789-8115-a73c306e50dc.png�PNG

   IHDR   d   �   1�S   	pHYs  H_  H_#�
{   tEXtSoftware www.inkscape.org��<  6IDATx��]	tTU��߫Je��!$�!�g��6=Ҩ(.���ʸ�8�L�����l=����Q���s��TPQ��i!�;�RI*��7�w��QVBR[.�snR�������/w{�Ig!V�X!���wEQ��ɓ'���	Y�|y���{G�_}��$+�#�#!2\��p��4�S?N�8p�6��sj�t�S�}��r:�)���#!�/���6��ʢ��zr�\TZZ
�3�����Fs�)�Lb�0]m�p���jNk�>;N�8A---���S0���|�6m�4z��7�|�|>y�^
�����!��n�t�r?炄��|�k$����B��_TU]��|����I������/Snn.�z��S�BV�^M���'��!�BX+.b!=�?���
5M�&H�i��Ʉ�p��Z1���_��]>�[.�_��ЪW^y�***zĜe�����Ӟ={Dś��A�(n����n���V�����aw�\$��M|�B&bV ��˰��o���-��Ç��W_�;３2�����R|��%����A���E��@xH �
� 9�����"���l�nf�y�_h��d����L!#����k�q��,�k����	5FK�u�h�~qq1���B `����yp�0�@GĘ�CC@^��\�����s=��L���//���8�;�t#��D�YC3X�N�l~ɇ�����yB���d���'O���ǉ(� �ȷ���(H9p� ������q=�%k� N��5Oq�ebC��2k�,J'�J*��@,�J�ϯs�����(�'�B��۷/4HwӦM��{=Fk.++�_p�"��������} h-�ǚ6��h.�L��H&HI!(8BZ�<BN5��-p�0��� ����Bv��I{��%�K��Q�����444M>|�gw����{�}!&�J��Ϲ�S�~[Q�t��B�X�Ͷ�H�誉`�����O�>�a���Ӊ�o�����I:":t:G�-|��ݻ;5_&p-�())!��al�V��k�N���������|�r�Õ��������Q[[+�8��BP��������9��t��$��ѣ�̍5
¥cǎu��({�����;N�0��k�}J	Aag!�p6ˬdt�`�]�0=<�����Dy�^�)n��ܐP�V���7�	���K��P�s�k:$L������[Lu�dR�q�.�su}뭷RڳO)!f%��y�%9$������oX����}t~�TS�Z�:ı s����c���Hێ���R�)��+D`�u� u�bs���v%׷av*�2B`S���t��g$�w���)����EQ�|�]�o��&��שūS����U�0?�*ˈ
rw��̢���bX�~ɑ#GD�мD�:�������a�宻�T %�`��O7���E��	�9QY�E�}~ꗿ��P	-�p�y܇p���$��O��6���^���u��' H4��j	ꄺqg6[�/�����7�x�n��6J)!�6�Qͅ{
�3��5Q8�S�W�@{#UV�Q}#n�n�\�+9��0\d�7�)T��Ow#��#B���@���Cc�Kʇ����}���|�sڇ@&H���p��>��{*��(-4y��- tA	���,��n�D�񚮑檢��

�7��{���z�����s�Q�)�#� y"��5���aʸ1>��݂����N� iB�a&�Ӡ��k���ؚF�s]!*+R�Y���ߙSN*GQP$��8�F������H>
E˅ԕ��3 /ԕM�t���l�>46�AR��E �*//W�I�;�~���
T�n��Ǡ������k�{���J�F�[uD��t򴅩͗ł�3;{�;Yᙦ������o%�'-Y-I�S;� 7rEǂ�TL(��'C�☪�TJ�d�~�(!Uk�l�@s3��9�Q�S��Dda*X'�X"R*l>�:s<�;�7����Z�H�L��Rk׮��c�>'ם1�� ��H�,�8�H���2�q��z����6K�"��;�ueq�J
T������ɕWN @�З0C��:�x@٠%,<��W_-7n-Z�(����	�v@�/�䒉�u
�
퀐�7 �g���.���m����)l�t��ag_����S�i_v�7�{�Y�LUUU"��X[*1�B&x��_<��Zs&$L̉1L2�abRA�|Ё1b��8�PG�O�Qaqmo�kj�n��bk������: L�uY��3��J+�d@���{��%F}�~I*��ct�-�,��+���w���mq	;���~C� �cr	-C��ׯ?%@v�E%���c�����
����{�]t�[ʡ� *.u�5�7�6l��̥$e�2`B��L��6%j�"�r�yMdZ��E	]���Fh�B۷o�0����D揠&��y��1�뢜�����:x�`��5��T��?�,8o��e��q%D����&#bId��L@��#0/h��\��x!r�0���-�9�p4�2�5���z���ư4p2�s�fA�����&e<ZF��J�?HA$MA��Sb�C� ��C�R���ŸFx�A�	Ȃ	�`>�<���{�uz�;���C̥;���)�~����ǋ��5W<Z��j.t i[�lI�߈�!�!�P��=�����k�s�4B�-[7����;����{�	����o�H-Z<�4���������B�t�`"���퉕��8���u�]=%��&�:�3��?����3�7�J������A�LU�x&�2��
!,BbhLʁ^=��.��ݘ��Hq/L;3�eA?J��4��Y���巔˥��~ʔ)�x&����l�;�9bo�h*Ժ
ӡ�h�y�jj&��-#c0�ep�L�t��C����돂�v 4���s�wqk�nS�:Z&�)mMVY��C�?��3�Db�ΡSd ���8ab�aN7[s�)BdF# �9=����N?�_YC�O�'
B��'�������ZN�8M1��	��B`~�]����rz��~;���n�d�>��"�ŀ��ގs�ߓA��.��q�A��I�my�Ld/V]X	�m3�)A��]��l͎#d��VB�Q�#�v���$NKc2J~YŹ�죘c�m���Ed/`u�`���o/prsZ�)��?p�����Gǈ��`a��sـ�������Y���ԁ�)Ia�$��p��(F�-� B��"۶���RD�QB0�`?�ɩ�re����C;��.:�����[N�)"s2��!�&M�vwP$>�M��D�Ctp����d�4��8<I��9i��E�&�����	Q��^����#��f<t�Pߖ-[n��oc��,�!g,;ǜѣG/޼ys��!����.� W̰�w2��*��UU�eee��2�s��x<~M�6�[�N+..�t��)o+�J2މVO<������B��Xw���d����ۇ��3�1j�0Smmm������T/r8[�imn�b���L"H��ọ�`B�Ҍ�c�2 c��Csn&$�!�l��l7����q�\5[��>Ȃ�g8��E�S�E�^��(�cV��,��> �n�+�q6�\�r�-	�pxf��z�[���s���y{���p�	!���pbڭ:~���>�o��5�e.gR�.--]�9�d�	_9c�z�����1̅z��2������I���N�<)�,�� �T����r��d2���Xr�h��l�j���&d��:���9s��6W~֌�q�ކ��+����Pw� �z|���A���~ayy�=�����^���%�^��Gl�b!w*�u҄�E`(OG`<�-e"kJ^�6���Tq]�l�bq�e�xx@JF�%X;�v���>Α�Ӱ����#�1+DS�e"6�<G%H	!x�/444<Å������TR&����x�,����L�e��@��͡�x6!
ȶ�^:z<���<|FV�OR�mc��
��!�)�Ȁ�¶n=�l[�s���)�>�� f���il�q<�CF)%jk>M����tS[[����fR̈��Ҋ:1�憠d��X�|��?��1�۽�+3�+�9�����fpZ�tnTk@B�t<d9-s��' ,G��*�i��e-r�JUH;��ĉ�8�z��4���۸q#�3&e�����(M0Ii=q�<�/\�5�r���hG�?��m.�a�Mrk�WБu���J���	���7nXz������8��h�<\RVJd��6����$/9�������+��<3���"Ӗ��� ]���/B}Hw�4@�P��% YgqjS��VHk��u%�4��(�e���U<�R��z!},��T�6�blc�I��n�N��և*�\��f�$D�K��9�ݵ�.Z��3L�Y[��n�$^ܒ���]����$ܟ˨So
��8�w��$�N��=���x����v��Q07j��s���6Y���â,f�,�|�*�2B*l�:�����NJT[�	�O=&ܺ��JL��K���EM"N۹k-O�\�>�B�� �t#�,���n^��[�Bx	G0�r�6����b^OtZ���yM���y�$t.�/K�f:teI��uI72�!��"����n�9L�z.\�����ƕNk��-=�X<$��|%�n������B_Z<��2����ES�#D'�9��QB!U����wk	d�@�7cd {��Ӕ��qf�ʜ)��$C�����MO����Ä�䫄!�0��;�B�=kP{����+������+�)�L�C������&�'D���PH���R��N=����)b�{Z?�A�+�C�'�o�K�<$9\J�s��x��QB��s�P�|m_8���ZN瑍�G=�\��q� 4{�⛘�0M���o�)j4KE�_��{�>�q�-��˚��+��@���˛�x����?�*�I���C
��%��x�~w��Vs���+�+P�թ�r�JP��Y>$W�ݭjaQ��3��	ӝ>���RtEՂ9y��3_	5�t�<��wؒ�JVӗ��.��(!���V�	��>���ϋ׾��߯�|�y�;��Mu������!��
�]v~�ҟ���4�aԘ���ի��ʇ�EU��u��~z��'�0f�^�<�����C;ʎk�>\ê�V�=����*ǰ!~��nU �SC��N��3��Eɧ�&Ћ����$2�C��
�]��-�3}�>���UolSݰ1L��9��]�+!�Z��Z�~�|�Ps�x��<���:Ԥ��NGsS?�m�Y�z?)��������{����`4��]�����c.<�W�w(=�����e�Q�L`M�W.������r�vD�cq���a���12Uu�A�Ug������E�tjϊ����Y��_.2�j*�� ؈�&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!�AvB�F�7^�c}em���cx��f�-������bRU�9d�2/z�G��(d���Q������lRH9���E2���i	i�T	L�_�=e���ƽ4����;JS�v�\�H��7wDs�9�@_V6o�[��5��ѼuPq~ۃ[G����|���yb�纮O����F�νt��=+W�++#!-!�K4�!eǶ:�G�Юk��z�ӷO����˟�y߆����Z<����^�վ�R����zޮ�:��}'���y�-j�5k��Ңy��K�������O���~�j���6��R��P;ɩ����ͭ��IΓ��@oR�P �@����'������.&�&r45�F�fo���].��m���X �]����ǜ���{<�:��C�z����d섄9�9�5��o���9揓�t���)S�й��Ǵt���	    IEND�B`�PK
     t$v[��� � /   images/f158dbb6-f78a-4fb5-8a82-0ff8626242d4.png�PNG

   IHDR  �  W   ��5�   	pHYs  �  ����e  
�iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 9.1-c002 79.b7c64ccf9, 2024/07/16-12:39:04        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmlns:stRef="http://ns.adobe.com/xap/1.0/sType/ResourceRef#" xmlns:tiff="http://ns.adobe.com/tiff/1.0/" xmlns:exif="http://ns.adobe.com/exif/1.0/" xmp:CreatorTool="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" xmp:CreateDate="2024-09-25T10:15:37-04:00" xmp:ModifyDate="2024-09-25T10:18:25-04:00" xmp:MetadataDate="2024-09-25T10:18:25-04:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e0fa026c-2b50-4255-8fae-7a1c4254e60a" xmpMM:DocumentID="adobe:docid:photoshop:cdda18bb-8c9a-7446-b932-ddbadfa4c834" xmpMM:OriginalDocumentID="xmp.did:8deed1a6-5431-4e06-9973-719a94ef57a4" tiff:Orientation="1" tiff:XResolution="1920000/10000" tiff:YResolution="1920000/10000" tiff:ResolutionUnit="2" exif:ColorSpace="65535" exif:PixelXDimension="992" exif:PixelYDimension="855"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8deed1a6-5431-4e06-9973-719a94ef57a4" stEvt:when="2024-09-25T10:15:37-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:196253a3-2d41-47d0-8e52-c694c2a25be9" stEvt:when="2024-09-25T10:18:24-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:dec66016-6d56-4a37-be9f-5a128ae8d7c3" stEvt:when="2024-09-25T10:18:25-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="converted" stEvt:parameters="from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="derived" stEvt:parameters="converted from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e0fa026c-2b50-4255-8fae-7a1c4254e60a" stEvt:when="2024-09-25T10:18:25-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> <xmpMM:DerivedFrom stRef:instanceID="xmp.iid:dec66016-6d56-4a37-be9f-5a128ae8d7c3" stRef:documentID="xmp.did:8deed1a6-5431-4e06-9973-719a94ef57a4" stRef:originalDocumentID="xmp.did:8deed1a6-5431-4e06-9973-719a94ef57a4"/> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>}}�.  ��IDATx���|�u���k&�S�6i��)M�-=rj+�R��"������곢����*�쮮xXaWwU`9�
�Rh�-P���4i�&͡9�d2s?�u'�4�I�g���_��L�ޙLJ��\�����߿_��ls��v�r�=TZUXZU�Uj.1�.mi-��4J}���:1��    ���Hv��2�M9��m�ە9^�V��X^��y[i.).H�[;��d��!���w;�9�b~�~�ojIQ�W0�t�#��!���j�^j�R}����ˬ�]+l���PA    ���:]��3�.4�}���V�>�\mz_C�q3�[��j*/��n��ʰ����'�C��r	�N!�Gg�
��}���w.5�y�7C��A|��r    �I��&���Q��H�Z=�Uh���e�lFV��E�O��+���#r�1�m
�䢴�
w����,�UӹlwMg���?�T�   �Qo�|�р����[�b^3�<s��+�gʂi�����z�O��}D� �A��3�[+ޭ�\j��ң]�~*�    ����*�wUw����~��2�L��'TƣF ��U�n�J7����]z���˨*�    �G����U�癫�|{��´��Ȫ�s���ֳ[Z+W-�D� �ߠ�;*6��-5oK[C�~*�    ��P�q�3^t�9X���b��3ff]pz��Q ��׻���J������˪�*�J7   ��uJe|��y���?�ܾ���2~֬l�o՟V��K����_�[[�_x�m���+vU�7T�   @����l�ak[��th[��-�NE��T�VŻ�#Tjoy�Ͷ�������*z~�J7    �_e|���Zs�o6�L���<1WCyq�[���f�fH�K� ޯ�]w2hU��U�ǊIw�{�P�   �H������Mm�ɏ�o�g6�[{f^��ޞ_O�x�p��]]�U���m�¶����j��    v�W�uǞ�ԪA|�U?#�A�����Wu�lI5���U��Xom5�}o    �����8s���>�F����E�sk��MɊx�p����*��k-��k-���B�    b!�\��5������isM>w~�\�"���Y�:5�*��'[ x�w��ҶR����.�O�    bgЊ��J_��s�ve~�c��DE<�x�9�o��[��|���7    ��)q�#�qW��]0N>|N^�����U%I(������@����<�ص���Z+��Ҫ�N�    �cЊ���`�ߨA���.(,���_�6f��Z{n^�p߳�;`�=�z���_kY�����u*�    �^�*�[����Kn8�����Z��u����$�D��`]n�������k-�ߩ��0N�    à�'^k)ܸ����
�=3�g�/(IP	O� ��=�W/�,5W�t�r��    �*\/�9ѵ�_�i�n��3n��0{ʄ􄯄'J ?e��������y�~�xk��    $�pE\��V�=f�K�w,�v�%��Us���fI�)�����6�s������k���    @��1׌�[ϱ�.�?��ĸO\8����VU]�����h��Õom-� >�W/��l.�z   @��t=�\Z���k�#��,��3p�%�I�)�n�����#]�zZ���    �!\	���M�}��h��s��^�87����5���|k�6��,3�[Upa�7    ��p%||��<s�ם��ۆcf?��K
fJ�[xo��W/���K�'�{�    U�k���͵�7Z���]Z�=cr��+�n��*���<��-�g����7    ���S�C��n��K�>���?W���13�Օp��������4�w[Z�|    8%����7��}��\�V����U�������N�    0��S�_��~�o<�m!�u+�]Y	wK �*߁�1������!?�o    �H�U�����皌�`��?X�Jx�xo廥#4���V;��)H�    �S*��J�O����qE��*���V��dp���|T�7��q�i�r�������I���<�)�!�v�Cޫ�	    D��J��6�f����&��� �[��s�s��?;>_��7��$v��bYf��
3p��M��O��ȷ�a���O    a�J�����i��|��\�Jx��U��U�9�K�����T�U�$t����"�Z׬,�������v�W    ��J��=>��_�g�wK�V�����b�{+��'�4|S�Nb�X=^n�h����`�ן[(k����/7�#�    ��e�O���F��^3^��[%<�ܪ|7��f�GǨ|'��^;�
̑:\�)Y�^�T8�I�_Q"�g�ݿ<*    0�����o�Iq�7�g:z\*�
ཕﮠ1�������|'�o�8Y֞5n�_�}ݻ�������~yuG������r���AC�����߾X._�I�    � +�Z��x����fE~\*�
�V�[�<>�DK��w����`�[��3��#�ַ�|��?~a���/�O   0�p%<[z*�?�c��{=YW���J�����m��w��n��c*�I��������5�vq���lO��p�g �rA��O̲ޮ��˦�M H9�J�W����o��4�_vf^L+�N����}O4�zs���w���S_Oy��f�±V��|�{?Y֯-��s��ֽ�C�� Rϣ�,5��/
���ny��Z ��\s͔>{���ឬ-͍Y%ܩ ޯ��������v*�IL���j���ޫ��=�:�/�gex��ˋ	�  �P�[��<� )g�J�w�l�*��Ƥ�T �|?�zˬ�6�R�Nr���ߟ���߱�p�?x�N��R+|�i3�u�'��6\�����ig�T�� �rN����3�Z��:}Z��p��np/}�����<W�|'5����_������j���n�7�m�p Ha_�n���[�O̶>�	8 ��S*��F�Cj��}j�?+��h%ܩ ��yf�������
��$�jQ^��o�I;�������e�3%KN?-۪� R��j����R�� ������<�b��qE�N�t�nw ��w��f�������f�e����@G�>�k;��U�/3�&�@�y��%��x��kh� R�)���mn͘]�a�<�~;R	�;�k�^�����Ooj]m�=��}Hb�=���"=��o����J2 �Z��az�hC��&�����R���+0;S.���y;d��:�t辵��vS�ȱFs5R��}?����?�bs`VY�̝��H%ܮ �;���.0�g߷~����w���殘~�g77��o��{�l��'� �D��M�y_��H��,����"��t��L�jN݅4_gw?dFͿ��~А����c�JxKG(�П���}jb[�Wj��dv�����f�.=������;C1����:{_�TD R�V��gt��}ц�����{�G�T�,�n&�|�8-;�#�'��.\���H�	C��Q%�u�!G��q���������}�2�Å]!ٚz��w�*���=�^0��|nj�����WFu����� �C�L�hІ�
rDV/��E�EV�u�ϳS�=����#/�cȺ��O�U�4׬'_o=1�4��%�r���MҽO<jv��-{}y��瓓E�z��i�x�  #��ȱ�,�_D:��Y6C���1÷H�8w��d����3=��wT��X���qIF�Zl���If�fd�,��nޯ����pk깿˘����o  �h�}tê���ӕ����5�<��L�T�Gcv��\"�]����l�-�D��ia9������-���Ȅ=v]<� nM=�톖���VS�SR�=؅yi �St����ε�������l1Cww�_�x�{0���ֶf�&���I*/��.+�e˹�r$'+���Xx��󃵁ُ�������o��M��Oˎ�Y�}���< @��}�c9rl8��pR���>��;x�MH��=�3=���B�"�ZgH ��#9A3��T�-�f o���5��N=��k-��~���)�HC@�L���¼��׎7%�Kn �^�.nǾ���K: '\��#��֣Ē3xT^⑿�����z��+�&tq�w/��cyl���O�0��c�����vvT����B�z��ޭ�Ʌ�ޟ��lfN�>�'V��w�G �Rw�y�Sχ�~	Ǒ��N�e�G>|Nj����n��_4�RsBQx/���\�-u��S?�<S+����c����~�ZS�!��k��\R�[�^R�#��@��V�?����_��j<  �8��uL�M;� �uù�Uo7O5�}"\���-�鐫���L6C���{c�~c���n,m ����k�����d�9,�k|V��Χ�b�yL��� H.v96mC���� �����z�G.^L��K_���U"����yC�NJ�	W�+ֿ���ⶶ�K�ȫ��F����G�V�������s���n[� Ze�T��a���x @��ȱ�h�;m� �B���z��?�������N5C�s"��J�jx�tw|k�hzlCˡ���(���bc���>�����5X!L=G�7�_�/;����G�� �䡁��{����]�d��S� �*4�٭�x䚕�HTL���%�/����&L�#�t�T�\���N<�����.)l�1LEuZzc�O~��6zፓ�ɋc�A��¶��D  ��8��{ 8�ј1Y�n���2��h}v�������Hp����-r�����eo�(��G��{�+���Z!L=� |���b�vs H^���=�V�iC	�߹�#�J�c�z�G~|�ȗJ���'�W��fۡ/]Q�g��4�[{�7���4�ja�7  p���X���*8��h���^Ɍ��ˤu�L���oDn�ׄ	὞�M�Y�/�%���0�
x��Z�o]��  ��u�y_+h}� `p���؆o�-�C�b�ғ�������xB�`ϭ�<��9��~��3�_��R�<{��U�&L�*���Qa����]R�g/G�<⸾i��Z   N�G�y_��iC0�e3D~r[�·a�I�Ȓ`(�Z��}�}�_�hl��$M��o�#$�V\��W��ȅ���s�A�^����5+�3'�K�x/�H�w�wO����  ��l=�6t �)�O��2�Нin�u��u�P��T��/^3����XIO��7=r�]_	�������߲z\�{�G
���  1���hC�W�x������̗�P�F�7�CY43f (f�4�q��cs���|���K"����Cx�z��Gz.x$p�~  G�4Co<[���@ظ\�|���kZ���22����ٕi�\I��Y��N�_�{o��aׇp�^��*x�G�+�h/�����  �v��s�M4�?A RZ�W�[7��1������X�����JxzZ�xnM_��#����߻���޽�:�����������  b"|���\wA�<�j� H]_��#g�v6|k�y��<���k5\�x�Dug\��#W���Y׆�޽�Uu]�^�珸|� ��o  w^��kц��kWz�央`����Mw�>���������\��yi�kCx�����G���*���v{���  8DC��&�����T�x��/w6|wv��:���@��:�,#�ɱ�s�%"�!�H���U	�U�Y�v����.��5����dP6�ʹ;  ����/�*�h� �S �������̉_V˹�o�Y��5����iM����M�ȭf���\[�o۸˷�K�(:d|�n_���`�7  pL��_�|~�����{�tg��:`M÷��C�b�{H�$�ʨwd@ۚeݭ�O����^�qw�t3���0�Ї��qW�2�V�{�e�+|b�xq�G�5
  1�����m0 g]�̹}ߺ�[۵��G�������ȹ�����}"���[T�w-6Cx���9}` ���WTl���~#�_Q"nB ������� ث G���\;�{��~���L�Ho����r=���[���
��J��]�23�9}` ���o��[*T� ��ܼ�@j�e�Gf��_�N���S�u_xf����.;�#w���[����6��/�V/5{� p�XO���w���z��tp�"�߲"�������M���{��q��v���j|�.�6���Uol�m���Zz�������Z��o�I�� �BC�����m���~ټ��\�V0mP�Z�� >y���;�4�'�]�|k(��{�g�y䖋D~����}��wl�������T�{��T���7���N�5�F>� �ŗ��n-��t��'���O�?f�F��'�����9Y1�� ��b���5#)��?+�����e��w�]#n�g�o���ʠ��O�n~0���Z:q��󋆬|���U  �hPuS����p ���q7���Hjkϴ���G��/}N�3�̷�Z_��#�?�*�*��2�i�׬�?ez8�X�Ϸ��U�ta�9\��Ӳ�s��򹹃���N��s'�U8�$�����u�u�ç*����Y ��j�G�ΰ����U$!#SПa�[!�ΡlW���ﶸ�
��J�[��ef ?ez8�[���	0��s��b�fe���M;���C������{   Dkł���Y+����">0�[�]|�/ ���귞��
��P6W�����������9���o�ƪE���k&Ȝ)Y���ۇ:�G������	 �L��_��r��+�����9�N~�W֜Q ����ҙ�R6>C�^]ACZ�����}����J���K��.IVKgtW��U�`�`x:�-���Ǟ��.��[���`�[�����﷑vW5���߼q�\��@�2N��Q��?��IY�( �
t��JW�#���:=���yG�.^�/_��D�\�	%�"=�#���פ!�g���,�?��]���io�yW0O}�2��˝.���NC�Q��0�{+�k�u'�T�WW�(�O��0�5m7ߴ�M���Q�T�{�ux2L��7�<��7Y�0_�uK� �\��������I2)2���^(����}��>W�P�x��t]�D�E���-����vTuZ0�s��S�{���9���s�C� `h�YCx"LB�D��_�_X�ǵ�
xD�s��חL$��^P$��wZ��dq����W�
Q�-}�2m
���<o�����
ny��/��D�#�z+�k�󿁘i��o�7ʃϟ HeV��
�4��
n}aa��}hi���Z��^Q�T����]K���脟7�n���q��MV�ߘd��;���wG�F[Z����IC���eO����N0d z�t�����K�&�����ӕ�h%��g}f�^����
"�d���n^y���KO��l�E"�ͷ�����1��ή ����"C���q����A�Ҋ����5���l�8H�͑F���/5ȳ���V �C����	SK��܆���{�꽯o��h_�����U��ǭk�ϥ�t�{u��zq ��4�1�3�SA񸴤��.�H�Ms�ȱ�A��X�s��a��=�k��T��OmtUz�y��er����������oĄY���"�6�������o�ȷ��  C	O�r���Z�a�Y;��������|~�U]�4���k�^C�vK�@>y<S�S�V�wK�w̞gc�yW�3���ϡ\������:�T���ƪ��[�g�9���7_4^.\�?��=�_����5 �@��K�xx��@�N.�{ݕ��N3���֮��{}�A��=��dz�p�.H>�]N�������F�u�7��ϡa���}w��
��,�v��NdU�C��;��/iG%��9�X=�
߃Y;��g653d F)�����kxr�=��L.� �\�����Uu]��>�D���:����ӧ����Wf0D�]��LO�>��dy�n���������=ܪ�W����v#Y{eG�<�r#C� `�m?�h��>\P���cU��g�ĒU���ƟZ̺M�0>���7�������o�t?���t�����{xu}��
xKGhYck��a�ᆬ�ޏ��Đ5 ��VkW,(r�R�FO:0�\���.x�*/}[�-�nw�,�.dx����:��03�'��ĥ�I��^U���߰ͪE�r���Y���ݒLG�Eb��gtk�u�øq����y=���~�N��4O��-���kCB�)�w�����O�;d��'��n 6�0�����:7%B�HG���>��n��a\�Ɓ�[:��^{�eUla+}N�8\_h�����*G�W���HC�t��#� ��M=a,��W׻g�m�Ɠ�x3�N3&۸�� n;;�Ӳ��&.+����,���T��ۯ(9�}�n�iw���ˣ p^�M6��f�����x��͢�$���N(�iF;��<�ⵞ[�7�ӹ�Ƌ+}vM���T�� $g�̑��iN�?�y_�+ ����h���ԏ�K��k�D�x���fq����+���h�C���З���Ք޷��`��  g���da+��D����6��]@���n�����[V�����Otՙ�o�  H���=,�{Z�V�u�xyI���y�<x��9`XR]Q����i'�;ɞ
x�;+������  @���~p�7��ր�v�0���Z���:B��J*���*8R�]��t��]-��b������"#�#j� ���~����;�=ɺ4j��鶅�/�p��p���H]ٙ�]�
�s�|qC����-�
���PYW��!� ���|j��Ь0~o�54��k�G�b�p��^ ('þ��p��UW��]��=��j��p  �T���k�~��ʈ���Y��u��{���r������=��쫀{l�ԍS���j�E�
���|�T� Hj��>�}�w=���6��xm��G�Y"���F��+�S�v���<w���4� @���~�p�}����z���֠�Us��_wA�`p?�,p@�3칎a��ʎSb��[�/��� Hz����O�ie{,!|�ǫ���H��ڲ�;�V��{�|b���]w�OT�p�[�Mp�'(p����Z��Ղ����8�  Hr���!V�����F�:?������#?���7���_g>������M��M�����:vD��#�=�.�֏�t  R��Z���:Pj_y�+�f8�~���hh�=\���i��o�@�`m���|���Up��;���pZ� H-��(5��m�7���-ת��'D ����\�l=�}�Yw� 6E ���+[":��)� �!Y[ӫ�}��q�c��ײ+|��p�^p�z�zh-���jAWV�֝�.������
xG�p  �b��⹿9ܚ��\��dEUqցsv�=�n?���J?����Wl���58�؜��mnW� ��۱�J�������b��+�pD*T�iA  ����;���[�J���8E��~M����|~�맞�[�	�@d�4�w-�o��5��Ő.��  �8r�/\��X��vmנ����6��������W^��{�w<&Ï�ր�;��]y�Ό�����a�s��o7#�  �N'ץ��譡X{��{�Z��D��q���\K�b(�%�O�׾S1�Hz���q��W  cЦC��nz�C���;Xk_ O��$$p;���� @"�j�{�+��Պ����m���0�p�x*�C�+@t���Q��/�1ND^�}��T���ug�H���b��ޟ���ṉnk���9b�n>0�z����  ��p�s���в�vu{�Pk�ܲ��7tj�O�q��������E��t��1 !#C=������G�}P;�a���l��vߐ=����튙�ﻣ��4�k��K�	� ���=�v-j��U�7�a����zҴ���m  ���!{�g���`g���yX\� �p�޼���r+�߶ź��q7����]�ĆؾZ��E2��?� �$�:!݉i�#M�����h��	�a�>@���g����6dA�=Up��%���i�.��r2��gܐZl����5�"�t�a�V��0�A���Se��	q��ΐ<�.�/>�|�  ��m�z��"	�+z��F۴��ߝ�ǩi�_��� �o�sz�ՊnĩhX��^��;	pJ#bl���{}'���
�3������q� ����=K9�+�=��G����[���=�)���ƻU��W��	c�ϡ��:$�G ����֊w8����nM�  �hip�s;!�c��S=D{z8�~����VC�{��wm���m��P�F�`�t�>�vz렻�)�=��-��}�[ӟ�:�
�T� ��d��t���0R�./��m[C���L8��D�Ȏ*C�fS��d �vȱ�·��E;�7���GI�����;1������-'� "�T۹��(*��"�H�\��w�}oˣw/u���Sթx�i��ܾ륧���Ī�н����ic����Qp�^�����+V%�s 0'÷V~#�묕�HG������������nE�ϭ�U'�_wAiTa\��?�t%� xm�!�]c�>p��
��ߛɪ����vq��&x����ıb����! 0�v�T�V'��8"��#ǆ�cmE���N���]+���
��8��l��}~9�p�=GD�0䌙6cKk�`(WB�G��	�^���~o<n��=��{��jI?\�)�&fZo�oc)+����?��|��h�t�1�LGn�ˑg!�j�al���?X�;���k许�8!H,��3��{�4o����GD�+���4Q�G�L�;��J�o@�]�(_^��*�2���?�Ǜ �H�[GC��G2��ƵE\ۼ�����|�
W���������NC�t��m�T�#�D�[��3q�p�ah�y���0;C����̙��{�����V���G F���s�y��i5���ȰH�еr���P�����@⪬��/|�{CxFz�t���`0�d��?�\���=M�!�i�D��=�B���>�pQ~��e3c7m}Ɍ�?H� �ѹ�ֹ�������g�׆���u���!|lm�}V	�x~��� ��݌�F��*�*3�Y��Nۯ���DB ����N��h��?��Q>sI�det�%��"GN?-[ޫr�:p���~���  @�4P�����ik�{4m�}�נ�ֆ�:͎�G�k;����y�f�l2Cx��}�i-���6����L$���o���Ym��p ��s�x,��}�ў���gﰛ//w��8I�����V�b   rZcAö���
u�e�n��k�����sp?'��J�fF�W�q}>:��ők'Z�[���ǜ?�[+�[L��x���(]&�I��t9P�6�!m��������q9m2�й@�a_��iE��W��pmI׀��f��y��ta�W���+ H�cQ�����k�A_�,�����~NU�UzZ���L	�b�w�i[~f�3�D�~+xי!ԩ�k����#3�vI��5+[>�:WJƥ��f[Kw5o=R%�s�˴��<>mE�J�S[�����е�u��^3A��;Ҋ��k'�r���]�OT�d��w,i�ׯ+�i�\�����������&�a�I*�HH�2������oE �������p��Ξ*���@N�6�s�'N8��#|��v�<Y'����M��Os+�V��M�������~�L���Q[C������_A9���?! �ȍu��5�܉I��������w�x�3!<;�V|��)7��	Z_�S^ܞ��oE �����?�Xv��0�b�\�О��P�����zS�B�m�Ѷ�k�9�/k���L��_n�e�7o�,k�:u?�^ �X��ǃ�p���������$ۑ��#9���f�s\eg��jIO�^�9��C��/'f�[����m���\.��N�>��^���3%?-_�f�M����h�����2gJf�V�q�ir�%r��<y~k˘��߶�X.3����kj˞v���(%c��@��g����k�[{�$�U�!�c8³2�%�U(]�<If�iM��f���~�ΐ	�xD {�ߺ���/���͖-�'��J��@2�W%�c�d�h�}�'��o_,�����ˋeW��\>i�����3f����V����i���o�{r�� NH���xУ�x��*8���`�EK�{ӹ���,�`����������:;y�Cy%q��*����o�z���\}� �$�%���r����m!܎��5��.�az��\k)����N=��Ig��@2K���x`�؎7k��9�Jg?OzZ�x=]�i�p�H�(��tZ-���rگ�%v�V��]����o�|/�71f�;��(���)LӶk���0��a�~�V��/�u|��C6�ns��q HV��~�Cδ��f��1�HpZ_1���y�sUp�U�,�	���ǔ�ߙi�"���K�	l�#	/���6p�t�N�/^^$�{]!\�d�6�+m/ץ���,���<�w���i�:� 06��~��z�p}|��O�3d�_�L(p6��p=�,ʑ�`���I$Z��j��X�Qeȃ/&~�[�t ��s��-m=���供�K<i�K�kK+�����O4m�}�p6]W�(����K���S�����>���G:�7N:r�8 ��Dk?�}�:�<0H|��j������i�ե!\����pm3O��Y�;���!��$�����X��fE�L,��0v��G;�m0:���U��eZɩ���t��4- 0�Dk?׳���D��� $��2�L�㫜��������Cf�oR�GBV�N���wb[�����~I)���j��Z��qd��~�;�C��
n=?/��h%��J���
��Dv
�$����U��~�-=#�Y�<V5\��ݠ���j=�X{}�!�|99Z��R:�k�u���}����a�]gHqƫQ_��6t @|%Z������-�	RUf�\~�GC��D&�.�+��S2�2Z%�4o�b:��#��|������K�Vk����U��6���rh�k��az>xa�6[� $�Dk?�;�LCx9ǧ����D����a^O@�i��M��ĳz*��>&�if����ѳ�Ր��0C�$���v��~z�T��<wV��|��4���p ���<�*�a�@ $��w�|�qC������0�'d��wOo��q#S�H�z�лou&���U�q�qaz����6d�n�nrǿ'g�V)��������*5x��-�I �d�h�������7L$�����4$����o��o�K����_����{�������?%m�V)�����s�d�u�\�|Bl�� 8+��ϵ�|�Φ~�۲���g�H^�}ݐ<3�����=��	�a��qr�o��<�=��{v���Xǋ������� ��K��sb6� 3}ߝ�Nڼ���ِc�zFx"���󹟄dg�$����6��lw�ǧUp� %�j�y��k��:m� �I��o1䇟�
�׾��!�u�R6�GK����N���ʩ�@�K��s�7��ְ���Z�����}"�����w�G&�� �v������?))� �|��.#�
8 ���瑄��k�82 ��N��W�Ӑo~Ddv!|,��0�[��디B   ��=�j��`{��r�}oˣw/B8�x�{D�+?7䋗�\v&!|4~�ΐ��`H*"���'k���Ͳ�G ����~�U���<e��H����ZWV��K�y2
 �4��U��L� NI�ϐ���so�f�V)�u�y4������<��A�' @�rcPm�{���]_X�
�-}Ր}G+�Ӓ>��Ն����վ��R6��!'����bq#�~ �P5t7�|4hE�6[�����!��L䊳	�}�q�!?yΐ�vIy)�k������c���&n���ז��P����s�Xk۸����ͭ� R������!w��r�ȼ���w���E^ޑ�-��l �nȑ3����)'��J�,��=_Y6��޲�  S<�V��ذ������m4p����E>��#ii�R�A�_�3�ak������[L��Ϯ�������ϕ�l �ڴ5;��ٱ������xɐ��3�{��S�������n�`)��j�>x�����&v�������J��R��)i#E=r�#Sj[ݳgt\V@&��%;=(2¿ˆ�%6�3���=[C���}ʸ�����!�ڙ.GZr���8k������=���%�r�*w��@_D��+CΚe��3=������"/n3���l?(F����'D=	]�͚��ǭ�劳��-�3^��Z�iAOj��Ip5<�ԑ!�.��O-)m���6�$�k�F3��qd�l�/�2c|���� Em����}�v�H6*��7�0!�S�=�,��<�߿�x�l�*��gh u�B�@:ܭ��G%�k��_�!�m0�r+����M�0^U��[�Of�>� �@�p���� ��sM ��]�9�,9������W�"���ĨjΕmG�dg�8���?"'���o��ͪ�B�3;�H �j����<s��V�?0��)n�g���-��`L<)W�?*i��TY4�YN7���e�����yJVvp7�����Q���y���EV/9w��9s'�w�y}��k���;�������S�5����m�ߔ?n��ng�[�$�f�h��1���
ۭe�]S$��}͚�*ם^#�yg�ĊV��	�}����������ӭ��X����Gl����W��OmG�ߐ/�ז]MQ�d'B�HC���r��s	� \�x����2�}-5� ���0���}a<3t���!���(��R:����;l��V��Ծ!u����������i���O����i'd��:[�u���u��w�%���ܮ��Up�&o<\,N��U�|�
�r���1{A䃳���P>d^� n?�w^;}�!4C�@��W}e���/@B�L�/3Κf�R3�/�0��t����	�5'�v@dG�ț����m��n����c��k�s.�����.��px�R�a[��]�jUs_�r>���o'hK~,�YS��� �����V�eeM��o�� ����E{�t�����KF����NK:�D��a]�������@���Kg��))�L ?�`Ȟ�"�+���!kH� ��jCW_�t��z�j�iul+�Z����G[�I�yrY^�Lp]1�l><!&����z,�"�����mr���m$s���PH[Ý������@ �_u����S��!T���o��l}L2Ӗ�'��F�B ���ú��ٙ�̘$2c��\b�=.�|���HVϭ��#J|���ݓ�}�̷����ȡ:s7��;��)�xi�\{v�-Up��-+��{�/�y�bS��m��0}^�t�����?=�jNI��+����_y�w}3�;��U<;}��c5ѡ'b�9b��S�V���d܃��B-� ���պ"�:���pF�peg�;ȿ ��DVΟ(NҶs�+��G��2)�������^�«�Ls�(����`#9�΍���R1|��/Dh�=�  �B ��acvU��^�c�'Ol;G�Y�T��������גKV���&;�� q�>w�n�  ��&6fg<�3�"������YsJl�fxؚ�:A��_ $3���޷���Mg@  ��=쮂�-�Zo�gdwm��X%3J'��:No����� H� �5x���a�&��<yJv-�f��KQA�tC��O�#Y�cV��|�0� �j83 K�>윈>�e�����a�olϓ�@��fy%'�#i�"��6���q?��|`�o @���p @,���g����oq4��5>�M�K�ē���� @*�% �4� N����7_,   ����zγ � >�p+v*�p�z�y��� ���%}ˮ&����W�7�� �����!|�����IV�� `hO�Z+�v6ˣw/�(�?��V  |ښ]>�CV�l�d��}�  O�ז���׊�~,  �!�� <�-�B8� ��	h���+�q��?����; �H�а�ݏ����o  �FCv8h�8Uo �h�#���Gsz0�\c�7  �#x Ƃ >
^�����X�n=�[_@`�9    �|�4�j��>�NB���    ܁ >5�9V�����%ݍ�p��    �.�(<�u���%}Ŭ�q�z   ���m���f��jx<���'�N�*�     w!�ۤ���[ik��X�������    p/�­�Z��ܼ�
�]��p����T�    1�����R��p W�P��
�:H-<D��    �� C��\�t�k '`   @r"���    �    � �    p     b�     @� @J;cCP �A   )�������x�j�����/8  HI�o r���X0:?�� � ��C���L� � @J����ǛK �t��L"� ��A�+�'e0  ��7�X���� @��в��?A�[:9�Al�   ��@��1� ���   i�ē߶�@!��   )�1��?����(�;��vH 8  H:k�0��M�o �`Z�|��2�Q�!���Kmc�ԟ��&8  H*�o n�b^���%]u9f�ڦ�u{�1`����>��c���1H>p  �4� Az�G�K2�5��k�|�a��u�CvT��x��DG   I�3|�_�7�$Q2.�Z�g��Y﫮t��J���ɞ� �� @�#|H��猳�h	ʻ����/��d˞v��� @B��L3|�� ��ɪE��R�uʆ�Zeûm�n�O�>p  ��.5���G� ���LsM�O^<A��0�x��[�p}@�p  ��� 0�e3s���kU|��mV on
� +f5������=�}U7�H���r���6  x� "��\�0�Z:Y����"���aם]c�.��`���H|��	��֩r @J���O��Qөꟻ�X�<g\oo���C w���h�@z]+�kޱf�l>0�
�z�ټ  U\v��o$|@4�&d��W�ȕ���.C�<��4xk@�#tG���ͷ5�?�u�ĩ� ��eg�3��d �㴉���&����Yp|�����=�����/&� �� �3�,K���I�zq������0G�9� �x��n��E�����VU �d����$|��Ξ�+�:-[~�\=�p���@�vk�y���&���A\_��oS $4�7 �V~�ת�/0��}��
�u ��2mbf���G��W?��5�ZQ(9^��G�5���io�n�/���W��t�� �D��l3|�� �p�9�d~y�|����v^T\�s���r���G}��.,꽎N��{��M����mAil}����������|'û�������ʪ�p�� ��f���� q�{�_��9rۏˎJ�����\M�:j���������o��&�U����z��Sߟ��������
�������E��?�En��rB8 ��� �.~i�|�����D@0j-���ao��DT|���~�_x�eL��[�v����m[$���pB8 ��� �N��B���A�k���V�u3}��Lo����oī;Z���:{�?�0~s�%|���T�W�BB8 �u� �n?�s����*insoխ�Nɔ�W�G��o8>T�)v����A߿jQ�L+�轿��3%K��l�/B8 �mt���%|���K��>Y&��#��+���PN����-��v�V^��7``�}��lG���N��F;: �-� �8��̑�{S����!��~o�}m�+�N��a���9�$���H�'�&�A����r��}�ݟ�+9�L�Yg���w"|@�`a�|�����ߎ�����r\m�}9�`�ڳ�H�pqE ��t���У�R����Ϯ�^�-H^A��Y0��t�=S�T���v��&_�������L�P}���_ՙ�c\�3�Oc���>W����� ��>��P�g{�l��.�G��{V��>zۥ��{��*����>���ic�N�xW� w���s���:U�[r��ȗ�l�t�%'�c�i���&9�2{b�,��c����!<1>9��Ԙ��&��,�;�/���?@�����빆F�˴����}������~�x��E&���	ێI��ٿK�����؞a��kȓ���q�f\/HW.7��G� ��>zA�}�ʷV��O-N�s�ڢp�#�AQ�������b�ثS}��O@�5m=�Q'h�>vr�d��̲	r���a?>4���9v�JΜ��,�v±Ǧ_�>>Z�Oס'F�s�s�vL��$���KWu�r+o��&�D@���pނ<����ӛc;�:Ʉ+����>3|�2!�]��*�斨�����!h�r���N��?=�} �{�j��H{�Z�7� .�3��E��H���ӧe�K+ӳ����R��M��;�8iE �� ��V��=����|�k�m��[17[���E�JjT��m���q���,˗�8)�U�"�����m�����}\������1G~��L9��מ�-њ9u���ӭ �p�k2���V��  �}��� |@R�_�m���~�QRT����g����y�T�â�f`�_���%���G��c������c�����fe��?�F>�&_�A������	�N�. �� ��� ��4�?����E9��R�^<=�j=�A*�aQO���K�O���_R�#�~�L���$���U�U����ˋ���V�v�E\=��^�i�vy�/�d���5+,�{��?�g�U|��Kj�vl�?A  �ˇW�7n�$ ��s�V-̓�o�}15��U���o_[�nv�g��wX�)Q��Ͽq�_+�~n��Dn8�H�vJG����,���;�����Ay��ط-\{v�m���b�+�y��q2�`�m��V����� �q���N���w���T�z�M�t�𽷯-�7gJ搕�0[ʴ�~�V�gX��4h����{�D̫�:�ܮ��[��c��BgKk���g��zZ�煽� �h� u�D����r�X|N���o3W�ͫ�����ܽ2L�;̶>�/��Z�y�d�xI�dex"�}Z������f�5��;v2Wڼ�"���+�+�In�=������  cE���s��|3��;�څ���$ݕ�=.���W���f�Fe���d�_X$�f�5xo;�a�����}�/����ZU��mh?�i�o�D��rx��CWHg��(�-�k���fS ���f���� )gբ<���&} �C�u����3^���E;�;�G��Ԩ{�u�O�/��?�������R���z��~瞧a����.�@<�̷޴�z�hC ���+��}=� R�Iv��\ٺ��#�]"<�\�����d��k��
>����eۡ�����Yѿ2s�9G&��hΑtc���Њ~�Y5LC �
� ���y���S�����[Ϙ��E��7G:l,Z{�f���4q��wy�Up�� )�7 @-��D�S�]�2����Z�uhJ� >զ�����;�K�����p�� "u���F� Hw /�K�涠$k��Y��k���h��vDS�J� n�����\).pO�;L��#_2<ѷ���� Om�*  �� hIE��7���.�z~pRaڞ����z$���d �þ��RV*��M���= �������#| �[\��L<<�|��k�^�>1cTS�J� n� ���)�Vm�9�oC _>�
8 `pך��o	� �A,�H�}����>���+���zΨ����܎=�ǟ&n���r� C�N���6s�������y��'Ӽ�0o3�� ,�H�9R��{o�p�ѫ��k%|�S�J� ^e �=�+�)�f�>p��� ��;I�E�G��#b�.���m��g o��ѧX�����x�@j�Z�!5'�Ϋ��|k�{��g�����W��H)�������
4 �f��<,F�N��*+pw�m�^d��^�w���>ϸ� �>K<�ͷg�a�P $�������������ͷ�5W��a��@I�o[[,�f��~R���ԑ'�j]F��{Z��F9p @���-��s-�;!k��3C�.�vww�;ތ��cѵ��`nU�g��|�y;���t� H�L��wyI���^e��}�:,c�z>P��V�EK�e��ʈ��kG[uF�e @� |'���b����C�zZߍ����������D�� ڔ�ཕos���G��O(H����P|բ|��m~y�����5��q��t�mF  )���b���%o����	��	5������Af����4øw� H<	T�W�6׮��R�vY����0�pݫ��Y�seR�;nQN���T�h��UucRL/ ���f��*��]BMݡ�\��:iu�C���wW�5�g�+LYǄwd���|����ϙ�m{�;̕���e�eg���srd���ƍ��DJ�e4��K�ۥ�'  $���-2��D�K��Y�s�s�\)$�*�����x�.4������ �Yn��_0;������<G*�a�
��*���l�3%+���н��'�tȃ�;��I+�]�;'��Q�V5T� %]���!|�B8x��I�V���k��_3�!\ø'W �SN�돎�W��hq����*p��� �`>ojvD����5QV�Uп[$�lq�����\���  ��3|����ඎǺ�x�"Αf���f�6��R��>)c�=��h�;,.|���tk�\�I�rD�z�]�M�p H)�oV�����H��� �DO_#�}��GpW��U�u��s�|��,��v�����[L��Ϯ��S�����е�ܮ���� H��83|���3 z�|�S0
�F3�?n��d��pg�"�jFsTt���Uk�����__.ݗ��u���h ��G���!����Iy�ʙIgv�m�w��箿��j?W��� �p���&|�M�kf�~��X1�]�>1Z$�y^wO�& 0����P���|�dwyq��A�;�� >�	��}i���axY�v���sM\+߅�o�r-� ���3|��;>40j��	����{���������L� @�D��U��n����Һ�ݞ��{v��]{��9������vu�[���SWw�]�U[m��UA�(B�(�;	�g������0�Ʌ��w����x�H&��fB2��|��/�/hm5C�u"%��� I+�'�d��O>T�rɂR�*�I��L'���G�>;�6t�*����'�4
 ���=b����"�r.�o��hK�f7�x��"�%`��u���c�/(�p�����n?��x�̽��ٱ\��
ng�[�� 
��#�VZ�Dw
\�C�z���o)�=0)%��k�k]<�x�����^<�����LҎtFekK�<�B��{�'�4�=׶�܆����r�g!\�����v>m?g�7 ���������,F���\&9�������K���@� p^_$.>��O��w5N-:x�g��نV�a�wtP��a{��^�pm={��jC�(���=��95�Ѷ���s (\7]a��	߮x���<4�Q�����^�H 8�hg�뇐�|2�֪���?�o3u�1�|�^�͒���/&�������;���jCWs�^��hPND/7i�.��=�8 
��Fo��|�w����o!���9>��ʷ�������ܵ���ck ���W-���Oh�����[��M��Gv������BW��g������mL@��C��@l����}��!x}���� ��G�<�)�o����_5Z!�<\�z>RN�����`ӏ-�Wfw]7Uv��o���]�d�����6��U��p'·�� �����y·�����3����3b�(�] ��Xg̫�N�|?􅙭e��+�I9𻾿�z����a{,Zo>��:4�k��s[�}�>�>3p�Y�f[\M+?,'�������N��d����_�Z�~��s ((�oDw���m}G�s�_�?!���j^
 �x0�{T��?[�2sJ�������w�--�<��\Λ[*^^-��d���1�;�M=9!��amvW�Ք�^�ϟʑ�2T�{5\��Vם�z'}�� P8n���7�]�a������V1:�@�3� {���� �R�����Z�i(�M�;��5��*G�+̀}��
Y��\�kƾ��j3����veZo��.+��m?w}�a��G� n�W�A�2�0^�%e��Rrv�:���c P8n1��=�ow�,F�?�P��'>'���%� ��} "��[>�����׵�XP��w�#ې)�h'��7�����Uʹ�K�
�X��q�{c�<��˵0~���C��lk+�p� �S�����,j��ޢ��J�(�c�]��B���S���q˕�f��&p��O��L�ߌο�@�W�'c�@�\.��T�?wݔ�,+�]�;ɱ >�^K_K�ox�Z�Pbk/�9ƿ��G�N�v�},����Lbw�x�� �����/�����j�V$H	�-�o.U����5�V����J n�z�e�J��=�d���jk[�����:�ݜlE�+Z��p�=0�Rb�o�����"����AC^����]�T�ol�h��k�}[�Nr=�'_/�a�c�՜q���m�n���
���+���q���f�͗68֊�'��@�uU����	߮��)F�?	
�џ��W] d���}r���-�FU�W--k������|'y��9�m��jθ^|x���Z�����zp?��}�7W	  ��=�/F�}�f�W�_ ���|�;��}QSI�_�4����$_��Fo[����Ň�1nW o;Y��M�
2�S���A���ѕ�|��#�.Fߏ$P~� ��PԐ�v�9vzQ�^2��������|'�.�7rx��έ8�zq;�hʶfE[��p߬����	3|���:�������$"�#8]��	�3�B��!�N�R�^�X�����>o*�I�����5=��ۚ�ɜ�Ŏާe۴��`*���7� ���F��[UQL2����f���	��m��H����w��p���ϫ�wR���ů\Z!�/�w�x�4�p��yh{=  �}�*3|�����E�LNF�#����E+�w8R�N�|ϝ^����=#�*�Iy���^�)m'��oޖ�[�i_?  ��={G��G�X�-�+� �=���Zn�Q����gf^V���:�g� ��$C��mɫu��>v�<��Q  ��f�����>c(���+��n����7
��v�ȣ��ZFT��kB���̼�|'L wK����x�>V�{@A |{G���)�2�O���/ 	�n<!��U��W�������`˿�����|'����V���؊6������h&x@!|{(���� �}�.��y�L/��+�n���+߭Ue����ˆ��|'�s���zh5|��vσ�V��B (�]]+w]G��D�U�F�c�g(�M�����O�u����ˊ-O~�A�x�W���6Э��qm5O�  (,�oo���t0��:������LV:�k��>�N�R�.
Z���F�|��|'�m��Z_���Ѫ����hśm� �0�=�{}G6p&V�� �ɩg nW�{T��<Z�����I�T�������5��u�f�m�Ƴ��7�I��� �����Y·�4XzC$�^��*&�z����J�|������1��*�Ip��
��NLC�/��?�	� 0��} ���#mV\'���,^��'���=�ӌ�|��-�~�0+�Ip0� 0�?��߫	ߞ�������yVe70�ßے�S*ߥŁ�g
p��Hp  |���3��T����g�@�!@F�E��KEBg	P�~��q���@.�U��(����]�N"� ����}'��{��"�_�#�A�P�6l�G6��"eJ建<���
��D  �C�o�0�7�����_��[â0�w�rm=U������_N��w  ��}$n>��V��E��(��[(D���m�yJ�{ju����g֤�|'� ����?�0��7��mL��pJ�
���<��K��ԙ��GU��kB-���&U�;�  ���>c�y^��Y�K$P������O��)��Y�E���g3']�;�  ���>�k��G�ũ*8��"����{?9*�}�ln>��={jQ���o3'e�;�  �K��D��2�OV����4|o7�-�R*�gM/j��{&o�;�  ���u��#|���"���Ut����_�.?�ҕ�M����d����~nƤ�|'� p�ۿ��ݢ���h� �h�����Y��d�{�y�.�n��]3&}�;�  ���>G �C�ŝ yhϡA���d5#Y��5߭��������YO�{8l�ɫjS.w��sٮ`�s���_�|/�( ��O������K�w�� ��yh(fX뾏tF����5�-��)n��3�T�G �����ȴ��=�����y��J�u�Y6�l�����w��w�<" �G�o�����yH+�[[�2�٨��ҳ�[���zmA��=����������ٯ���e��^^=�������j�ya�|��T��ʧ�5���߾G ��hCG>y����Yu��T���U���OO�q�cT�G �#g��-��%){zsV-߸c��ZZ��u�L/���>K���AB8 _�c3|��������#O���W�{*�uߣ*�uE-f�f�����+�T�\�����wdu�;WOM;|'i5���̐[�� ������.��=�&j��ڎY뾳�R��^j}�O��{"p�����Y��h%��+jG}|�����\��]C���WZ��$}_?�K�; ��gb-�"�B ��i��l(����|�V[�垙���1����Yӌ� ��;ٵ��s�4)	R>�����i���>7;e@ۇ�W�x��g�G�I�F�U�J ?�����[���,��]Yl�ߟ��QV�+T�'D G�j*B)���zL����v����3N9��������$����V�W�ض� �����<�-�k����~�R�<��D&7U�.-���Ե̝^D�;Mp�,��N?��ͩϻ�br���^�Z�5=i�٥p �ѷp�v\�>�Jk���X�R*ߡ��~��u;�/(�+T��F �������me2Yh�{�zn��:����m�J	�f�  g4�M Wi�>q�+j������M�Ҧ��w��Sw_vn���]��m2���r~����#��p���A|{�0�n�Sg�_h�|����ZχӐ��OV�G�� �"vP$μ�ˈ�@�U��}O����ln3]0~����}�2m'��!��4t�sm���x�6z�lJ\����5�on��Ƿ4�}������X�:p  �cD�~�!���_��/_���fZ����V��C����**�Y"�8 �Н��M�֡��a�	3�o2�Wa\�}'Ct��\��  dL��n3zE�fV	N�+����U�V��U�͋go���)�K"�#p��n�kW���=ƕV��_��� ��3x�}�D�~��������  d$���!��pxf�A�社�%��k�i�,�2÷N?? ��ߺi���{,��p;����D\C����V��tF�~ �#��#: �L /�o���'���,9�\�n<`���ų��9!��@[Ϳ}��&�j�!o��hM߸�WV/?����ҚN~���[fHI8����mv�,ë葡��9 &�8K�#~@�O��}��ln��z���+��~��r�|gu"�F ς����m�Z��Hן��F��G�w4�o�ޓ�\��5`�ãB�V��r�����"�������ƕ5)����E9 �8��{;&�'bt��}�l�G6f��$k����-�����3���ie��;7K��	�i�����ְ6�<m���#��5i����Ζ����������\pv٨ʷV���xv����.M���� ��%8\������~�L=_si��o��ۄ ����ΆVõ*~ߺ��_���_R��\�v�9�g�������hZC��r�⊔˻
  c"��KF��=�%��<{Lz�������_\�����ۈ ���>���-���)�ʩ��u}��o���^����Ԧά�O��'��Nҵ�  ��` �?@ �+~��vy�5�-�uM��p`��.��+L=�<���4�7�owd]�V����A���M�����Ϻ��÷*/	Ȇ���e]I L���1�Y5p������e�����43,�|������!rN��?�a�\��Rּ�Ff�I���Վ����7&o��e���y�  �68<G ��4|F��(��{o}Mh�K+�z� �b�N��+�g���:}�v�$ |� �Q��~��>y᭬;B�k�_6����U!�~;� >�V��;)�&ܩ�l  �
�#��A�}��K������ztaCX��{��ߎ ��A���i�"� &8<fC���O�w���ϳjI���Nu
|���~W����Qf���o/��u����]���hw�  � ��cZ��#����%n,����~����畱��A�t8��4��+����RW]#�4KmEH�JUYP:zb��3.G:cٵ_���ʳߕ�)Άq]�~��	� ��E ��3�PW���E~�x���;����+�m�=��5a�c��|����}�b�y���7�NV,-��s��ʐu$F�/��!y����=)��:���ڮm��� 
^��f��w$��.�[k��C��{��ߎ"���m����vz����[(+�i�E�ͳa�\�Ϲ��D�Ƿ�Yu�o�5�� ��('��S�@� �|�<~w�b�pˬ�"1��	��1����g����Mr����6�6�;'^����2���'T� +PA ���@�t�ʈ�<�r�\׀�bq�3x�
E ���:X�{.�[��/N	�^"��l9ѿ^������*8 �`i�P@�+� ��Htwʇ�ր�������ߎ#�����M{�do�u�%�ⴁ�,���x��RWn�+�T� I+���p�$�)���G8� ~j��EM%{��߮�����V���N.]�|�N�U��AN�?c[%�*8 � Q��ఇ�z?6���S��/=���[�"r��8m�p;�߿޵RV]�^�N�+Z.}[��ܞN Pp�px�!l�C�]�1��*�������-��i��?(p֤�kl
��y����=�sdJq���+���y~�Ⱥ����;f��|�G �QhA�稀#w���������!Y<���2������׹:�U.�f^*^;�X��.)��|.�]�>鴡�ZZ)  �^��W�� ����R�)�x������o���dRp��Ϸ�L�	����R.m9m� �BNC ���5��c��z~��X�dN1��]4���f���=�f��'~���U�W�8�{<�6t  |/8M ���p�D֋D�<�U�Y��f�pm��6�\m?|�45��t�.���ܫ����'E�9rbH�T?%,%��< L&px)� @֌����	d�|JEP�u}���J��e���u���nj<K�F���W�4�{\�N�p߷|�]q�#y�̙�� ��5�}�w_(,��#V�yl�Bu�-����ۖ�+��~���wL� nG���C����KQ�WYw�|�F�� �Z��[<@ G����_H�q#��T���6�Q��&m �ì:�~�"�R�=�77��[|�c @���H H G�t�y�HZWM�����eg%���{�� f� ���
)�U��ǎV}  |�u��
pd�H��m]7�5���4�doz�M� �kk���2�*���cc���C�t @!	؊�����S���V��O��ƺ"������s�E�����gZ/
t�t��p @!	�+¯6���\�aD~���������"�������諐�j  �$4W$`�7�pK�h� �ʷV�3`d�\�:x��#f ��9W��������~MEH  �ş�[pM�
82����L���[�y� ���r�K$u���ɷn��rzxđΨ  p&��Eb��]��龵�/�z>�Y��u����W��E �RMi�􈿕��f�`GT�L/>u��W����;\����JI����`\  8#ց�M�qd�Z���gz�8�7i������M�蓞)x�u�ȾcC�<�w��3��-W,�H��/  pFZ����i82��;��s�n<��͜
ޤ�v���v�m77�~'m��'k/�9u�����R_ �  ����A8\@ G���\[�3�I�yC1�+��+ߖc\E�|;T�2��~�gҖF|��k�u}M��Iׁ�ц���KS>�/  0�@x��pT�|��l2adY�N��\wQ�m��� �@+�L� ���LV6�v���	�4��ش�{sk]Z�{~GoJ����x ��y���4v}1  �	��Ϫ��-|� �mǢ��Ҩ�[���ˍS��
<1i��=u�vE[N�h��#m�K|ن�� ���>yD�����t���Y��9�8��}Ͳԯ��{�� H����x����8%�@�L����m����uE��zd��tZ�ӡA�'� >���εiOzp��*�����5�V8�����>+������޺w @��W�A �S��	�%@���͈���x�5�ya�~�7���<	]E#o�n�F�M��볩5� �A�yaYʖd��K�7���1%�wr�y��]}�� 2S��<�����n�ϑ!C÷1������*�S*���Ȥ�ʎAl3*��]��G��]г�����ᳳS�ӫ�W�R38��ώ���\=U>ziͩ6�$]��ß  2(^.N���̭�5�5�U��OL� ��V6��|�pl�zg�b-�]�o�9��wқ���~rT������p���Y��@D��; �m�;�+�Vʊ���~�#��I�d�t� �(��f
�O��#�Q�|�P� i��co�t
Øps�Sk������-�rϵ-9����Wzz�6Ю/Mo�u����-��vOm���u��Q��%֡��uYd0.{��ڔeVm��T�F�~��_�<u  d,X'R�,aK2�'�/� 0�r�����ޙ�\[��X�*^��hPND//T�vY�]��8�NCq���|��)kKV����3�V��� �U��r1�Kh�H�*2bG ���~���:��'m�����W�'���Vt�Į�o;��%W�~�w�w�v�t������ `�V��|�� 9�������iCo����|�
x^��\۬׬h��
�*��Ho�z�B����?���Z�ζ�|,<{�:tK�e�J��L�5��[�c�9 �nV� �\�f��KW
�	c�u[�7��`�peg|JY�L�G��Е�OFw"|+;��cI��[�]�T&K�*��ʐ�V���r�}H�=2(o�� �*�D$2_$�*@���ȼЀ�,&2��-g"���$���YW�>�	/r���s��pvV�Ǣ�㴏 |��r8����odN���c��� ���$���YOj�|Mt�ʲsm��k�)z��i����p� ���6���'�G�T@�w�B�L6U���@ ?���I��K����#�B�FeVq޺Ƿ��;���  �@�H�e"? #�vv��F��H�nx~ ��D<����gb����L�ϑ��,��X�\+��K��k5��7 `���(Ft���H��:3�O #Z�����t����0Z�m��.+����)%��^��{=��<�Ͱ�M{��	��� �?Bf��A���	����"%�
�)��귢��#���f�͗6�ފ>���^񊶞��  $�'x�D"�`"V�Ȕ�ok��"�������򭛶�½��/  8ͪ�mc ά�*��22m1C��������6��9��O�5÷~�����乭��� (��D��g������Q�s��@ Grx!�p�fǺ�UK+�c��Aټ���]�� �%W�D�|Y����E�3�J� >Y�Ϡ�C��f�{˱9Ӌ���K�����^yx}�  ���7�1����s�%"T��-k���OK ��	hHm�헵+ڤPh�vr�wI8 ��Y�mW����y��NZ� �'4We��A,�
�{�&�f�����
x~ ��A�ꁎ����k��}.��]]��sʭ�HgT���K�:  ��D��n����wh� �2�o;r^x~ ��)Z׬h����=М����|��}���ղl^�,l(�z�5E����xco����_x��  �w�����I�I����s Q��ϕa�G π��M{��n�2����6L;�V�����Za��%V�O�E����Т�����Һ޴����c���i�*7���¡�̪r�s�ho����I�k�$�Ћӝa�p�t���́�#5ʑ�R|+8=ъ���`�*j�������=���
x~ �gHC���\e��|X��za��O�\���<*d���q�8-�	_��^�(h�]�w��I���F�y�J�v��n��b���mxg���o�c�)�O5�:v�]Ǫ�7s���Ln5�~N�?��Ņ�Z�e����_	&�`"|��I�-�NM ��,i�}rk�o��Z����NU�ӡ�dU[���}t����[�w�ȋ;{iQ�A}��/f�0��F �Ξ?������b�Í������z��{���
�E�ȕS�<?�s���lE�5��/A���ηeo;i�����bW_̪��Eג�q����;��7z�M��̕9l�>? �J�R����f�'lPz�y��C�p�!�ph���� ����������U���%����ھl$�X�E�S���֖>y�NZ� �	5�!�sbt�|��-(`��@���������ө�ҽF �Q2 ���n�F3�;�u����{�j����wX��s�T���l�0�-꫗W[-�  Oi���]_��+��}� �q��\���!����0����z_����m�[;¸N4��o>Y�.$�0���~�m�hQ xNCx�7ᅨh��?-���x:-�aҟ��'pX"���Nk_��n��l��x�P������嶎�9ֶf��d���Q��E�o9,  ��^x������!��.%��L`x�h[�d�: �*��+bt]��$P�=�7�ng�!�
8�kp䍑ۚi_:�t��8  �*:'�&\�!?����w8���2��T�#�#�$��ͫ/w3  \Wt.!<_�Β@��p�1��������7�����Uʹ�K�  �J���m>���2	T�� ���9��p�����y_MZ���/&;�G���� �p3���d>#>!���%P�'8.�| 7���8|e�Ak#���_^���~�  �^�y1�~h>�>(���(�E ��͟���4x���98<7�Vc#���;z幭]�&� �;E�����E_�D��� Rr� �p����	��������˲y����d��o1ONB ����%P�Y��B3�?!b�;�S���;t� ���w�n�iA�������j&�-� ��P�	X!�q���(���kp�A������)ᴮO�9 � ��J���D�Iq]
�U���x¥
x�Nx� 	�sp8"9L���imF�9 `�(��d5��"�7*�"Q��
��*�鴠��G �m2�2����^yx}�  0i-�@ս"?c�i�s��F�9(����x��q�hA�p����S�¦2Y6�,���;:(�w��b @�u/K����6(���o0�Fz�K G�T�V��@ G�n��n��h���{4tw�b �p����˚�m��A<~H���D�.Z,�o������@ �ch1  ��@���jx���b�4�$P�!����N��{wE</��u�Wo�������<��7�����*i�qz]������?��T>D�9  Y
�H��6��k����q^�Sh��/)6�@� ~d��Y���T�����kS�oi�·�{n�6��b���s�壗��C����1Z� �Qr�,��F~��wb��4t�O ߋ���jA��9[�EM�A���{������w]7u�-������4�Q��>��78N�ǟ�  ��4C��I�<d��D�.�����^"@ވт�T�p��òV��2��|�ں���NZ{Y����>�7  .(�����D�6��V3��G����_l�n�� ������т�l���.M��÷��~���z���ЎtF�}�s.�S:�:�_Rͺc  P�tq���V7���h C
Bp�H��f���\���� 6eP���Ʃ�˯����<������i��?���M�)��U���M��p�;I��񻾿_   
Z��ZеХO��WE�-�w�u��aV�����{1w;siA���ڊ�v��w�f|m=סj�i+�W<8fU[[����r���O}lQc�u��  `������(��|�n�p#�j��7���N��|�DE�Xm���+��px϶ >|��N��& ��������x.���^QujR�V��XRA   ��V���% �"���
���a��u�F�ˏi�yL����#pcR0��V�iA��NAO��e|�Z_�(u�7���5���-�)[��;�T    '��0�S4�k�#v�
GO�Γ�{2�G�|n�d�Oz_f��%whz�-��0��Wg2�9������Z��p"��j|x��Z�|Z   ��a947q����H"�[�./4��%�k�I��v��|�Tǫ~o�ޓ�9�<�_?%,~�r~�4�&�57��y�����=u��=�~[G�   �"P�8�V d(��d���`[ �uߙ��=\.�ﱌ<�|lE��5xϮ�lB�=���0����T('�   ~c��4���u�w2��6�+�V�\��+�z��=��P�A��u�   �_�\���Ҙx�>��l�{��W֌ڷ{,|m���o�i[�=׶�Z3x��
�wn��|K��	�   ��\�~[w��l��L��[�M����^6��|l������5�q;x�E�[������q   ��T�l�<{\n���Zn����S���E+��_R��Ȑ!�f�m�F�!n�ן�`��}�m�*��K�j�V�	�   ���pJ���u
�Ko�ʪ���.�~M��U_l��7��>�aY���^ңϟ�^&�X���<27�@��N���V�׬h���f   �/Z�l��u���5���
�#������)�«�ѝ��g7�:\�):q��7m��R   �gЂ�q���z�Ͽ8.wdZF���}���gu�:E]�݇{ig�8E�z��my���jx��vֆ   N�m��c�p����Q��w��w.�[���t?�t��g��-�I��ꛫ�   �Sⴠcl�p��'�Ȗ�}r�)���I��Rg�m�I�w��=|�!����g]8   �րӂ�	�j����t��EMer��b)/	Zەl�:V�v��V�Y�I��!�   63�[;�t8	�{��$]��ds���w���$���}Sk�    �����]�Y^p<��Bj;�~~�	   l��
8��{�q��B�I���m?h&�   93<��3=?�ǡ[�M�G�nSv���p    �o�n	�y� >�ϛaԍ}���(��W'�P�Db�RS��Ҡ��[��)��e޵�����vE�0��}f   �%��-��� >B��j�S~��ly~��;�N.8�D��ұ�	f{��u`P^ܻ_fU�JӴ#�0ř0����(@   Ȓ�8	�s��j=�ٶ9r��B���3d�9�����b��&�&i�딣m/K}�a�Uc��_׃   ȂGܠ����~�v��o�S'�ٽRV��%K*�9����F����3�&}���W줟�~�   ȂGk�����0v���Ћ�H���u��-�ť��%�JG����n����Vt��Vt    C���O\�cp��O���������XC՜*�F�uWK��%3���Ϯ�tt��   @��<]�5O��+kd�٥�85,�!�1���Щ�?���`\vDe߱!ٲ�O6n�q�1�Y�f۹�t���e�M��WHY��Wl;'m�   @3p-��7�Tn��V.j*K	�c��I<�9Ӌ������X�|kK�<�B���ހ��M��vm���ˋd��o�u"z����Ȟ�Zp    s���~	���� ��;fɥ�*�$�������˫�eU��7��o9l��[�ܞ�����ʂy��W4�k+zy؞n��&���PUVVJUUՄ���g�� ��x�iA��pm5�Եu�*�v��A|��r��͹5]��^kC����2�q��r��x�#��F���>]�.��[�06    m���+���X �����?��U�}G�u���q���C�2�6,Ӫ!�iF��O	�y���3�{?9*Om���q��i����g�����5�$^$v�g   ���S��#�L�[�r?��W��ڕ�Z�;WO���dټԀ����Qن������}��Lꦮ��V�"c�T�ЊN:   �Û
xz-�$p���u��]�M�#C�<�|�<���ϙ�͕K+可���%��.����r��h��5���󑢁sĎ*�v|��   @:�[��{��{n�6jʹV���������zo=���:�$�ּ�`$��h�i�yeM���V�횈�_'ց   i������WՎj�+|���"��=Y��	�mξ���i�ǎ���z�ej����I��(Н�yX?��=������W��}��c��ۍ� �+|݂�����(u;m;�;|'}��#R^H���ZZi���:={ۛd�t���B[���o���?jc�;?ʏ�;|�qR�@X"Ѡ��9�Q��>jJ��9w��  w���0�-�����k����v"|'i%|�y�s��~b��}5ip;�E�_�gI�`��p6�v���̀�!mz���Դ����B���x�,����g�z����r�R�9����J � �݆���=����U����g3p-S������;f��|���U���"~�����Y+otG��Pw�̬r�Ű��������s�_f��yݨ�o=P�H �m�����{��Y9�]j��}b�3X$��_  
�GېiU���^�-�/lH���Vcn�j���S�wȦۖ��s��~��\���bΆ�J	r�X�5��y�N���~޷�VK{�{�	�8T#���y�]��s_g�<�w���`w�u_W�;f�9��B���_���Ǘ����44Ϊ4 @��s���9�xmE� �-���-/��Mi?�ޝ@ʃ�Av��7� ��^?4EL푅S�k��d�;�@xjg��֎��r��[��7��{�̟�\67��a��o���^)O��y���LR�ٮY��h�  P8���+-���� ^?��@��� 4���~Mݩ�M3�	�'�+$���Q�ҖI��O�� k��ɼ�ܻS4|?�f���o8��/��!��3o�ꊄ�S�}S��N���2Y9�]��d�b�N�����i�`z��#�r���z!�B4t�h~���
  �E��p�
x^�-�k�wґ�L��z�ꋝ���m��!Z&�?t�G�ͱڟW�>.E��~�e���{�����G}ED��G88�tq]���W��z鉴�WZǔ�!�Q9 �Eo�eH����^g��@uj����X�/���=��,����: @A
����xܘ�Ey� �9[�!�Rg�� �|봡�!�F����D@~�5�/��u=R_��Pz�U����57�|��Ho�u�+}!��3r���L0 `�X�b�=?L �������7ה��{+ݳcG��~�PX���ͣ��!   ��7]^���I�s5��O�"�5�����   �ˬt��6n�<6��u����ɗ���\�p��   wy�����l���^G:g��kD�Oaׁl���Z'�W��t��m*k?*��<�u �Cee�TU��¯ޗ�700  ��t�϶ ~�#���\Z��Vd��-M�®����GXy�"�ۖ�`8   ���7�!l��� �s��4�S~����/�N��/�c�:Y�c|Δ#�\���Z�ip    =>�$p������+�_s:�-�W*ny_�����[��7m���#};%Tv��I�M�oE:   ���7k�iA��}w��ހ�>����x��m�z��LznkWڷ�u+2�T���E��M\+�5E��r.�    2��
��k��<���ޔ0|�)�p����E }1 ]vbS~���Y�~rK�    H��8	�s���=.=��$��^�HJ��<�ɭ�9�W~����s��ߊ��   @�ܭ�6dy��
�ww��\�O+�v���*��\�Y����?��|�ua�7   ��8-����	>cWzui�=���V^�I��h��h?   2,/Ђ��b_��?u���T�_��&��~n��	� �;�hTҟu2�`0(���^oppP��ܗ�e�D �[�^#�K��k�W6��r���פ=�+�r�+�pm;�;|k�y��w4|��+++�
��HDzz��
 �$`p/�n:p���'ݿn���s�m�+�-G��DBW9�uͷ�o����    ��p���'�9�-iz�a9���Ċ��@|��A�2���5�I_   ��f��=��Ѫ�n�fk�R�[�m�#�3�(��
���]S��U�v
�o    K�����F F��:���k[l?w}�a�ϟZA����
��q�%�CR<`og��i+>�o    K�����!{� >�N�^����*�p� ~Xj�?�"2�#8K¡�D�J�:�C�15����aw��h��}f    �� S�1>�:�۩*�H�%ڞ�ǡ��W�z   �ȃ5���	�T��G C�
�F�Z�   ;��^m��.��1�-Ȅ ���O^U+~�����n�!��Vt?�=�i=   l�����t��k��?2M�$� �n�A�<����uݷ~�    lb����A������5|_��U   �F����]�
x� �O�PC��o��   ��\��W���^#����Bx��\?/    6�;�ؠ=o8���[���B	�:p�5�   ��\��V��=*�h;�f�[7m��+�$�<����s   �i~]N�s�,h�ݼ���'<_��=��>�   �hA�8�YzbK�h�}�6Y��.~�U���-`�7   �3kE�o�����x���W�o����T׵���z   �6t�pJ��#��@C���؊6���5xku^  ����c  �����rW�������W+��� �V�V�'�6R�   � 8õ��=��!xSkb�/�����:q�:N�5�   �B3\�q#�����{� ����Z� �l�ͦ:��������   �1+��A wQ�2^'����4�'5�������  �|�a:	�sp��f   (@���a8?� �?�����y\�{�SP؊�}\Bg�  P�
u>��߂N�    ��7�hu�nҭ����G     �3]ɼ�8-��¶ ~�_�    �I�zW�)���
8    8!����0�-�   �	E��?4;�|	���     N):[$��ѻH�}(F�    �r>������   �!���ň8{��(p���e�E1�(��aX�Ѻ#E��
  2�p��݂%�{� �0�|P��G$��~���A�[1�CV5��_�{�\�84Ev�  `��l�@�L�ν�gx� �'-��)+ۥ����3�p�� ם5��:Ϋ�=K��B  ld�����Y�?�p�'��M�����6u�~�W��˛�d|��=`�`2�_�#7��O~}��:(  �&p�5�y� �i@��#�R>���s:�K+��USdټ�Qw�3*����>y$�s���fVȇ�*� &���;0~�|�k��3��Y�'�&.�|q;�OÉv�1���͠ѐ8e ��Alqր�8w�EU)����=������z��kU�k�d�e5Ҽ�L����3V�/�u���p��N��V+�{J@���A;vPܱ���c�]�<�֚G"���<4�dX&�����>n�׹�p���������=�9����;fɪ��i]w��b����+7��h� ��;�� �;��7�z�zkU���H���<t���IE�<D�&�`�yL1�O�p��鷠<F ���XR�rY��^�]�s�Դ�w�Vÿz���;����ִs �ͬ�|� �i�;���o%vH|)��u��$.k0):��爄/6/�	P�B���/;rj��p8����[[�{�]+�7_Q;��D�ŝ��Z�5�_}~�U�N����#�ާ�
����y���F{�1�^�#ŏ���17��Bx@�x�"��QPE����Ɏ G5�H�o��]U��II8���/t���![����m^^=*�{��7�/�5���k��W��-F�2�)U�/�a�E��D/6�x�b���b�����H�O8���t���i�o��?�󻾿_���MR]��mE�qe�m[� ��^3�nIT�cmR�>�3��"�f��
��U�_��K����̴�m�����8��J��g��ԉ�]}1���c�n�k=�4��eg�� �G�������I+�G�ȯ$�!��J3�0(yHC��붟� �?�k���ή�?�����m�{M�~_ϭ4X�ik���v���J ��A�-�_���E~��z2�
x)P4_8-��� �h��v+lk�]�?�m��\C���:ٴ��
�)��U�>S��p����*��vx  |��=��a1��*��%�$Z{�9�8��A wP2p��ߞV���A}�y�{N~LC�&3�?�����x��Lt��Rց �[�cb<k��_
�?.����/�!���k�+2x�\��ng������fZپ�ږ�B�D�Pn���+X��(��[�� �뾓!:�
t.�o  ����,�C���!3�����V	��A��\|)P����y�@Z���&��,?�ݴ�d��{=�WA��7f���Z�����Y���5�9W� ���;�S`�z��ڒ%�x�V �	-6�O��T��<GZ����۬q��cX��������D\C����V��tF�~ 
�Vl#f��l8@;
̀(]m��
�+�sEln�%��x>m��n�7Ɋ��p�^��{e���a��+���g
�_�e���S���oOdu�ë�!C  �\d�����^�F�������Y��V���?BsG�=�NIz� �gA�ͭu�>�z��>�f�zٖ�q{O�:pmC׀��G�
�Z��˵�[�w����3_w�ʚ��GN	  ^2��Akp���Ĉ�O�������1�S�����=�d[����/Oli��1<��K��ȴS�5`��gg����K�`��XYqP.8�lT�[���y<���eg��\���  x"~4��Ы����o�~�Hɵx-^,F���� �?�x賛}_�Ϸo�fMO��%]���_R��\�v�9�g�������hZC��r�⊔˻
  ��.F�Cf<(�RT�>�w�/�2mI/�3Z�q;2#N ��4�s�N�%������o���^����Ԧά�O��'��Nҵ�  �*�.Q�������Z��H��������Ȩ����4���y���v�*�W<(����V�u���Yמu�V�%ٰ���eǺbYW� Ȇ�����S����s�*>c>^$��%�mG7���@ �@!��$�|����]���6�ri��y_�̪-��)a�]CwgoL��;`�vc��a �+[��.����3����.|���5`�L�)��� ~��v>��'+�^���d�ê�  ��A�ȯ����;	T�)R|� �
N5C��"�/�|*Z��|���������[�@  @��&�/F��)�� n
�/� >�����<���.�-��  �����Yp�˨�c�Ik_�@��p�V��?��ihA��t�[�|��(�M�u��N��7��?���z�&��|�؞ �Bat�!( C[������T W�k�#���4T��|m=w��֣�d � �f�ɪ�c���qy����h�\��M���s4�{1� �B`t~AP@�^��_$P���!�X��?7C��0�z�T���ϑ���g��K�'�~UYPV.�n��9���A9����W�Y5�?F��Y @f����:
�l#P-�������Y"�w�>-��� ~�S��O�:[v�\>vi��g��(���J��>h��N9���L�8,S�ⴢ �>��"�]�5�H�N���m�9�4+�a�n�q�<��#��dw������B�7�'�m;oUy�H����}R��L����Up  &f��������f��H�VQ�@��b�8�ۧ�+�c�y���f��>�#kpIT�5x�eӞ:�~�r��j��V�M�#��r���R�k�y�� 0�ȯE�LV���Hh� ��tmEڑ���lA�u�V�hWl��p��wo���E�U��5��3p��]�K��T� ��v+�a����������9�0�,x�C���	�1���k�����2�,(n�\/EC?��p�-��
~��R���L*ͯ�Y������!���S�:  W�O�A��������@�'p��<*bf|�L׀ꈖ<1�����7�^.����V�;��h��.���v���S�B3t�3wuyh�����z�wtP���v�� ���wl�`���<ц^r� ���\,2�R�752[>x�D��'&} �����֫�}K�W4�E���^��|���E։���}�յr�
)	g��5gz�u�ZZ)�X5E���%��  l���xR��b�?"�EM8!�H�,~���_^o��:�OL� �hӞ��ۦ��{�x�D�b)�]RZ�{+�ʦv���T�'����w:��th��#���j�ǟ����i� @�^5��
 F��	a�`;��k%<~<��e��#*�Ƥ�v����|�\0U|�3�JJ姶�˩6�o�1˪Z�K[�K��R_3������������� `��Qk�/pJtW�^~� ��vt-x����0����L� n�Y�����傦i��Y2��p0�
�m����ٲl��U�Ȑ!o��k{��}�q��7���%���X5��j_�˷_S'�!��G �lY�;~X��_�Ϣ���n��K��0�gZ�w&m ��jm��ա�+d^��J{t��(ν
nw�V��
�]}1Y�ZO�ay��5]G����r�%գ�����0�p @V��*�X����A�bI�lT�0Qz5���Ǥ��r_�}��\�ͨ��*�`�R�m����Ɏ �k��j;߰�G����Y�����㹭]r��F|�[v��& ���
X��ٻ8��2��ϩ����tw��	da	�-��EDP2�8�0��wT�3���2㌎3.�a��¦�a�BBHB6������Kz����s*����VU��NU}ޯס�TwWBR�z�Fi���<.F��8�\,f�43�S�܉��֦�2k��R�9U�=��qjQ�.\H���J�c�i��g��u���ʷҪ�ǯ�!� b���AF�Nti�ץ��t������C{����V���
v3�`�T��/0Mܪ7:Yʼ��s��o_M���ªI�l;w2|��YRd��%����lZ��2 ���wǂ0�;V/�C ��U������ΜF��l w�}B�q���R�.��q�~�������ޕֹ�>�$�O�%mE������ ��0{5|G��DtܿD G.�U���c~�M(���:�j]���%Ș�੶Vj/��@�/;H�~ҍ����z��'�<ؽO��#�/f�*���hE ���e�Z+@"�*8N�T�Bx�c~j�p��-8�b��l����ሂ��S���s6��g����hR��.�_2�헷u����A[�4�����%p ��̞'HXx��V�-�Iv��< '*໛B;U�<U�]���aΤ����X���xas� �������$�-@2̾�� ��i��V\�����Q?�Lr	[CsH�Y�$�s`gA�,K������Vm?�dZg�?������K��q^"0��}���c�>/@��;cO�h�0� �
>F O�qm���P� �x������;�gd��zb��{��5�ϰ�;�g���K���Z{�`x����F��o f�j+,��0�/�;��;�?%�p����zI�Qnϐ�UY�)��nٮ~�M|![����{�� �mif����7�[�X*���s� n&>>Ѻ��n
�
2�`�����ՖvIg�w�e��O�l}c�\4#�[ف\�\C�tЂ�B��)�N 'س�p8-pq�H��a?��h塖� �x���0�q7��=>�7���5R[�+ D�h�����PH��pL��H��\c����Hu���_�.Ȍ��R���P�1�ōʼΜ(p �
xs[���4��~M]7T����7�ʍ�KU�-�(l/���
PP�M"}���Yf�1�p���m� n���{q� s
6��?V,�I�6���ui /�4:r;kߚ�ү��;9_]Q╳f3r�ү�_3n�%p�;�����bN�,��&@������/ԣ�ڬ�C�!lj�d1!
Sh� ��*��a%&��a=�_a=���)J�޿ݺZ��K�v��� 7� �ۘ3a���um��~t(��jW��-��%���jeƥ+��m�b�ޞ6�CjK�����r���U^^�?A^[s� �>� �t���؈�Eo;�4rpa)� noC��:h��`]{iW���C��4�vD���j?Wkv�V߼�G�/<���ҹ�[�6�k�;2v����;��Ϝ��6O@�h�9i�O�p$�~�
��w'ق���:+�kܹ �Ql _�ք�7��@t���)���W�^s�v��Y�b�M˪����;W��O���[��Ty���'ֵ  ��H'�Б&Fp��m_̓9&�%l��Q�s�]H�R�\9�����S�BW9�U�]�vǴ�l�|Y�<��3m��:�}�Ճ޷�@O�Z� ���s�m�H�d��������]Qӓ�-�π?���D�q�r�1ӭ��.�p�1I�?�*x��<�lZ�^zFɰ+��ۦ���5:�5|�m\��~��U  �G�92�6t��Q�B�^���:<�f�Eς����?ܘ�1�BR��7�N��?�r�"�)G[��'x�dӤ���I����I�:��z�s��2�A�'O�G�8�y��e���ԝRu_��C��.  ���	v��8���OMl![�C����g�'ZW�[��zazFt �k'����ץ-���y��z�����)��q�$��=���ڥ��7�*�A�S���E�K��gZ����[�/�Wz���w�O>�3wl� ���&@�izx��� ���Y��єf��D%|������lCO���귯Ns�]i�wGdn�[�5x;�z���d|�
���)�_}��~��3]ן��uK��g��ް�{\�4t_��TΙS,�O	ު�-,_9�u 8)*"�#3L+�p��Qۈ���d[���m��o�z�r����
���j�#Up5�����N�N�L���t�V��m?_9��m�>��?���g�)!\i����uۊ	�����Ȱ_���{ʌ�P��1c ���s�@�E�3H��,��V�m[����F���[�p�Љ��GC�KG�I'm;w�򭒭~�Ϸ�2�!\�"�m��U���B�H�n�O��  0�0���8��(��%K1��oC_�=�����\b�ƜX�6P��9��m��8�KKK��|'g��R�~��a�vr}�Ev�;j����#�Dh���nul�[V�~7  �`j 2�9p�S`�L��(oL����������WV	҇ ~��Up5�l���!}�%vK�A�̻]*}��g�tp���-��}�Ȩ����Z��y��^R)��C����u���g6v�v��3 �Nf����If�M���>�_��=U�~#�S���o��W/lCO+�	騂��N��Ɂ������jRA\�w��5	x�w�����D�����\=C|�䀔y�8��)�'���j�_�i�7��r�  1�d�v]Ё�4Zq������ؕ�?n�:8z�m�iB ����"��εi��i�����׏tM`ډ�x�����\��>��~Y�ݑ�V�����=w��g[�����Z  F��cȊHC���( ]n��Z6�$� noCr}��.*ۮ�QK\t�� kޚ �}�t�[ч�-ѣ���r��:�J�cR��NE�7�N��T��q�� �V� Y9h=�-@�,;�T�[Z)��Mm,SO1z�N�B��y�!�Պ>��@�d���;U���SΜ� @ZD�QݐE Gz�ze����CZ:"���6��'�w�[\�<��#���,��?�6�!<[�
�*/� �W� ��0#�v���^�C�XːG߆^��5�X��uy���,����8�R����nt��:�z ��=֕�SD�1E�?#
HĪ˫�͝�~W����6tU��k]7\X�C�(z� �� �<�C����"�7 �p�~�l���9��-� >HcKX�X�%V8� >�|�l��� @N`�)�KjM��w��Ry�ŕ���Yp�\�'^��cpf�D C>�p�N����}a�,���3��ꛌ� @�2��#۴�K�q��V�#��Di|�dwSHY���2f�B �xX��vt����YVоlA��3�X�'���+  H�U���?�pdȔ	��l�y$�'΂������VtlV�_�m�3�{I#����p=�K+���9|�rϨ  �0�D��Ȥ�-���tʫ;���O�X�m]щ�?{|��3�L O<:3�6׎([�k�|�����*7  apd�I G��rEu�<^	�据�%�u\s^)�SD O���+��\����9ђ�O�ީV���� �8�� ��[zF��ti���ń�p�z7[bK���_ݾ�ӂ����RA O��Z�,kK��s����C�;�*w{WD��ﵮy~s�l�K� 48��
8��+�奭�r�hB5+VIl}�i�Z"G��x׻�u���I"��@��׼�T.<�����pE5\��V�su�;�*woȔ���dcC��f�ܦ �YfJ�CȐ�>�����ϿnN��oE�ë��dNп|a1[ѓD w��]mK� ����o^�&���s�;�*�>+po��#w�ȣk�:� P(��2�
8�H]/��iw�&h�V�ձ������'� qᙘ���\j5O�ʭs�M}v[�?* ����-瞖;,8��
8��+&X!�K"Q3�_noE���x�Z����lEO<bA|�='�K��Ӭ0�j ��}�
��2WBw*Un��nh��h+�Z�>{B�#W�V ��,���<�O�N�c7^	����]��b��7�V�ZoG�J����,������V(���|��@�}`�����z���Ɓ�ܫ�<��Y	W�w앝�����)��`���	o� �t\[ѷ�M��Ʒ��K㡗;�~ەEB%|����^�Va<@O�ֶ�7����==���- ���rF����apd_0�[���獉���Vtmg�*�y�3���2�q��T�ǉ ���
��c!�����`C1�<B���Ȧĺ�tY��L�|~�����d~��J��?��3�o.��>pd�ܩE2�. S'����g��l�	I�� �6�p��t ����En=ъ��I���R	���f�ß�f*�c �#+�����Z���^��u/���X7�^#p	*��68\d�Ā���I�&�+ᑨ���ȯ?7U�IT�GA GZ���c2zP�'db���t3��3J��8�@^�����MB�KPG���.�.���%[�3�cU�[;��'�����5Q�*��X%<�mo�� ��X;|a��?�D�NȼiA�
>]ަ�V�?vm�}ن]��?3�8�wb!ܠ���#ۨ�Åt+z�<���yo��w��|��:������7���1:�=p���V���AY838�t��/�/�/��Ƿ����+���̀y��p��p�#�<u��g����U��{!�S"U�_o�5��'�������}�L8�p!�#�4<��YV�lA�ݮ>z��G���+�d��2���u��@��8�'���b� �b&<�O-�s"�|p��K���N�$����W�_�ݫ����Jx|&�J����V>��<ޮ��>hoL�]]����xI�]oh��q��6̄g�����N��&�{�WN�o��)��Z	���O�����L8�p!�å�kW�h~�̙�]=V��������}���׺��ܨ�3�=f³� �l"���޵��>�luꏙ����{=T�#�#'$Ӯ>�Qg+��K\��H� 0�%� �S)ͳ�!�8�O�%�V�P8���J�G���� ��3\���K��)ERY����� Ә	�����p�3g����	�~y��ה��=>ڙ� �̄g�݆�� �*@.����%[��|����W-f�?��f�w>2��+��;W��-������
3��8��t䈀ϰ[�ﾯѩ�쯄o����ۍ��R���<J.�g�=3|8:����gU�z̀����1|��W-2�;��×�� ��XT&＠B~�J�77����^����G�f������J�c��Nȼi��!No�̽�� 
3��/@���9��+���-���q�&�+�)��z ��OL2g���N �k��V��
ܻ����]��� �0�F���z��-@��3�53�r������nrP%ܺ��n��n�5�?=X0�p8�&�V������D袵+p�r�>~T  _0��3��,*��QX��o������W­����	�u}�y�҂����1z~�5K*�������8��ĺ�Aǐ@�a&<��|1{� #�	� r�-WT;�O�����ᶈ�y_	'�#��X��N���9n ����4�����/$@�i r�%g��{.���_v|�sP%��϶���"�gn���J8i��w����`0f��D���H7� �<���/l�#�a'o��J���;}����7��.o+�pds� 06Bx�����~FY����N��!��9���T	mWo���2���伬���q����݇��g[ 0:B����b�<,@Z��f�y��˪��͝��8�a�T������A��OͻJ8���+�Tدk����������=�����ΰ�#� @��g�#ZOC �T	�쉆�����>;���̛7�p8�J��c-_�#���P��������`0B���1	�HOu�䑥g��k!�:�n]��}���M��>ů��/��g 2� ���᫻��e�&t=~l޴���?_?64�o;�c?��.��(x�����_[�x�i`��	�o�{i��a]���t}�A�p}�G��T�[kk/<#�����ih��}a�,���3�2�.0��@���ؾn��r�y�r ��s�b�Z!�|����i�o��&���U��i��4���d��}���w]_�vI�V�t�΄��l8�m�[��\Y#���H*J���Z���@�u��I��͝�eo� @!��pg�m�p8�S�1 ��Z����j��uF��e������~�E����zE�o]ɞs��pd��#�����2�.0j���@��(zݶb ��� �3��/�ͱ���1v�����X2�?9��P��+��'�.����������ȡO^W�`���sjK:�2\��E�KdΤ����J��50����G6����3 y��p.!��Q���򜶡?�j�j	g�K�[�"�y�έV�~��:������j��Ϛ�����]]�y�,_Xfyv�gv �f�Sc.��q��QRX� �\u�W�k�����H���V�&J,pG_�����6��s����L%� �����[�mW�	y�# �Bx
��aݥ�÷GH�Q�\�B����ߒ��@���_���)9S	'�#gmW��jY0+(g��y��k��4 ���<�
�����pFD"�.�]�!@�(x�V�o=���;hK����y՗���{�����hJN5p�;ޮ~Μb��W�: �Bx���cU��gH��\�B�U�߼�j�a��p��]_=��''��j|�������kW�|a� @! �'Gg�p$˿$�U(@��I���u#�p��n~����}{����ȵ�p8
��vu�b�C8'<	�:�!*�N�D1��B��g��q��p�2��p���M0�\T��J8pf�8�s�g�]L8�P�� �j޴"�h^����3_��J��~u�w�xĸ�r�U�	�  �1Bx��g����� ��C�� n����A��<�>z<j���JWU�	�  �9Bxb��ub�6�D�0��Jo� �N����G��#��o�J��^<nW�?��T�	���0 M�	0Jb!�����;��7pBe�����-��ʠJ��6v��n~��uE����7G ܄p iDO���zC��Fbh��( 1��"��R	}w��/����o'k�;*Y��� ( �npD�8�U�£Y0	7ҍ��eथg�ș3���q�A���G¡�v@�{ZV+�p  
焏�w��¥�~���� N�x�k��Jx�����������[^��J%� �	3� 2�s���(�J��6��W�3��o=��+ N�pV��RZ�E�p݆���C7|�����ES'�2^	'�n�8�b&||���V�!u�JdK`��0��`xg�e�p���	�����C�wN�?-��J8 �F�X�����y&�Q|� ��*�L��ˁ�!q��#'f­+����Y�q[m��3V	'� P���Pt�Hd�H�s��e��{j���L�1�[	����x>ӄ��%��[O|,m�  �>���FA҅|����&U��ņV���>Vq�;Zw��e�7���� ��>OU,�w������Q|� �Iծ��C+�������u���n��B���L��ᮾg  @f���@$����Bw �� �IU93��)ܳ~��vi��}|e��fI�y�9q�  ��!���(�!vh!<��b�~�
����M(ˉ���W�x[y�o��Qu�;z�s�� �귣[�s�  �E!�0eg��zPʭk�u�<��k�½_��^�X$V�	�  `X����Bx�
����s�#��`hОd]z�y��m=�O�W����j�~̱J8  ��>:=�ʌ���� �F�]֣�@A�ߒ�yo�q�w����d}�#�p8  !|tF�b��"����g��*�?[ �A[���7��A��?7U?�#)V�	�  `L���鬰y�"ᭂ�e5Vt� HMcKH�@%��3j����CO~y������+�p  0.�����`���B�A�1Jn���� u���"���G�b^����'�8��x���� ���G���̎^���v+|/ �8��<�_	�F�x�W��{���IU�	�   !���e���D����O�ҿ	\, ��'-�q�*ᡰi��}����F�g$\	'� ���G���4J��cO
\�3A��[� gmj�<�_	��3��}�1���5���� @R�3J>`��b���.�;#6�� �Z�V��"��A��Ξ���o5��k�QR4�J8  $-�+�O��(��z�5W̞ߊ���@�;�ߗ�Y�9~�7�tK�믄�wG�۾���''�eAϸ*�p  ��{�:j�$����P�ݿ�%=�<5��ͼ7�V��'u<v.T	o팚�n��G��$���3f%�   R�&��#1���X5�
�FA�Ϸ�+|{&��ij˚m]R �+�G�G��~�)���N2�JG��� �#�	���j�����P�>1�� ������J�T	on�����;���Ψ.�X	'�  ����S%F�G�GagZA�1��AA�Y��:�~�' 2��7:� �W�[�Ƨ|8����̚rﰕp8  p!|����_,f��̆;ɨ��
�EW��ymg�ll��l�T	�4l~���}�t[�QWyj%�   G'�,6�A\��ᭂ.�U��S@f��Ƃ�~�_	�s8l�}������֜T5�N   iAO�nJ�.��],��=�x�ł7΁��w8$���.nP%|WS���/�����ƘR�믄� @��|������HߋV/�m���N#p�H�
�T d���ڥ7d
l����!�?x4���1����J8  �!<A�Yb�̲��J;���V���g�K�s1� {ں"T�T	�����_�Z!�kF��   �!<	�
�[��kbA\+��R��<�"+t�� ����ǥ�-,8E���u(���_m���'�	�   #�I2"EWZ��J��:+����:���3�܆�w�N ���V����w7���Խ�   2��"�1�K��� ���%�S���5p�����vE�}�{u��<�+U�u-��N�z�   2�� �D1�׊�~�
��ba<zLr��L1'B��V ���#!��g[c�g'Y���XL   Gw��V��&+�o3�VlV<����Qn�m����f�gX������$�   ���0#(X*�,������N1�[���E"nؤ��1|b���t9iͶ.y��6A��   k�i���4������X�1��������>o�Sm]uv�a��.�u���ܧ�o$�   ���!z��^~c��4��a�5��}u�9�u�v���6J�/c�����_�61���s߯�p�I��ߎ   ��Y���;3v|� �I/o�{~D�<8  pB8 �WskXQ�8  pB8 ���~zPzB� 5p  �*�p p�/=pH����   \� ���?��78�   \� ��/�i��9��Qp  �Z�p Ȏ�y��ic��Yp  �j�p �,�w�� ��� 3��E   9� ���������fp  �3� �7z���_"��   ���9��M������#� ��C��h����C   9� ɡ�<{�   g� 1��g  �4B8 ���-��Ț6�%��   r! �G�v8  ��p 8���Np  �7� 
����   ��"�wn �g��I�5Ѱ_��?�Һ�O�����3������z�G�n2ews�m  0:B8�B����7��M{8R,���]/r�lC��Э��p��c�q��
�Mb���w��q�H{�  �!� ��x����A OQiPd�,�E�Y\{�!<]&W�%r�|�\����a��r�Ȗ}�n   �p �#5���a��ޤ�<W��P��t�!�X!��3E*J��p'o�Lú�o������U䥭�4� � ��i�C����a���F O��5x[�{bevC�h.93�=��+��V ���6Z� � ��#����u�ͼî~#?������\�ȼi����J��E�u�iyt��#kM�u  
!��;�Wwtɫ;���eskX�����=��
Cn�Ȼ�� ���Mv7��B�����G�;����O�{��A���M9�!  B8�lz}w����-��� >��3Yu�ȹs�/x��.��K"�~єpT  (�p ���=Q�o�6�匩boC�qn���X�O�S��Ă���� (�p �m�<��M����Y��W��8 ���Zf����	�3�r��D�����_2�7 ��G�������U��s�,���ְ^^�{4�5��O���g�� �!��~�J;�#*� ~�E�����}�Cf։|�1S:{ ���!|��n1O<��/�W�搷e��#�<����S>���O}�����3����??:]�=�X �,6�O`$�5pk�� ��]��
ᵱ��~  ���m� R�����I���&�|�Z��к��u�!�yԔ?n�%   ɟ�v	0���f�|i�!�j�ɨ,������p   `�)���qF�����D�{�G�:�����  ��6�ꖾ0��1���������m�iz����|�<�a��gE��a늜x=2��h�{~��\�~�_.   @����?V���m ���������h@"fP"Ѡ�Ǿ�M�
��^��qÊ�O�x=�֥�ɳ�/_`��!�?"�   ��'"�X�2�_wA�·�w�
�E��b+P;����<-�/�A�c��V�3i�i�|y�ȗ$�@>{����xvPj�}2��'E�L���C{WD�:c@[�r�xXv곏�ڲ�3-�*�����!��7f6|�B�V��D�ԙ��VЗ"	Y�u<F߉�xg�Zկ:ǐC�"?x�`d~v�̨8r[�!S�[C�b��GC�qw�<��M�t����w֊�;�'���'�_�Ε5rΜb�7-(E����VQ�/5����-,M}����� ��z	�[^�ٓD��2��%)�����T���$-���#����W
���iB8���0��nF����bY��B>vm�]a}b�q��U$笙A���j�h^iB�{��j���3J� ���7�4(r���e�������v��mt�[(Rq2�{�,���x�?!@6h�u��2�Zm���i��9�� rۏ�xT�}� pF���u�!gNO��2k�[+�n�K�B�J�{-���}�δ~=��m"��B�=�Ϝ��X���M��5|��� @z�E �������o]�>QU�5Q+�G� ^b��+�w��k���"����n �ms���u�������vp  �99�߶ؐ��*}�[��Jrt���r�~�}�j�{�vO�	��9#@�i+�����s�Ch��WMJh1ގ��r�XH6��}GB#ާ�1���#fe��L��Q] `���s��|���~$R"}V���f�t��p=���mO����,y`5!��.�̎q��s���N��G:
+NC���S�p ���Jŋ�2w������(٢���n�2�}�t�����퇚�}��uh(�rq�̟^D ���E~+|�˰���`/2��I>ҟ+�K��XZ6��y�!�����n ��b����t~��eU��I��]7LL(D��oޏ�mO�I�8��`�Ǜ]�(?�m `<r6��q�!��IO��ל8�;E�"�M���Y#��m{�"��͐O�WnV����.��J�CKQH�y��x���3�>�l$W�SV�|<�[�X������ӷ�㇏�/  
UN��N�����zB�주
EOh�|-�/g;�tCV-y����Ô�5�uڄ;�g��6yv� ϝ7�E���+��C(ꑞ�Wʾ�b��Z*�hn��|����pm{��k!�O\W;f���#�YZ @��d ��i
�}����B[��q���^i�K�L�{X\��ʥ���E3
��92�$���>q���N�ϾȆ�*y�@������>vD����#��3���G��VM�C��-,w�����  d@���_j�ҹ������q���c���q.T���v�!_��{��~oT��:"N?&@!;gJ�TC����ז{GSix|��NY��b؏O���,�u��2Y��|ď�wE�  dPN��Z�v�vÑR�D�R�zõ�È:v�+�h\�O����'|'̮���/��N̽v��6��ǳ�;}��{�p����8J�  �r�ɪe�o=�������pg��r�pq���gp '�Y�.�%�zc��=nL+�u�[�G;���Ϸ0� @��L ��VS�5�v�9N2M�}�|�U��O7�sD���*x]i��^����@!8���"�j�$��]��bď�8�+l#  �r&��<ϰ��v�iz$�����
(�׹����4���Ժd	�6S+���($�97�ƪ~���7  dCN���~;{��H�]���V �aǎ'��úLY�]\C�8U�/b��ﮎ$fق�?����n�  ��\��+�k?GJX�6�H�������<�rA$G��X5���p�P�538�c�X�*   ;r#�;\��DKc������W�cȃ/��u� ���ȭ�6~7���P\�d��o��  d���%�EN��d������>o���3գ�+�N%
@�\�p�'W7�Q[s��<����p�  ������N�A������[����_�P�GO��� ���̑�~�3�E�đ���  d���n=��L�nO��z��OZ�<]"F��i5�\i��?n�
�9_�Д�+��k���~hn˖�T� �&W�Q�~;�|��P�N�>ia�p�3`�X�\ �w�0Q�/,��}�M
ŹsF^�v��p�� p+Wp��vJ8ZbI� 9���.1�ԏ�Z���9�L��$ ��7^R9��Wo�G�N _0k�>Z:"  �˵��H���1���T���l���+V �@rt���WM��S�F��}����?k�l�C�9  ��� ~���g��#f�oD�E��E� ��+�t+p/�����;���k��3)   ��\���~�������H��qq�H�/��H"P�^������Ɔn��=���;�_�  d�k�4�hΈF��k���"�!g�6e�v G�wE���䇏��P6� �f��>����;S�F��;H���J�\�3۰8s� R����7;�m��  �̕|�L�s(3GL�ϝ��7�֕zp>�^  )�!S�����x ���� �T�[i�4�����M�vΞ���T�$N�Xԛ�R���P�53H�   Y�� ^?ə�����8+-v$��)�"�- 	[\_,��ϷP�s�� �2W��������B�W��֘L 
ڥ��1���رų�����X9�?WZ	�m�)z��5  ���3�Or��4]���<S<���##���)Ն���0]�f_�Ε5r�e����C�xI�t�D
����Of���ɜ @��.��v��\����t��֐pʷ�-� 0��o�6e�j�t�	縭�Ք��|  
���5�=ѹl?�>��Áߪ�p ���w��(���T�(9��w���ښ�������e�~�~p  ��}��
8<m�6tP�����Q���uö�k��VM��>�$�h���?��lB  {��}<��v/�p,$�TN=�QU* ����l+�T�����/�d�ԟ��+2l���ƺ϶� Ȋ�߅�ȡ9��͙'7� ���3��.���go�(�o{�54��G�gq=��  �-���m�����p'T�h)[�$�{8*_���a[��N-�[����-�s7��1���r��2aQ  ���t�*�Q� K+�:<V���'�w $DC���:G\:v���Lt��\���юl���Up  ���-�̀�s��1��_mC'�H��ϴȹs���y��i�����l;�3Jz1Up  � �+���SԱ[��9�# 	����/��m+&�q��b������*���  Ȇ�g���fC����=} IӖ�+���Mb�ԟwc�ȳ��~\  ���t����2���v
 �D�}�CS����ͻn�(�~�Y
�XUp=�m���X7  �~�nlA�&��'x@���ںFZ���*�u���Mۻd�%#~Χ���_� H�^�j���`��v] �	9w[�9�,MgxG�sc 
�h�t#�'����ݳ_
ɏ�<*��2�r���~�^^�)�#�  Ȁ����u���������S�ea0�:Z:9�3���Ԇ���a?��؅v6��'?y��G:�L���w�ʂY��o�ׅx�_5A����
  B+�M%�F�׍p'��D�]Z8Ղ��7 '��ҹ�#.d�iY�Z�W��O�Z4�qھ��gg�ck���4x_��|�  �݌�X�v] ?���́���Pz3c� �߫[�s7M�cڊ��M)������
��ąVï[Z!ϼ�ao�Oŝ+k����2wj�  P��
��Z�>����a�=}�)74��b�<����gaq�����
Q 2@+�W..q��E�J�l��p�A\�V���j�v�Gv����Z���2e�OfMȜI��  (0����k��V��Z�l?螃��8xJ��(�m����8w�j p�.;{v�s���s��4�w�D�`=�L�@�9:;?�L��   !Zהk�����M���vG�M��p�
n��1�$j�,���|b�P�{�/ �]>��W�G��juVۣSm��E�37ˇ��0�vt  ��z�MV]V�n��Xܙ��jm4B w��~{<�=as�t i2�B��\T)�o�,����M_/��ז��TÝ���[  (Do��~+����m�E����mi EJ�����&Z���n��mZ���5���B���Κ�[��N{����խ�� (lS'�,z�f����ɺ���kJ����bgnK��2���'r�����mj1� H]�lAi��P��M��i5�Pi@<�_��º���m-�q��
�=�ĺ���4  @�:�t�Ʀs�c]u���rn�����Sg��p����]��^g�T���G��c����׼�3;$�h@�o��Z�
Ju�W�K�Ri]�50ToȔ��ة#�-a9z<,���y�  �dP �y��)վ&�M�J�)ҳ�w6�r�gB��蕰�R����܃��Y��<)��7�64���� ��k�m�^��㵣���~�Yk7Y�S� ��mi�m�s��1�~Wv7��t��+ ���9 p�����   �f��m]�f����]� �x�좦��vM\m�+r�����vJ_� �,}���r���0�1��߻ZJe	d���E(B   H�y�R�:����cH���E�*��Ϟ]���+�E6�uv�����D�QW��9���6�W�z�\�Wtˤ2�J��ۏ�   �6|�e���Y��]�3��TY��m�tn�7U:�қ�\r�s!���>x´�\��p�of��<n_[����F.�?,5%T�Q��"Y�X%͝�=	  �"�~��"=ul��:gv����l�JՋ[�
���^,H�H$��>qᤍ�����ƶ#�5Y4�UΨ�|Z��ǋ嵃U���R   �0���nπ[\Ok�R��Ϯ/j����i�)�!C�\V��t�k�wv=�3o���8Z&;��ɼ��2��K&��I����q��'@&5ueױR�z��~   I1d�uoI��l�l�I�G��Μp�y�چ���W,r�L��2�H�D06�g�;{Lyv�;�χ2��L�^�i��?�4�\7;�߃����W�C���1   �-�Y$>\ή?Y�ϝh���6i��j�Ko����M���<]��s'=�)��
PȺ�|�˜5  @>�?�{�̀=�������w�mϼ��QSN�6����2��FH��V	E�6�D�#��]����~   ����^8�����W������&+�����%��z�U�9{�>�>��B8�����M�٭���6���    ��|B�w���q�3�ֵ��ם������s�8���DM/��C���N{r�    @�[0+0��V��Ϝh�Y�k�{8<U\�}����h��;��V�	�i��H����:?�p�)\O�9   ��;��~���qC�<:�����{�qWmCW���U���'I��zzş��o�c���   �M�|��+t�w�� ޽���F+��yச�M���,�w>�F���Z)Tz|G%B��    ������Ȑ��p9cj@.8=(�����ݫb��ܶ�<���r)�!Q	���v���5e�a   �|տ�����G���+��N�5vJܺ��U�dpWU���_5�y"W,JO+�.e3��􅫥Px==�K��8j�ϟ��    �ٳ��e�Ƌ����ΞSO�:eܺ�[��ާ�V�u9{������)�����n	�C��S<����1��3�_��ϊI�X9    ����48r���]Y�i�Bx��_�t�6t�ѵ��WW��
��
�Cx�H>Ҫ�V��i�fS{��7   ��gW�/�v�y�o����Э �m���Ϙr�<�3��U������J��!��Z�餋���	    
��鵾��Ǎ��/8=�x��@���}��GcU��-�\�}mbD��TJ�ӊ���*������ys�    @>���x���q��>�쬠X\���-"?x�^���sҺ%=)�H�Dr�V���N������{a�)?~��7   ��7`�y���=��x���#V�E���Y�p�������U��J��3�D�]���!6�k�h�K��2+���t��g��.Z��Ք{'|   (�����F+xw���#΀[���u��k�+�'^��r�,���cV�Y8+�!\i%<�9fp��F]����0"�wf��=�g~   ((W�3�N��*�z�^s^�,+��K,ٻNgO,��vC*3����zE��vk����oO��F提{`�)O�N�   @����Y�k���Q��������3���E%����N�.��Σ�|iUf����zE�+�Y��(�a\C����>!`�#;�Oo��=Z��:K    �Z|�{���JW|�&e�y�Xܞ�漒+�7�Kg��7�2���2��m8ښ�>�y��i�� �����-#d}�^+p��_7�4|���o'xg�(^�Q    ��=�=�ʫ��c�y�Xܞ_rZ���yA���΂+]ʦ!��������gް��v��x��[���$�r�ۑ�]�/�ط�m���[ll |p��f�%2wj@�K�2��/E���>�LinI���౐���K]Ӗ���Ε5r�e���t�gv���̟�)�>��������M{{�M���!�p��r���{�Qw�k��+"M�a�ߖ��C� ���δ�bϸ?<��ॳ� ^/.���ׇM�)�|AvC�If�M}�q�S�)+d�w���ǫ�Ք�����#���/s�5��:#ҢWGD6���m�Lz������rY\_<��j����S�d��2�h~�|�g�z;)���go�h�t~�[����敞��@�_��K*���-�Xݚ� ��7X^5(t�O���U���/��?���L���x�;�'���G  �����3���8��ӥg˹s�d�.W�o�?�ܔ��Cd�in	�ËW�s�{���`�x��q�OJ���Y+;�f���owL��gdp#g��a��낊QC���j҈!w4��żiA��#��П��K*����������t@  p����k�-]]W���w�x��Y��+�7��g����G�|y��U�;�碶NS��?�o ��xU��q��~�)2�r��+g��O���g�Vk������=\[�����cϠ8�G
��s���N��̺�)ߏ>���MIkWB��� Pp��o�߫��	�~Ǎ���=���%}���-��\=��M9�*��+�N�{ؔ���@r4�j[:�X��`�l�����jK�p�[C��ݲ�`�)aRC��s�e�䀜>���p���Z?�g�f-x��'ֵ�x_�<�M˪��?|�G�����@:{���[�m/�ªI�bq�� ��ھ�����������cG P���-�k�?�
x�,������q?xPX����S�F�)e�(X�7u�Y�԰5��/f��H�Vۣ���iu���Я����<:���ҁ�4>7��M��Y\�g��-�-�Z�}l�q�������O��=k ן%�n��_[3��ժ������O|��&ٸ�G>w��A����d��85���gg
�/o�t�	$ @N���+��︄#��KJe��nY�3w����ӱ�HO�[L��}�o ���+��|��k�Z���Ҁ�L��0�D��hs�k�w���=�ls:}��	��o���~Rd`X�'R����������1����-��������ez���s�nl� �U������W�>ş��w\�ܞ_����
����q��b}�Ȅr�x"Xm��'|H\�ʬ-�w���i�V睍�IU5��{�=cG��Ws[X~�B��{v#�����=~RUj3�W�[>�mݲ>����m�_��4+\;#�= ���.��_7��Y�۾��]���w\���ڳ���)�{��e��?w��,x�c���io,���2�jn5��E�~�� 5�t��p˸��YN2EmuJþ[h�~~sgΜi��`ߠ ��캎#m��#��⛝��ມ=������A����r ($]֥�{�Ċ��ŞP�7�L\�⛗�O�����ƖH���@�����1e�,��jC��[H�j�r~���=, ��xp�uɖ6'Ο��\����>y�
�٨֦��%����|a頷�ɈD��48�k�D��Ї�8��� ��bo=�����*�s����~�%�[�)�v�|YE�wmy�z[��k]�?�3˴�z�^Sn�!�N5<��O俟3����i[Rv͒rGx����.�:O�,�,?Л�bD�<hp��}���tZ�֍��mn �5ͺ�>�4ݼ�|��*�I?`I6�۳��:����[���l���=Sr��E>�_��Z&��+�*����z��;�+ ��}�|�CS�O�sB�u�IՃٚ[�����|m��:���9��	�@p��i��u�x  ��[ϭ�(;��s��n9M��d�n���o�|Yy��;%��@Nz�S^�f�mW�rI�U�7���-��&�� 2C+���k�q�g=k�����t�<9s����l��q��G��ߕ\�^K���zw&�^��ǧ��
 
J|���9���W-����z>T����\<���}�������Ӭ�=�#[ч�Y��J�����r]���A�H�)�z1�r%{Ȱ�p�GO%�5}����Lkk��W��]r�3��г��V�dg�>ɒ�b�D\4op[�����Y�>�h�yYy�$��|���9�}�e�}��m�?�oEϹ ����u�\�Ժ.�� ���ѵ"��5�� �B��={ZM�<_��yJ\��i������8q�zfy�3�C�Sie�>Y��e{����7O� @a�rQ��mq�8%� noE�,�߲�b�?��X���nEק�sb+�H4�>�6��8���h��`�:��b=��/�t;J��ϑ��i�ux�.���������-O^�����Y;�}�/ �|��s�� PP���e�����\+�]N�x�<.t��%o5�����V��%����d`_�P��3r/�o�o�K[	� ܧ�/:��U�=o{�}��ۦ�µ]Y��uK+�Z�X�X���{S��m�;��7�Z���l�)�-a�C7�k�<�o ((���w\]�z�d�#��qNp{+�_�����C}���z5xϐ<�'�r�|C.�/r�l����M����V��� n���u'���k���!���&Y�w�l}_!�h�)��#�6k=�ډc��v2ty���.[0x�[G  A祴�I[�޺��W�S�84��T �g	�{1���ʪ��w���+��[�G��)nX-2�iqC�Y\��G�ll0e�>��;LY�] ���n�N���U��c�N]�5���� ����(�|8w<UZ�Ր����N���E�# ���m滬k�9�����*͸�.1�x|+z�ܩ�+�����-S%���������n�kEܔsfrv}f������[z�y,x�q$ �AR�o�j�)��q�~=�|��5`�s����
����/s�����Bm��'fң�
�� �x�[��~��س�����=���L�+Ywٖe��`
�n.	6�BH$!xS�f6٤�tIHҝ�4�d��k�lg�N��v�v���v2�K�l�M��FHS`��`����e[���>�ΑL�-Y����F� c$3�s���q.K/ݟ���� .�ykǶ�����ơ����F���ƭ��3�y^A*q�Q�ԅ}L�g����蟯o0H�~"�^�v���}<�>K�  ������l��F���G���8x�z�=����g邏�R�[4�\�z{�,�0���(�Ϥ��m�l����  @����%�{םwU��A|�Lc�<���ǇM|�%�@��f�&vE����|�&:d;H���0.�oh,ps���~  �����C�'nry\/��[��,�y"|im��/k�9t޺�N���q�M�x]}���?�E�o,��ŋ2  �h��h�Q���v���x+���q� .���][m�����?��]��gplP d����O��G9�?�����8aS�g���3h�ky� So��k�yS;^W�	�ϱ*�u���  HM��{i����5߲DpiW�E�L�]w��_y���t�'o��qM8  D���*��U��<�'��m�9S�9��.�3����|�|!��~,֋��r�W���v�wO�0��^��'��=  �!"�o�I�޵%�%~$���%*��iӼ���v��kÆ��c/�4�`�&  �i�j�Vyq_�<��wD��ޑO�:���v�|�b�>���oc�<����Kbqom�[�x�^�B��c�]c6_SK���  �C�|��N��a�lSB�oY���+:_����z�G�����e4�  @�U�-�w��L���!��槟=1K�~r+?��W+>8�Gߖ�����rK�i�Uٞ�{� ���7_�S����ۏj  �E4�|����]���|��e�&����u��Q�����	 �pz�Y�%�u��?\��7��D��`C�"�3�)>�׆w__O>�.�7bN����{���7�*���L"y�� �E4���9n_n���[�� �h��3���t�m�	 �`mrF��=y!9+o��_O�T�bg��X��E�hK	x���L/�Q�U9�1D�T]����%L=��ūӳDR��Dm��z�ӵu�}ښoY��,Ԅ���"݃/��zFЄ d ^�ގ2�V��)�ܪ�p��p��$�_d�y�mR��Hـ7_�_ �6�����|-9׎�&u�$vsL�i���gi��~�{Vۧ���M�;�P��'�ϟ,
~�G���GM8 @���������ϫ��ï�Z�`�XK�"�NfZ?���!���~Φs�tï)dpHcr��Na���_�q��fO{�-��K�R��}�=]�{�����	 � ��������3�4�Tr�;s�pn��9�dv��%����Ǻ�ۭK#w'�'�E�V0����x���'���l������w �Hn�]�ýu����͎�4߲��&���`����O��
��A �a|��76D����̿\�d�P��$�ݓ�k]7-S��Ɇ^n��Y�z��������E� ��x/œz#�x�/עN�"�g�S|X�(Z��oq=[�LZ�-K�"7�	_Pf��D�����& @�8xs���6���U۔>���f���Sjп�}F�c��)�~9�畏_S�V�����K�  ]IDATyC��Jk�۪s�7�t�P�G�l	�' �3%x/�!޽����i�+����%��"���*K�K�Hj�-KV 5�U�&˾gK���M8 @�{p����Fijoe�)b���������)O�uڳ�#Ķ��J�WǺ>�'Y��,��Mop�����ƴ���(�m�5��:M%��=��Z�����K�/�{���H�Q_��	����=ՖB���A��|%��}~�Oo�}�	@Em�7W���3�"%���%{�W�	����{�R��=Wm�a4�  )��4ʟ���mh'­-�]]��A�I��?��en>9|���h��!??x��N^��s�׽01�,�ŜC�T���O�*�=o��!��>�F^^�G©�7�;���(w?��u���|5@���B{��M�,�������$�4�|��n���y)�|˒�CMx�Eo���*
��z��1�M8 ��p�k++��h˭�s;c����I��ZP�����Qv���4���W���k��*+0*fp��yc���yƨ���[]oEyʷ@���2�\�S��������eX�%�݃��#�8?H i"j���Ws܏nv�L�-Kv �IM�!K���#3u?~�c|�X?�p �4�A���T�D����=q=�*�L��q���w�Vq�6_0�h���	����ܴ��^O�Al�x:~}n_�C_ߐGK�a�C�r~���!E4�Oޕ�pߚ�j�e��CM��g�<�)���>4�  i�C�o�<�#t�j�N��M���X�u���/�+�ǂ��C��K�εr�ԫ�����h�������}	Y����7�"m��f��K_+�u��R�ʹ��a��{��W��{���(���a�C/���	R�p�j�K���S)�S �LD�m1�\���toZfK��[�*\&5�b���;��h�w�M8 @������x��<e�7�Sl��;;�7���*7�~񆓏��������_s"??����h�Zg^����y�7?��~��q�����#[*nç��p>a�FwJ��D����sHD� 0�w����a�\sJ6߲T��M��[w8(Ϯ�b�����X�y�k  �J������Z�m   I�|���zr[�{N�1e�oY�pY�	߹6��JM#"�{[���c+      )��5���[�����ͷ,U��	��4���3Ͻ�����C}6�� �}�k�     �M�|����'�湶��s��ͷ,U�Ln-F�᩻�:�JM���s���p��)�X     �m�滪��zb[����� �E�-K� .7��;V�LUe�v����'k�     ��ww�qY�3"����aӧU�-K� ��O�ъ��������������{x��     О^1N�q�[w8�ؐsA|�vͷ,����C���\oU��ܿ���u��6      �ɍ������|Ñ���,�r��4l�e��e���5�-�e�ν��ރ�s�A)x����pp     ���!�31Z��}�d�ݿ6��LG�i+b���ͷ,]�bm�դ}�v����Ҿ�����g|��\n"      H5�ƛw9?�n����uٴ���Mw�����դ�����|�!��7���E�t���k�      R���Wbl�]΁�ն��_�ⵛ4B+\�6|GM��v�Ž�`��w���������     H���w�U/5�;��\3t�x��i%��BkË��3�:�j�[xmxI�E~�i6�     HE�-��}����M�gH�T蚤� �>7<�n��XSe)��Q/�s����4�      �#j�-F�څ��&����,��]Úl�մ�դ���,���M�TW��.B8�}��D����h�     '��޴�v`�*[Ӫ�X�����o����r����B�6�����w�f�s�_j��^�     �����NGM[W�i�J��%��cn_F4�jZ�jR#n6��;j�I������@ɩfi�:q     ���#��h�;��}�*����Rl䇤�>�~g�L��F\ٲ�n����8�/���C#     pcԍw�G����R��~mV�������[-���Ԉ�a޸�Fb�>㣏O�|�8H����4ֈ�      �)�%妎���6-������I}���x��#��*�Q���6�r/A�{��E�&�8     du�-߿437�^��f1hy��#k��i&���\-Ԉ;��h��l��}~ih�����"��_�=�8     dE�-x�.�r�vmXl�ZM:E0o�A\I݈K��.��y�vG>OM���� �q     В	�n1����/��ޞ�B�?�������^G�[�XI[�g��c���[��7���[ь    @�S4�F�γ��\�x��%���yE0�s����7��Dm���~Q^��|%@'���-C^1��<R W7�h�     Dk��ŸT]i>�b��Yn�c3�O��4�q� >I�N驓�q1L�Fö}5���/]�����b�wxG��W�XC�      �j��i�\�g�\�%�MgE������\���#��ڌ˶����!5������h���v;[����9��r     ����=ԍ6m��t4{��f�0J�bxg����Qǿ�Cw��Mw!�'HY��!w���(7ۖ��ߥ�`=$j���t���)B:�{F*|��������%�cm     |�"��Eh�I�/Bv���9Ǫ��a���m��]��+y���lf=A� �'�urYE��B��w���g��%��a|h����(�9    ��:2�a�d���0R�-ƅ�����h�S��K��.��w    IEND�B`�PK
     t$v[��e�/2  /2  /   images/0956fa89-558f-410d-92be-91de6d3dc59e.png�PNG

   IHDR   d   V   9P3�   	pHYs  �  ����e  
�iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 9.1-c002 79.b7c64ccf9, 2024/07/16-12:39:04        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmlns:stRef="http://ns.adobe.com/xap/1.0/sType/ResourceRef#" xmlns:tiff="http://ns.adobe.com/tiff/1.0/" xmlns:exif="http://ns.adobe.com/exif/1.0/" xmp:CreatorTool="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" xmp:CreateDate="2024-09-25T10:15:37-04:00" xmp:ModifyDate="2024-09-25T10:18:25-04:00" xmp:MetadataDate="2024-09-25T10:18:25-04:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e0fa026c-2b50-4255-8fae-7a1c4254e60a" xmpMM:DocumentID="adobe:docid:photoshop:cdda18bb-8c9a-7446-b932-ddbadfa4c834" xmpMM:OriginalDocumentID="xmp.did:8deed1a6-5431-4e06-9973-719a94ef57a4" tiff:Orientation="1" tiff:XResolution="1920000/10000" tiff:YResolution="1920000/10000" tiff:ResolutionUnit="2" exif:ColorSpace="65535" exif:PixelXDimension="992" exif:PixelYDimension="855"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8deed1a6-5431-4e06-9973-719a94ef57a4" stEvt:when="2024-09-25T10:15:37-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:196253a3-2d41-47d0-8e52-c694c2a25be9" stEvt:when="2024-09-25T10:18:24-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:dec66016-6d56-4a37-be9f-5a128ae8d7c3" stEvt:when="2024-09-25T10:18:25-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> <rdf:li stEvt:action="converted" stEvt:parameters="from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="derived" stEvt:parameters="converted from document/vnd.adobe.cpsd+dcx to image/png"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e0fa026c-2b50-4255-8fae-7a1c4254e60a" stEvt:when="2024-09-25T10:18:25-04:00" stEvt:softwareAgent="Adobe Photoshop Web (2024.19.0.0 2f12568b568) (Google Chrome)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> <xmpMM:DerivedFrom stRef:instanceID="xmp.iid:dec66016-6d56-4a37-be9f-5a128ae8d7c3" stRef:documentID="xmp.did:8deed1a6-5431-4e06-9973-719a94ef57a4" stRef:originalDocumentID="xmp.did:8deed1a6-5431-4e06-9973-719a94ef57a4"/> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>}}�.  &�IDATx��}	�TՕ���z����Ⱦ�*(����DM$�cT�Q'�h�Y��b�f�H�1�=j��"(�,�44�4���Uu���w�yU�T7U͚���QT׫���w����ާ!J;*����5�q��ƃEsӲVn�^�ׄucf0d��T�%M���MSZ�;m��0~��[����Kǧ�><�8��)m��k*0�̟��C���?����Ƨ�o���8=��J?3���/���h"�|!����F(r��m[�����G�o|o��4\�z�}�N\q�8h[w�Ɯ{kq�x'f�v�O�z�3���������;�]E�?B�@9m��Pg-��\��4��pĸ��+r��I�?|�?9��g[��r�[k��1L��e��Q����}#ͩ���Bg��w˻z@:����ϴ��n>���S����ZL����ƏG����5������
�z���_���y���c`�B� tb�>��q�ƕ8����r�@�9&O}g"?�*;a�N��
�Y���

2��U�>�|AP?̶���I���x�����3+�(��qg�W�,���8�@�g�ކ ���&挬4+~q�h�[�`j6>��՚'��`�z���g���9��� P�< �a�j�Acf����qy�/�v��n<?}Ȳ��{�\�Y5��|�k����С��;U���
0o���k�c\i��9J6������D�:����\:����]t�J}c=��R/�Eǃ/+x�S_]>��]�3n�Ff�W�acx2}��oǴ�N�����u]�n�t�S_�s�X�
#j�4�Q���s�zڍ,v!7ӊ��~�P�>��u��6Y,�~�	���D L2����y��p���/��]o����+t�s��k�9Z��X���ʃ^��8oR*�BSGH,��M4�0kl~{��C����!����ˡ��#;�
�q�-���0,4�܆��3�p�=�D|���w��m=R�EUQ6DL����d��q��醝�}2\���y
~��=a`%~�F749Yӈ9dd����B�^/vD�8�f���>i¥3sq	�b4g|����J\����C��2R��dVnn���ظ�K�g�X�MH���q4"'O^�Ԏ��gk�xn:���⏇A�s����a�It�L�&�Y��hxDt����r��T�_�?6t�d[��Ʃ ż<��n����|�N�?�[@�:�4ͷU{0yD�p��y}��|\v�F����� Ye�q�P�0Nb)S�c�n�rP1,Hw��I*����3��3��~{����rӂ��@��NS���t��f�0No��������m��8�����	������<�������wu
h쟨<��X5�P0:'��\�@��Sb������`XŘB7�lf��ȱ-����w�`�t��N�C{eCl��>���T��Dז�nCs'e�����u��3Y�+~x�H�t����MX��~x�9/9��Ė+�PD!㧁N�B\�I&���M��y�0��a�^<s�g��8��X0�
�J:��f���I�J!gЏ�l6��S:a�|&���~m�(k�m�� +U�o_���sPQۍ;~�m]!B0�����~`W�BNr�f��@I�~�H��]ĩ:��B֘=�S|@HT�xN�r=��p!����)toCA��c�>��R:.&.���,�ZB���R/=L��\�o��	�=
��7������Dw��u�-B�9���>��Y!k��+"4�SH�X����[�dX�cW��Ǻ ٗ��:bbI��T���tRX��/2��<㋺�X�mv{��u 0�(`�c!�@U�~�1g��>�7�ܷT���0�,n�Dpߓ����ONa��k?Q1-��+�������V������ҽZDkj� 1�<��Ӌ� �� �z�r,J'\��:��H0��ޝNQ��,�xЇgu�0͏ݭ�h�����<7�gvc{S:t��iE�s��`&Z��0gh\�6�e����fki�C���dƾ���6��b?�>)��dy�(tI�-V�hx��D����U0��k���v+>^^��r�����U꯭/����04e�C�d�f�6�e�����,まpdF�x��*��,$Ѧ����&�h���;R�B�>x3
R���,8�ρ,gF4�w��5�CS��0��z����#�K�"��S�\���ɍ�p�9�Ѹ҉%������e��t1�-]��%>r/q�f��;��M�w.݅��w��g�-��o)�ᎁH�J�w�>��s3��&�Ϝ"��;�a�ҏ~-��u���˳�w�����;���&|^�O��2�A���!o�PL�}��09��)�R�³��+F`3��<Lk�PQ�&�z0��D�*���Sǭ��J��9�ZW���.L�����c��9u �~�_�9eOc*vԥ�1�D8�t"�$�*��G�!�a�+jy���@^�Ev<�͡q'&�U>��������6<!��l�7f'�;�2�QgO�u@I���r-���$f4˩��'c$��[�%�6P���Ɖ�E#�2��#抡y6L�ā�6��aݮn������sI���1�:��R���OrO����!���L]�7O<�}�)"�"�
M#O����a�A!A�Z阕��P���e�P;>�G�١�ViG��΃�Z �Ȗ�IH$h����G���ǥHXfѼL�o�woƻ�E3-L�b�0v�c7��i'��(��<�O��4{G�f���0�����FS�],��Hu�lY�R¨j#'�)⺭F����.А� �F��aԒ)2���0�EZ�*��T���(�C`90(11��mF�M>�lb��@�ym���qC!��:>��-b�pJu�Oh��6W�p��T|^�GU#-x��U�H���2�2(���l���5�n�~<L�b!G�2����ױ��S���c�dM�ڡH�c�tl�禗m�cY�c�bvܢD���`�L!�&;҈m�����h`�, b��{��zao���A�~��,���>�{�-��}MSن�/�!'MØb;�50���P�j	9~!1O��H��z�g�J���,����	�0k�T��~PmQ�&��y�Y�>rk���Ԑ��;i�v��W����q5�0KG���'�h�A����a��=$�6༷͟䞳 "�ެ1.A�e�:�S�Z<�y22�LV��:/���Ӊ#������m����譚"N��b��e��ӎ+���㰩����u�!jJs��m�5�B�YلZUCPR�����7��R*G��}���$��G�}Mo�%�!'�b`<z[J��Ì���!@��G��x���k�:��Wҁ��)l{����1Lꢩ�@���>TU��&���b�&d�~^����~��Y1���ϋ�?-ư/�8
S��z<�r�$���=m�ct���y�����9��7[kp� E���%���![@�;x�}eE�Y���&1�2��;j�xq>�,_�x�)�cas.\�G\�i�~�t�n���:$$�YU6�4����R��簅���{�(�����8���Xzt0z�t���ȑ�K<�M�����m�I�,$�@`L��Ol��3�]�[9�`�y���o�� ��VFV��lّ�v�HL���4.;ycK����br¬GɅ�����\�%q2$�:m��S��-ů_kFuS��4׺����{�L��#���0rd����(VQ���䡝��v �m�����2�p��Q.��� �Ab�d$���8������v�ؔ���c�&A�kB[I�\�^��q��O���]�Y�!���W���VӀ9�E��_؁��kw;���?�*EmK�LKú]^�8q�O���\�r�:*Uf97W�@�-�D瓷�pL/9@8���'��"=E�yuSxի�+�=�����̠ס���`�}F+�v3�F�;�I�j�k#���[Q���{�Ȗ� ���׷�Nj
��$�������	�>Iҹ��t�Mɲ*�?���dVJX։�rV�3��7�hV-�t
� b)�.�����Կ����G`�P+����,X[��w����OdF+d��ϑ��%�'IqŖ]�C�!.�+[�v��m��4�}e����p(c�)CwBW2�Bb7�A��@~���Km�`�^�OJ5����k҇t�BR3��V�p�C���!4�i�o%L,*�H@�2����)é�wK;�g�{V?e@*v7��	�p�5���x�����FuK.����RD�g�X��'R�q��n�a�,:�$���� H������gx����,���<��~���[u��5�p��z┕p�Kc��
�O�.1�UۻE��t�%�b�'���� *���$�=fD�!\4EgX�\�1��:G�_B�6�O�%$�-%d&͍�P��(�����+��}�󻯛2�Y�!^ِ�[��IV�NL,�#�lSUy�㰹&�1W��0*j��{0(�@��3N+[���� 7%�=��R�� �چ�h�}��q6�kA�-����lIC�=$�8���.��t��I�B�����Xh�N�?jE����*ᗙ���⊬��^��r܏܆�ć "��K8=i�2}�e��%�Q�����A�!�6��aT�8Ǌ�fg��������{]���s0yz!ʲ����a��P �8mFe{���`��V[Sg�E~j ��CPY�W��fV�E �n-��=���%��!����Y���^3g��%���a�US	�[�;f"l4ЫMR��!<��DR�RdF�&ա��;���RduW�3(�)�u0ͬ��b�L�R.%}aU�pG�"Y!�B!DHt!B��r8;"9���=�ti���9����g��Rk9�y$W��V,�`�ߐ �)�b����Lz[H�3jp1,v&#r�!e�f>=�$�u �>\6��nM|�g���f7��yiL)�0v֧��o�����G+����>?����6���DS�D��5I3�f����͌&�.��6��k�aZeᐣ�l��Ɩ��8'��('3�ӟ\�pٔF��K�P��_�xmX��x������}�3�$�膴1d}��!BV���ZR�l�F�uO�D�JN���kd�����g�~L.�౯���DM����6�ޫ���ˎ��@c2��y����� ��BbJ�ۄa=%H�i�19$1Q�������!��B,|o�WM�@JJ�;�B�A�h�T{��ُ�7'���T/*l(�v�wѤѓy�ߢ�V2�u���*E��Q3�����nGGG�I)�3��&=&���sbg�� VluK�m��T���l�g�te��4R�.�%� ��#�K�=W��Y]��j2o���-,Vt�����f/x��ѥ���r���%U�r�x��N-"���U���k�&%C�w]��ujH�D=��d�ݢC�ZC�`�����U�^�h��˲]�3�����%o�5-y�Z�Z��3��9M��2��.j��;����ؒ9>�G�<���n�f�Ţ!##��-NVV����uJ8E�A3U��1��h$�Al�2g�zs�\Y����̩Ei�����9mU<�r��-A��r'�7n9�2^;�p!�|8FKK��8����|wj�q�|29$��n1{����v�$�˳��É��?p���OLݝ��e��QE^b9u�%Ɍ���D(�`0(\sJu� �������5�k:����X6gy�C9�_��,���l�kwȢ{�ضG�݋�$^)Î�ƞ%�~]��t4"kGv�9Ѵ|�X	b 1 F H5l�-���~������#�!�����%&�a�����bO��J@8��.[g\���!�Y#\�vw4bB���\�ߍw7n���N^�����>o�$��)=��'�sLe�D�Qb`h&ڑz0S�R(�cլ�9<H`ؗ��v6�^�I �&��x^�iUi��${�3u��ze�N̚`6F�e�M^�%)�43,�z}��,�6L ���06��PX&C�ۉ���#t�1'����B��f�pgo��X5�<���8.3�T��n�P��Y�a$&����������]v�)�%Nxz�<��8)�d��f��q�U`�˙[ba�d��f<	�\����%#����f)�D}-��H8��{F�3()w�'�|�I#|G��	 HPf�ϩ�T\9� ���]��%p�X@��u�� �<ϭJ}7��L(�������q�f�Oȁ&�&>����Q�"ax��v�e��r
�Q͢��,�s�¹˽K���]��=+. ,^��ZG�@{x!�!��54)�����z<�I	.��&u�]ވx�VwT	'����$�r����&��E��4L��@�0Z�mt�J�!�v��4uV.�+U�DF�
y��<�_@R�l�h2�X��k�T���C��:7]Ë��ř\tn6��ih�d���s��P�e�φ�N����]��SCL��B9.����c}SI"c� �I���2�s�%2�+tn������g�{V�u�$�7Vgc���Y��32U,ݲ����w�p9�����ٙ�Xr���i��;d���ZIt@Y$~�/�}e4pA� �M��8�A-￸�($��6?����R�������Y��8�B���ۂ�|%~*7. l�pN��I7l-2�{�ƶ&���S���%K[$�����C\º_�9���|\��Ћ_���/T��H���	�8D�@�Im�P��L�&��b�Ă���ٞƱ{p�?h���GP��nL�t���[���?���/ڃ�G6� ��W���E"�?��p<�+�;8-ͫB�$*�Gx��bnq4`k	��RL����/%%�Ca��H��w�.�^>#uMQ�����aK%fL}H�~KI�K:��˓D�� ������q�ɐ,���$�x�`'��/\������"��[�q���B���PE��Cѫ����+�p�㵓Wm�����3��������/oo�M_���~��c	�qh<�J���'~�~W����C�R��^{�φ\'��!�5-�<Y'��E7=oΕ�I%N���)��������H_sN&����%�t��`�sM����U��َ�.�`�W"?�(Gf�x]����A*���'3��)��n�D�`!�1��0�xve����X���l���AC{�e��צ��/>;u�u�n��_�_�9m��
�]�Y���F	DA�UDW0rr�V��čb��,�MHNlE=n����/�abq^�e}���-<N�o�
,[b�b�-e;~q�r#��>�,��٩n
��D�|*��1PRr8(�� �y)�	�"f��,�ц�%ml��3>O.o��w�Q��]o�t�F�K��}�m�t�>aP*�S�T'
kA�M�d�����:1���K̅:�iy4��iS��$�$�GF7vFޛ?������}��~rI@9�9%�/(���J��0,���|�,�*�a�����;]�{<��|��!ƶ���C#��)���Q�[�W��ʓ�@1����_�B�F7�*U�)��u&��F9����R�����#��JG�����G��J�D��N5�@�锡�s�$��i�~��WVֱ�,��ݔ���&.^���oM�3P�}N�
��/ �%+�42�3SM`xS�n����4�XdPv��#�MG̗̰X�9|�R�,�x���=>Q��L�� N-��Up�X ����ƿm^Yc�����$'�ؿ�3$�7ʃ�7;������_}Ay��"�̌��sv�w�]���w$�6��_�݃�>�W��h�6�>bH�y���Z�n���V2��(��Arød���ӱ��PP�XQg���3~�aFx�+�9���aAv�&��%��$��/6�(���ir����5˷?V+k!�hU��/�ƈ!6��kE�eW�}�ſ�8�%�����|}syGb��e���.ݙ�̋�y���B��߅_ݨ��uԷs�y��{h�3(rX�P�[1!1߄��Ŕt�,C``Z�6�H��zq�A)N{hp�-wc��T����d�n�(G��o��{��S~�����E�W̰�Of�� ��i�l��J\��}�%���@�\��K�I@�7Cve6��"�g�nA�y����l�U?4��фi��$�-�y}x|uD6N�Vt�yeM�2eB�d��Y�u�2k��^�����HRl�?Zp�Uy�����5�����&��b�W�:�ȎȢ�$S����F��`��J����u=��N�����z��7���YI�6^̟����y�-ҧU�ˁ��qŢ3��+Ǜ.ʦg�;��TU��3W&)_�M�8�|b�L/��^@H�(tӼMwl����U�����ʰ�7i*�Z��u�<M���a9���/a����pO$�2S̝$=�%�T���Φ%�g�D��r��L�X��d�m�~	���<Y���	�+�TE��Ud��;�0���V.�� ���SNi�d�<������fD���M��V��/�3�i� s�|�oD�NX�0�}R�-Q�&R��7�%1�;�m��%��b�G �~"OM���'U���^4b�4�6��8�M�=��M��� ��?ja��ă��\H�X�S�f�BeK�XY�@7�a5��C撄��Qe-+���v~"���7�% ��������5dV2�0h�, ލh�6� Q���Dt�k���%�_��7�E:���~����y�?��W����`t��y�#�o�=���xZ��(j�bfcϲ;
����vj�Y��Mf�F�b���T)��GX[b�(��g�X���AJ	�nDWm�� Q���N�m��i)/�uE�7|Ac����Z�y�s�m$*lt3f��E�]ʌ\�[�C����q��u�=4���A�1����$�Ń9��v�xO�W�B~LGK�k8u<�A~�,�l\̢k�� '��h[�э�\+F���1+�t#�(�m����%�t��Xy�%�t̺y�uޝ��<�Yy2s����7��g�ۺB�j�x$���@��[]�`�`δ�7��\���q?Yl�"#[�Sv�������M���3��`��� y�����"�������B��<x�ԿL�׏/i�D���߿�0��&S��A43l�����fC�~��Y�Û�E�zq�ޥٝ��I��k;�1K��;{��㍓9��F����ɴ���+�x�xV�i��:����>��8���O�wox�?J�m���U����g���ț�.�'Wr�Y��|So����Cbu�H�w�Z\�������\�ǳ�|��ږ�108N�O�\�nɧ��hX>��	�$���y+�殰�.o�I ��;���㑊 +��-[�_u1O2��.��U?�'�q��ڜ~�Zۣ�����>��ld��j[7
�5��x �_x��.�C��ƺ���6��n�C*��������x�Ǔ����\r �|"��	^�a;�'d�u��+�_�����M���0��v!�1�GI�]l�kk������{�ަ�t/��s��M:y�!ϾƎ���y�y�Z]�%�Tɳ7.�
��h�t0��<���z#�.�B�k��!اIt�-�Gz$l D�\ꂗ��f^��я�j^��
��1�?�U�Q�F��.gܽg/~�|���Ixby�k*}�8�B�=_$��l��2�0�'%�cJ����K�Z�N�<�(�j2˗������E�x��X�ً����ٙ��̦Ц�/��    IEND�B`�PK
     t$v[�����  ��  /   images/2c98734f-75db-43ce-800c-ea69461525e8.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx���	��e}������]�st�3���#�b�uT@�5��!�f7	r�?	��pIV�b�ML�1DA�� �r�r�}�Q�un� YM8��y���~��5�pL�4����y�O.    {�@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@���#�^]޲��o�n�h���!˖�Bn��J����_�j��$$I���$Tw�����
!�{�%�B��{��ۓ�?������Ԯ��ݞI��T�ilI��ͭvcC֙]��uֳ�  E/��n�=�*�5:�A�4�_��[�J���U�i��h���������'�����6tS���3���\ҞJ�ͩ\�ٙud�ƏB{��b��%��n?��� ��@`h�q�����S/it�G�����c�fZXZ�؍;s#!����LxϑVH���P����������y��l�����ٍ����ܔ���Yc��b�w�~���Љ�� `�� �w~��W5�ʞ�ʕ�1r�n�����G�?��J���3�ܢ�v!��'���J�oXw۶\��@!4��7f�/¿�z�Kn<+I� �7���K��x���Px�l(TO��7'ɮ��!��v�3iq�[��Gxn��ϛz?��g���u�<X���ε��
��_��׎�+  sF���N[{m�ޜ}a-���*ϯ%�C�K�OK3͕�!w�T(ԍ�W������5UhO�Yh�|���^1=��_X�� �=B��W>��ۊ߹w��|\=Wy�}ii�V.��\=ɪ�l�����]��}g߼��{
�����2�l�e� �:�@�N��W씖�y:���C��[�U��^�J��dR9<��<��܎�3o>���
��o�3ۿ�����  �6�@t�<���˷����������1�.�� �mL�m���+��姽a�m[���kK��W_�j�ߙ �O����^�d�S=��yͷ�ʡ�0����G��s��	ݧ'����˺o.�w��r��=�ȩ  ���^s�_Z�,[�������KG��
Β�f��v�ѣv��Gmmt�˛����j����}˅��	b �@`��q����5�(�"ʇR3$�ɴz�d�������n�A�>�K�v����[ 0�: s�m�^�����Znd�M��3[�Ţ�]Z!-�HG��Q=zˎ�o����+5&.���_�� ��@`μ�c�|h���};����nr�����3[x��]p���w�K~j˧>���� 0: {To���}��L��)[��n�N�I����t|M:2��7��M�a�����:+IL``	t ���~�ۇM���ع�۳܂����h'!��F�;F�t�w��;�}�\m�y��	w 0���s���������g�$���93���&�k���[޺���*�����/�F �!�x�v}۴ߩű_ڐ�V�G�U����;��߸��-�o��?�����@�� �_Z�Oc����OM��u{)7`/����j�}��y�x����*����#ݫ@_� <�S>��e~0,:��OK"SK
�j��M6Z�����.�uv��ŧ���  }D����?.;��`��nJ��V r��U�fco�:�_�����S�5��}� ������/_����w�g_�NR�+�;�$)l͍�1M�v���//�6��E<A�5/� �7��w��٬�����_�� }����m��r����~�u_)�n������[ DH���������ژ����b��Ls��a�M���׼c���>��^|։; DD��3.��z�u֦��Z!��F��[��5����ε�^�\|��_X��  `H�r�5﹭9���\nQ�!�Hr#�sK�_ٹ��O:�z�/��o �e`ȼ�_e����6$�B'�P�N
+�K�����𴱰�7/x�17 �K:������F�hk���$$�7�i���N���9��o.�l���O��  �L������������%k����NB�-[x�T�����%�{���t �@`�:��]�`�_gK`��C6�5���򎅯��k~�/N?��  �@��Sνj�L~�c���tz���VKK+LW^�f����W���S��
 0�:���Mg�VXvF=ɍ���S��t[n�	����N>�?��/��  sD��S�^y�d6��I�9أiaѦ��ߺ�_ko�UC� ��ϝ��w��އ7%c�5���9�;.�#]xl-��I�}�c�|��� �A����'�x�����OMeK����'YuSa�{˺�~������O�C � �ЧNYw��'�n���i<-c�,[�(��<�jm�l����	<�����f��WO:�[��%|�� <M�Ϝ���%[��k7��/�̴:��,��Uޛ���1�jo�j��O6��Ѿ��j)�GWYesq��9��Wv<����	&��	t�>r�9_�C�U4��-
��L�۝����h1˺�,,eY�q�x�����f��~��|`g�y��fs��v=�O�Mߖ-<�4V��=k���{�x�:@8����l��){c��k��a���q���\��^�/��?���[��{���ќiu,�ẅ́�������]��#���3�Jod �t����]WΟ[KF�0G6L6��,yx���Ti��k{����Φ�f����[��Fg�����������3����y�����w �M b���K~��|�9�;o���d�H.�{�pU��c�պgk�q��z}���n��L+����SϽ�7.��1_ �:@�N[{m~{�}jc:����� slG7�g�v)��O��;���}{�Ri[�ٺg[�~���\Y�'��ŕ�c����/���� �:@d�{��6���N%��C��a/�8�l>r�|OX\�e�G����K�!s�o�7��Zo4��s�[�_5ݒ��y��3�9���w x "���U�z(]�g�$� �<�0�lu}��s{׷-��{��*w���hܾ�Q���Rߙ}~�S��_Zw��.x�17 x '�����>�`o�T��`�D멞C�m�\���o�=z��o�X��m�l����kIq�����t�տ���$ ���E �^vƅ�W���|c2�� {і�f���t�,������/Y]���ԹsK�~����A�c����ͅ����{��;�7]��O� {ѩ�]���F咩������	a�t��ۊ>��n.K�×�G,+zg�o�0[�w{�1�K�$$[�����?��/�|�Y'� :�^���/?rK���gCn,@$��ܚ�@�O�U�:�l}��ٙ{�n�O���i�:�����e��܇��/ 0�:�^p�9_��l���Y9@D6L��9��1V�e�88W�S�����;����,�ZZZ٬�œϹ�}��q� 5�0�N���߿9�����08�a��
��ü�C"�s�?s@�rԾ����޺����*�F�_�����N9��r�/��o CˋC�y�����M���t�'����wG�֩Vk��E��ZH�c��T��O�x��3��m��)�{��6W}��s�Y}���D `(E��`P�y捅�����t���\�>����P��ʳW��>;s��z#�v���Uy�����O;�C���7_�Ar��kސ�5�V�6L4��XV,��������J�����w�4�l���f��l�Mkοa�3�����6��"��л���E�ѿ�JJ��#�;z�����ܽ����_��1;��o�wӺ��p�7�󬳞] �0GN9��e�K�f:)�
�G�����l�5Z̲�z׳�^�/�(�����k��i�����n\5����5:�� ��� sळ������KkIqy�>�a��I�g�(�X��_�Z�퍾�	�Xv�#ϻ��/�q�����S��
 4�����?/;hb���=
K�����!K
�Ї��4{�!Ց�w4��[�M��{��dZ9��������eo�ܯ�% 0�:��������K��(@[����V-���Y��u�gfn\_����ӧ����~��s��֋>x�� �@� {���\�����Hr#�܎�v{��i��I�X�%��+��C��o�=3�y���ג��?��N=��^��c ���Һk��!]~A#d✁�q��Z���ׁ��E�\��g����}����~]M���}B~�߼�/.�g�����"����~�ۇ=���e=d�����E!�#C��]��qwmz�t�/W�{�'�־�K�����[ C�<���e�7��?_O�Ð(瓤����a^v�ƉVߟC4�w����|����������z�7n	~����� �C�<E�{�w�]:�����%!y��r�ˋ��cj�����7��M��V�����q��v?��ڷ\^� ���Ω��F��&�O%���m��)g��/��D:� � O�ik/_�>]򷵤�"���/Y]*W
ٮ�ȯ8�Z���;'{������y��\>��m��޲�\�矵`�wO����l�>3�V�,\���<��_8�g� }M�<I���v�t�kii�0�F�Iz��rﺪ���|�WR�~񇓓����l�D�5ȁ�S�%��ܲq�~͏fj��)=��>���v^��K/}�֬��s� <L�<	�����Ƭ�7�Iy�0�+�ݿR��������,�Fz�+�ON�%��zh��|^������������ˊ�%�,�ڝ������=]������ }K��3;������٩�rp`�B��tu��ߢ���� ��r��?��҃�@���;&]Z�<^(,(fY`�������퍾��#[|�;�}�O��}��� @_� ���u7|jG���0�YR���\��v(س�K�k�����ο�� �����=�W��3����Aka �v���j�{��^���L?mٚ.}��k�}��ӏ�x ��t��������-٢À�Vr��r��ŧ�����O̶۽���@�0�jn�{�Y�����P8��9����A���~��Ri���_�{��h����Nh'���_=��߼����� }E�<�w�{�[�f�Nj�H.;��J�ZL����$	�q?��>Y��>j�N������곇���YQ,����zq����Hv���S�r.���ٖ���'}�k^�W�k �ot����O^q̶����}U>p��ۛ|�>��Q+KŰ���ɮ���p��d��iW0OCo��m���ۻ����[Q*�U��z}�������ё��]"�4W��������.��W� ��`O:u�o��ҧ��;f�|����Je��=z}�X%�wp���;���p��~߽�Ѹ���Q>��U�� ��sIz�a#ի�˼��NnQ�x��θ���}��#� �� ��w���t�s�![��j.{e7���tN�i��B��}ۥ�=8c���zo����Go���W��s��6�zG9~�J��O�����ZR^}�L��o���7�# ~���]���u7]\KK���e������9��}Ծ���Z�u׶����=��oi���ڬ?ky�x�>�R.K�~��#��F�iz����>�*2��>w��C?�}�� @�:��s��k�d*���a�di^��|�xa^���"�g�T&�S����V�X�����޵��8zU����wB�_�vȒB����wզZ}P��ұ7��3���Ͼ�E� DK����?u��M�eo�w���U��G���5?͒�U��_�ejb��v$}�M5:��==}��z��f� �O�����ӑ�cj�7�>�,	Ɇ���y����೧��� @�:���Һk��P���AX�{D�����\�K�T���~�A��n��lit��O4���ɉ#�)���O��&����x5�;��/w?�c#����m��O[{���~� @t:@�^_�}�|A#d�0 X����7O��ߥ#����_�\~��t�����������hyq���e��8���ȗo�����%�e۲�_t��B  :}�`O����`���=gE���U�R�d7�����Z��;��Ƕu?'������S,�Oy·Υ�,��#^I�9ێ:ҷ'#��y����?p�� �"Ё�����;[�ї��v�����×����E�ʥ��V��M���7�M��=8;���V�g*WF��{6�Z���>R��-�S��#}ka�/�r�U7\��/�� @4:0�N=���lH��'�4I�+�TV/�B�zg�_~P���LNn��Lv�l�j�����ɗP)0���������#�#_�ujrG�+��,�V\�'����.��W� ��@�ֻ���E[J��q��j߮�="���ՇT+�,��C�z�`h��ś'&��zͼk�;���55���b�E����:@�7�u�WG�tk����In��h�Ϝ��pV�D�q�����kgCn,�����[�c}����ʃ��/�69Ֆ�<�n��o�l�^}p���6��Ñ>R���'�7�V�����;ݧΣD�/^��i'�w��6��/}��O��v#���^>����R����Z�G�e����-��8�R]1����+�7�z�~��ɨw�l͍��=k���_�~̕���/��<o���-����F�q��#F��:T��bo�wo�4���E�?�6=�3��ˇ,)D7�pw��<{�!�^�O5�!�Ho�i�9]�gg\x�q=�ȩ �^#Ё��K/�fw�>���J��������V�Ŵ/��/ޯ\�1�j?����(zw���ڶ��I�&�N�s���\�w�+�OO�"=�1
K�X��� {�@�J��?ڞ+�خ8?�煴����~�A����<��k������5;��_���}�m��<�R��S��^ؚ.~���{ͅ���� �^!Ё��O|��۲�o}���n����GS�%��V������� ����F�ޞz���j�F��g�[����R�2��IH�dK������@ `�	t`(�r�W�;����N��J�r>IN8l�o�Z?��9�WR����S&��z�!�|���	�V��7wB�9li��c������ld"���ݧo �;�����2��C���������۴�'c����+˥��_�	�86M5[�x���k�v���H��i����h�M�����tq��Y �Wx�Y{��<���.��B�$'Z�8�sV�[gZ��V� ��w��o��|��#��Aw/?�R��ujr�t�"�#�����������y�� ����@�Mmߺs��uk{�$��C���J�/?�'�.?��21Ӟ�0g���3�v/�O�Fz��"=˒�7���o�99Y�D7 ��d����G�OO ���lˁ�?](�
}�7�U*�Gs�0D�$$�!`_�a7\��y\�H���'�N<l��Τ�V�{��7�$�wG��l��:��}��~! 0/:0��s޷��Pa�Ч^��\^�8_C�����K����qm�n��r��������t���\�����55"�	�d[q�o�q��_��GN �@����Bҗ��G�[,>cY��Xo[��X-_�������1~��#մ��I?`,_x�d�u��zt��gCn����ݧ� �sH'���_ߔV}�������-�D���r�L�u݃�����`������T�tBE������ڭ'��������񉯿�/��_ �)����������>���j|@���\z����ΙV�έ&���z�'�b2s��r9��$�Mv/W���z;���ڡ�N�W���.��e_X���F�9$Ё��#Y���4W
}��uH����ڹ��d�re�Lk�w�8�����E�,=dI�����Y����/�65َlM--�[�z��u�� �3(����lM�l�X.	��\�@����:�R��-��F��~s�+���V[PJ�e#��y�35�j�[�3V�e1ޏ�3��=�����^��6 �D�|��3���ێ��K�����Z��W\�~鶩�V[���ڝN��{�#��ϝ�Ύ�V��#dK���:�nm�l�fZq��TY��-����� sB���W�wcZ9$��g/+/�ujO�ґ\�����wOGw%�����;���p��H����t���s��S���n�o��؍�~�>pG���'��Ͽ�W^�� �'Ё��K�.߾sY�]����zӛ���fƖ�f�WR�-ӭ�w���du�2׿V���l�魈wC���Vk�z�~�ӗ-���I�fJ�~���� {�@[��l>�8��J!M^y�H%ILl�^��R�1�i�hG#�+���7��{o��w��΋��E۵M�����w�a�L+�>����y�^�� �%Ё�w��_�k~�χ>�+���T��$����"9�j�7��1��(�����ڒ�,-fOv�Cg��no���[���S��+ܙ_zƙg���g���z `��@ߛ]��[!�딎ܧTZ1����|�WR��͍C]J�F;t���6�sG��<֮�A;/>�f��[W�����? �1�k'}�k/ؒ-zq?]���h.w��R_�����,[�0��՝ݱi�ٺ�������a8/>�&r��<m�<���w ���������k�JY����]ê�;�f�����<�S�����~f��-��a9/>�Ꝭ��~���� ����_<�cHF��H��r!�7b�nu:7o��~���ن�N��v�3F��9;�coz�'/;�s�r�� ��&Ё�5Q����&�:�/�8���ݹkK���k3S�1h&Y�^\�[E�� ��&Ё�t��M�ȳB�N�'�KVW�w���h4��o����j *;�Eo8�ܫ����tc �i�@_�*��V'��b���A���j�7u<�4Z�����gn�T���qj��X�U�[�� O�@�Ω�\���قC�e��ˊ��T{����h\}�tm�vv���l�kO^��}.>�� �2������Y=�����ʁ�V���ݵ��@_h���H�n�� O�@����^�ƍI���'�ݿR�璾x3!wo�ׯ��V3����l���=��U�9�� ������X߬�<V��(ok�n�]������`��l �R+$��aQo��� O�@����\�I���
Y��x����a[�ٺ����3mg͡�M�_s�_Zp�Y'� <i���ҏ�˽�/\Y*���O������Lך�`K;�f�U����s�� <i�'������ʋB�d��ˊ��cj�:�n�O�g���o���?�5� ��"Ё��Z0vF;I����[��~�����J��Л��/wLMm�jz�h6��m��]ݧ�+ �D�b�w�q[n����PX>����1l�n5�����)w��@��-�� ��4/"���]��FȢ��KB��}�����o{�qŝ��Λ���N+��o������� �m�ڙ�N��������O�X)d�=�[7��^}_���axԊ��� ���D��O�ԙ¾�!r�|�>{y��)I�k�a�Í�� ��t�9����G|�W_qK `�t jS���}�+˥,K��i�+ݺ�.�a�C'���������"Ёh���ʃ7�#��ȏ,����%�|�'����9��l��N[{m��ӏv�"�n�@�f������=��pV���	���5�s 4Bnt��Z�}zq �		t Jo���ljb�+C�Vs���
�����O/�/�sj����x�t~A晴@��R~�o/�C�^��X�X=D�kwLN߻�)΁3�T��;�t��?sg �q	t J3����[^�r�.�;{���;s.΁�wTi�S:���� �K��9�_9pSRyV��Q+K�U���=X�1�x,٢��t~��$i �@��(����
.��p�,[� ��y�m���=8; C#�/����}����$Ё�L�"w�>����!ܻ�Q����Z x�ܢ��@x\��ɟ�ƫ6��X�آR��8�������wMO�`�Lf#�=��/-���w �@���/X"������^���_�kz�ݑ���i�$�Y1����u�G%Ё�L�#/+����POn�u��ݵ�ZC�O�L6�sA�<&�D�?}�[��Q�_"�̥�b�������h6��T˪�z��]��y�� � ЁhL�+oY�V�-�×a�ݽ�^�y��Ԁ����l�pr��9��@�Q8��I��ந��2�/��I�׿ͥm�f����<=���k�@xT���~�u��BĞ1ī��V���;������9�LuJ�<m��K�?�� ?E�Q���%Dl��ec�lh�f~��Zm�l� ��v�f�a�w'�' ?eh_l��mo��w�(D�ˆw�|�D�q�s��4�Tz��:��#Ё��s���Fy���|��2��N�wM��k��ZR9���~��#� �F�{]�0���C��\���j��_��ltlm���4��SSo�>�| ��t`���娷�w}(W���^oܱ�� s��U^:�O��^uʹ_Y�))�
�ZXL�e#�lضx���_uom: ̑Z:zd �t`�ʏ��B�w��Vϻq>t�ۯ{�6Skt��}	`�$��_����_�r� �t`��	��B���Ð�1�j�pSc6 ̱�b�M�:��	t`��]�v�w=+Djy5ˍ�,�o�W��-�󠑎 �7�kn�ؿ�l}�a�^�v�xa�V���֨?��� �`*)v��_�^�'�n t`/JF�O��:�Qn����t����L �'���;##��6�*  Ё�g&)� D�7��RȢ^7~��>;Qo���W�l�A��"Ё���3o,|;)��:`q~��>�]�v����yW����"�o�+��g��Za4�-��@���?�T��i�̿Z���9t���P �I��!Rc�,�ҡ���lY=��v����g�O� ��@��zR~^���E����x�F�����ȕ^:�@����tp����3���9�zRzn @���=�}��'�(�?/dI�l$?4��o�zD`:)|f����$n� ��@�]#�{u�Ԫ�\��}�u��sӦY���^�L����Ƒݧ� CL��n��a��ʅ�3���m��t�m��B'W�݇.Ё�64/D�x4�ʡ!R+F����x˦�z ��lVzA rC�B�C��MIqY�-�V�I:Z̆�����V롉f3 D���
 CN��Y,��:i��0mo����-`�͆⒏��N<�l`h͋Q i����#�q�y�j��7� "�$dߺ�����k����@<ZY����ñ���m�z��j5 B�j��@��@�U=�"T�'ɂb�C�޹��9�VRxf b�W���o�вJ������>���Oĩ�����@�ͻ>v���!��-����{�7n>bUO�|`�t`�$�/	�Z62$�Ϸ��ī�FO9��e}�����i&������Ur趷��v�	�ޛ�_ CH���	)�i>Q�;'���vV꽙+Ё�$Ёy�L
+B��+ñ���m���k%�`H	t`��;�x�s҇!�ۭNg�d��v z���< )�̋�\zu�Ɲ�j���J:���q��l���f�[ ��@������C��g|q9���MX=��l�_ ��@�E��<#D�N�&I-~�?��!Ё��
I�Uk�����hv�C��vmo�reOi�:�MS�V ��V���:0t:0/:�����t�W�{w��;Ο������� 0d:0/ZI�O�Т�pz �#�;  !�̋f�_"��4���7����vV\ ��@�E3�9�w�0�+�[:�gInE B�so���l�ά"T)$���V{�� :�_Z![ ��@�\a��e�\|��{P57�+�[km��@��d�(���k�{��O�_mʅ4I�$�7��m��?�NV C(���IC�ܫ�t�ϟל?�O+$ŏ\zu���[ CD�s.IQNp�擁�-�M����O��ܽ+ �̹vȖ�s������s�� }�P��&�t`�t`�u��X�P��t���N� w�O�C�Uk�����k�tQ�P1z�{����+-��!#Ё9�N�(�<�[�'-��@�ju:Q�/�K�s�$?"4�gЭ�}-��Q sI�s��	�a
�����zK��+u:0|:0纕��ea��m�;п:� ��@�\'I��B6�3��t�k@�jE��.�\����t��D�V��-��V����$�:�s�4��kM>	�-;܁~�f:Q�hK'Ĺ�=˒�^bn�;���>�S���0����t�	���������-������vb|�>���wi��9п:��@��@�\����,��>�=�ٶ�����T`���̹v'�.Ї`��:��ډ@��/|��KBt�g��m�ہ>�	Itǣ �@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t ��Ъ�;�N�7?�$I�Y�X <� �:�V6�c�ҽ�1���Lelņ ���  �!W�N盍퍩� �1� �8�#�vtZͬ935 `	t �'PZ0�m��̷��  sD� <�$�-�4����V� `t �ݐ�i��x���-��v `�  �)�r��ek�֯��a �=H��N'i�N���P�MҬ5?�V�^Z�d�޾~��#�T�>[�ٱiI���`Y�<ջm>Mׯ0:� ����j��/��2�|�V^�l����]���&�H��JgjS�F�i�/�gʋ�mڛ��� ؓ:��h5����t%�Hs��޵g�������5 � ���:�dvz��l5�5g($i�譜��=p� {�@�c�F#W�M�V͝5g8$i��xņ��ؾ�\��� ���lm��l�m�ex����\.�8Į������S$��L���z��:�N`X$I��B����N��ֶmX&�x::@i���3�E3l:��P����|א�v� ���z03=Yi���1t:��K7e��l�Q���V�Mp`O� �s}ì�`|s�T����K��z1 � �b��4�\ad�|yd:D��}�Vc� ���w'�����g�S{�]z�����E�I�k^u��'��,fИ��Q3
�fU�q���M4Ƙu�5�d�q��;�
B�i���]j�:�3��b��roU=�����*���Kso��ճm ��i�u^yn�+�:b�~��b�� �T: ���0�r�Zӫ�[b(��:���  ��t 0ǧ�I���W�b(��6��5 `t 0 ǧ"�W��[V�PA�Y{��  0": Lǧ�ٹ��8�mY�;��X  F�@�	y��4�4�a�ٮ��/�e)1P4���- ��� 0n�<�vsA��8���As�8 �� c��i�wY��8�l;�� ?h,m~^ cB���p|pˎK;�8wb1P�^�8 �� #��i��XVR��~�r�H�D�;�s~f cF��q|�(:��tr^(�o���n��
 ��#�`D�n��Fp��P���C���@����ځ��\ &�  �D%L��k�n�8�ǹJb�T L�  FΫ̯��R_L���o,mM��M E� ����sk^���8_K�<��+ 0q:  �\���*����X����  `   ��[(�󕹦j�\^��AI  0�  6��/u
�-�b(��:� � :  �T�W�綮���N���5 �0:  �4v.?(�m[C�f5�6�  �  `Sخ��/�e)1P�NcA  0�  6̲��hr�z�Ake�  `0  l��D�ŝ-�N�@��/���
  �#� ����4�=�s'�� �p�[ ��t  pj,+)�m[��\$�� �o,m�l  t  p*��s��b�$
������9  Kt  p�T�����|1�Jb�7���  2�@  '�P߲�J}1�J����$1�8 ����  �0�2���=1�0�W�oWI�  2�@  '�+ϭy�ZGL���o,mUq�	  E� ��ʕjM�Ro��t��-mMB�   d�  W�Xi��1T�yh1E  �t  pLN����W�P���B��� � � �Q9�B�Xߺ"���ksѠ[  ��  �v=�8��X���F=�� �!� ���7(�o_25΃n�v�s ��!� �#,�	K;�,�N�@a�]:� `
�  �0ˎ��y�(�~{uQ  �R:  H��J�8?h��H�� yhk��  �� ���q>�����B1P�q �:  �M�-9^>%Q��K�D)[  �r:  �K�[9^�%Q��V��8 � � �Q��[(��@*���ځ��9 `��  � �2��+U�b �$v��4�s �!� �1�r���m1�R���$
= `��  ̐\���W�b�a�/mM� /  �  ���K�|maM�o,m��AQ  �Q:  3��
����1T�qh1% `��  L9;��-�����|��* ��#� �b������KbYJ����~�&  �@ `ZY���۬��V]  �� �4�����cɲ�D����X  � �ic�qi~�A�vb1P4����  ߃@ `�XVRL��vs�(���As�8 �(t  ��r���(�T�$�e�bٶ�k�m�:�x��`�4���-  �A� 0T�a%E�|}ב>���n�N�8N����}��F��Ł���s  � �Pn�i�npܿ/I,}ӏc	����mw�����S��$
�a�+e  8& ��SN�%��o�SVE�x�u�>뎛Kt�;���%��[;�=}�  x\:  ��|[�\\�/�w;�����i��]Ǻ��{�$voe�vIb�7  8�` �Q��:i��� ����rK,+�͋Jr  N� @)���u�@JT��9� ��C� �1i��-��PV8�[*�  � �Q��q�SE:��  ��F� �ʲ�b(�k��  N	� @Xv��8��PѠ��yQ  �)#� 0���H�Қ�D���l%QI  ���  L�K��&��yX��"  `�t  �y"�Қ������`�~M  �� � 0�J�W^ˊ�DI��pPO�>  ��@ �0:�U��f��RI�Ya�n�  l*  ���n���T��8���s  6� �A��oY���T�Zq ���  B9��ع��H)G��|Z�  �� � 0�r��4��b$e�  �� ��);�M�'R*��h�ƹr  �� �%�ӷ�|G�DYv4��k�  �/�  L��݁�Zb(�[{�9  cA� 0ʲqM1�>JM%�  ��!� 3%V8<�\ꖊ�  Ɗ@ `����4��,��Ȋ��$QA  ���  ��+��\"�"IX  0:  c�y"^iU�J�DqP���,  `bt  Fl繲�q�8�  �( �R)��kbY��(	V��  L� ���8��nّ�(���b��<  3�@ `TrŦe��H%�gG�9  &!� ��b��H%q�
�si�S�  �@ `�%�׶��@L�׊�sq �qt  6�r���x=1�R������m  �!� �$�v{�x]1���s  �F� ��\_�|[�DYV�O�\9  �E���(��P��q��8��8�k�  �k ǖ$	�p̀4�b��n�*�	2+�#;�"�q�D  S�@�ͤ�D酴�	��e�*�sc߉I��R�'�4�>���M/�/D�R9 ��"�`��Q�0�D����ͣ,;J�|����Ѡn�8/��?p�(t
�J�h: L' 6A�vȨ��Pb�bp�[�_�$*�NǖM�
�(_,1� S�@��PJ� p֛ό��ɕ��6s3�+��E�T}7�#�X���m�F ��� p���>{�^��Ĳb1������e�L�3w��������o N
� ��)�Gǹʕ�,�6sZq�8�f�J��i1� �� 'A��Li�Ej�[��b�$,X�_�,=�=�B�T�2� 2�@�Ĕ�٥�BӲ�@L�Dy+�낙�D�p�{1�tvy�l"����V��`�('����@*�sVد��{F8LOy�ץ��\�`�^	 �c#��8�0�#֛Ϥ��ږ�닉T�Zao޲�s<֠���ql��κt � ��#�f�r���x=1�R��8���bc]: d� G�z���z�x]1���q.¬�#��+��q" G����8�����3J��@�|[���y�[�D�����.]o�y� `6 ���q�3KY�/n�)R�Wg��9!�q*������������������ � �fp�-��@rņHǹ��\%96@o����K�o+�|s��e/x��n��;^�^�@��LI�[VlY��5�j8U��pSXb)�zmS7�� ��(��b%���	}W)%Y��=v�֭�����߼�����K `�� f����8n�#n��J��C793�~W��o��Qo��6�N�]�;��i�r%��Nپ�;�O�~�����^~@ `�� f��5 �+|'Q�U��1\ǝ����v�7n���4~� N�`&�R�����px[�Z7>җ�m�/����L�/ 0�t 3G9��urIR �̼��ҳ��Z���s������+�/ 0�t 3exp���I��� `e&�-K��~ޯ��w��#���
 L��X�s}!*.�� p��H/�k�e��;9�����u������ �":��0��N�K��ܫN �0�n���t?Wu��_����4�4!�L=�(��� p\�H�<�ww_q�V���[��>|� �� �L�~���� N���}���L?'�n�u�^��k>���~� � �L5}��/4 pR�9�bY�P*;�<�l��������ο��^}� @�� �����& ������,K�Œ���e�ۭ��I� 2�@0��~�%�`�Aߵm[��X��n��ԫ����;_�� F��:�?p��  6Š��Y���\.CݩN��_������{�	 d� �JE��� ���w۹R�8���@��X�wj������� d�`j����  6�R֠��J��o�f�Z��-������>�T  �t SC�u�#]  #�ı���4����ծK^�_�u��� ��T�;�s�9 ��>�Ro�i����ʭ����]��Ȼ_�J_  Ct �ǎ� 0^����q������� �@�Eah�c; ��ސ�vs����ݭv^�K��O~����� @FpQ ��z�A�æp 0!�9�\��=q\��~U�6/ �:����l
 �����{�ʕP��n���U���߼��/ � @&����7* �D�=@ܜ���g�z���-���k�}���	 �@�9q�A���v 0Ġ�uˮ�X�m�z��-;w��M�+ `8@��DI��&�� z�Q/}n6u=��j�~�uo�O �@�)~�˺s 0�^�n����l��古� �@�zj;���������M<z�m�_�����m �"�dS��|��f��~�����X:�L��&�� ��S�C����vuo��?��w~�o���
 �@`���>�W ��~��G�����]�����_��g�V ��`<}|�  �C)����J��qSݻ�z��ƇӇ�( `.zMO���% �)q�Qzss�Dsw8��ko�񅌢0��Xz͹��v �,�a\�>�aznݽ��7}4}�| �p��Xi�;l ٥��M�0�`�g C�0R�����( �8S7�ӣ��?��/���� ��/ #��.g��4PJ/Wr
��q����SzG�0��8zS!���  ������;�c�(���X|��������� �t ��=�� `���[�TC1���U���\0�=�X5 �>Q8qŎ�u��!g��/������]�i�	#���s �^zGwǭ�eˡ��G�ó &�a �`� �[�N�P�L[��/Y8㗯|{�Ϯ��+ 0A: c0z �/�]�\1j-z��vl} }��	�b�=�٠G���Rdڹ���O	 L������ f����F���-�_z����' &�b ǱŹ� 0;LEW�%K�w}��@01:��ӻ�
 `�Da`��X�?�c'w E��8}6�  f�?軦���:/x�;^�w�� &�@0Qz�\%�% �������n.gԹ�Ka����`"t >�� 0���5��@?��� L�`b�(�h5 �a&n�%��W]���~�[ ƌ@01l ���F�E_
���;��� &&�8Z f��(Դ@_U�� @���1�� �R�8�-�q����s��/]������_�	�1"�LD��p �����X���H#r^�>"���`"�� X�_�b���d�1#���� G�����I��7���~����7}M `Lt c��� ��a�n��Zw�t�M�J `Lt c�w�  �`�n�l�1"���ީ��� �G;<�]�e����� ��`�6� CG�k�1Dˮ_�w����W� c@�+�A�  pq�nΜ@���u������� ƀ@0VztD  8
�[kE��@0&:���>FG  8
�[k%�Y cB��$��s ��қ��z'�W Ƅ@06�? �i���N%��W���g�_� 1�ذ� p<��V$�+q����� ��`,�ٶ�? O�ƽVt맅@0:��H�ب ��������ۉ� ƀ@0l 8Q�a��}�� ��`,b�, ���n��1 ��E�q ����6��}��53�����X(6� ��8�g���9����|���ݫ�- 0B:�� � 'j��a;b�A��LzG�)��� ��q�uì@�i #F���@ �$�����j� ��� FN� ����Y�Al- ��`�L�� �O)%&�,�" 0b:��3�<[ ��L[$vQ `�t #�w ��2n]\O `�t   Ǵ@��	 ��`�ҋ,F� 'ǰ׎ز��z L'�ș6
 ��J�`�t   Ǵ7w�e� F�@0r�7�� �]JA0z:   p�8 �F���X��J�}>�����J,�?�Ob9�,�2��,"�����)�����6�R�V������ `
��)�la� p2� f�`��Y�\f N����!����� �>�,A0:��S��  N� f�`�� �ś� f�`䆛� pG�A:��Sql[9 ���Ĭc�X�`t #�$��  '.�#� Ɓ@0rI� ��G#� f�`��0t�� 8i�S� f�`�(4j `�$��
tF���`�8&� 'L%1ר fO~ F.��� 8qi��u	#� Ɓ@0I�l� ������Kt �@���� �G!ר fO~ �"
}�� ��o�5*�� �Ũ'? �+�}7_  �+
C���@0.:��H/��� p\*I3�XS �F����R�mYv"  C���@0.:����Yn~   C�f��N���D��y: �q���S 3�'@ c�9�T  �%}�0���� ��QO� �[�%*�Ա�( x�$
�J��A�'���.�u�/  <J���b�� �C��(�= p�?0s�8 �X���:t ���Pb���� �*���Y� x4�ן����N:���8I��\�/  <,�{1̑��M0:��z�B�N� �k��zb���� Ʈ���
��� ��8��(4���s �@�;�� ��E1�`t �4w �:��s�9�I �L���^�/
 `��Q`��v�t �@��=�=E���l��^&��s��q �L���KLs����t21��u �@���~��j�Nz� `�DA�Ǒq���s �B�����.{�ZK  3g�i��0���$�D�ڭ|� �-*�]�w�0���$�D驍l �GϠ� &�@0qz�cy�@�Y�k������ &�@0q�~�)��e;�  �^���IWÎs���`t F��b}qM  S��nw���:�I#���m�
�9ײ�H  S+���0��[�}���X�9�1�^����5 0�z�qG�i�7�]��>0z: ct�M/_�;bY�  �N�&�����vK�Q#�Co�����|y�) ���o7�<Z�x��Z���9�Q��f>_���C 0E��/����s�DF��`�t F��w�5֢�t�6�*b��m�ε��� ��i5<�T�\t ���sSG�Odz��J��( F�@`�^k�Z�ۺ* �LS��Nc�ȝ�Ot�\�ي7����H�^�-Vj�� �YA�U������'�DGχ�ľ ��� ��i�Vj[v� �Q*I�n�Q��蹖��� ��� �������|�+ ����jz�O����Y1ˮ ���h����b�c�  [�(�����dG�5�N ���hI[��j�X_\ @ft+U1ԩzޖ; F�@`<=�/W�0 2��6kz��Hǹe���u���9�#�dB{u�Z�~���� ���8ʙ�1�v�k�5K%��� �� �(��v����5 `�nc�n��p�2�]+H�ﺗ� F�@��V�����8� ����9�];��s�(A  0:�Li��U��\��2sx f����n��P��Z�9b�X� 2%+�4�� �1yj���T��ke;�O `t �����^��x���Ncn���+��W ƀ@�I�ե���=�XV, ����~Q�q*�ң�r�ڑ
V�� c@�Ȥ$I��zp���cY  ���i�.W�`=�+?yߵ��E�1 �d��N�Zu�Tk
 `캍CsIolxz�t�ot��n: cB�ȴvc5�������N��� �E�A�����n���� Ƅ@�i�͗��E���*��i� 0rq0(�7H�`�ھ��l`lt �v������]K�͝��[�{�  FF�w�\9h��s=r�ѩ횕��T�� �	� ��ʞ����5b�$�S���F�[���� F@��n��S/)�a�Y����y�� �	� �.:}A�"�����3�s�0��Z�8 ���Z����M�͊sm��� #@&r�\�����H���Uk�������C< �1��ڜ?�o|׵ڬ���j��Y�1"�dғ��Iε�z�%~����*��F'�� ���n���6sj���/�\�; cD��'��'�?���"/�A�9�ϩO����	� �*�{���JQ��q�դ�����) 0F:��9wgM*����a�I^s�ҏ=��>sG�K���K"��\Y*��t�o��vm17xP `�t �s�'��)���Ÿ�������j p(�7�����s}�l�^�? ƌ@�){˲�Z8�a�$I�3+QMΪ����� p\���ơ�ue�6���|������$ 0f:�L��GϏ��H?�nׂ����m 86����9��=6G��v��v�K_�, 0f:�̘/{rƖS[
F�}�B�Ǖ���� p*��4���82��sm���m��$ 0:�̸d�l�j,C�I[ܺ�J�[���  �����|�����֝k�JT%
_' 0:�L(z�����ᏣG�u��V�) �!=r�<�?#�Zw�n��^{��l� �� 2�){����o�(���z���毰���Ҵv�uG{��=��� ��� ����Ii�o&�N�T��z 3J�֮7�#����k�u� ��� �w������_<Fql�H/��}eY��)*�3��n�V��|��/~@ `Bt F��b���j'*N#��i˕�@,; �I��Բp��6�ۏ�3��� D�0Z�����7�ϑ$��i�
i����� S,����JV�|�;�����	{��u�	"�����7��^t�������Vw=�7 �Ba�]m��%#F�c��v�ڷ]��� &�@0rz�c#s��^j�?�r8ҭ�q�cI�N;_*W�F�qN:���Z�vc� ���G�)�#�K)Yp�� �0���я8�R��Ǹ�`[�閇��O�5�H�zݎW*�,�� �DY���\���IF�3εmv��'���g &�@0�B+��E��Z�#מ������~/�ő](��X�	 G���Y=8���/��D�sm�|T � :��ٌH�����Q<�����H#='��R�R�6 ���0�\>X��1j���%	���y���- G�+=�]G�FܳԑO}c�<��Ӕ�6��$���f��dI��ʭ�C��Ծng�?��֭�=����t c���p��~�rG>���/٣r�h#]��a+K!���.����j^2fq�X�{�/ �@0v���V{�H��Kv�|��U�^��Ob;_(�.�q�J��ڡ���zsmq���5��+n 0�`"6+�Z��_�>�Oݣ*��ȯ�|�wү�T*Wb�9= 6M���ʡj�֛k��sW��Q�� �At �Y�����/�t��̥{Ԗja�Wyq[�V��Fz`s^:�	����G�T�k����yߛ~� !�L�fEz׏��r�p�����ȯ���n��y��S`�;�I�G��-�gqJ�6�8wT"���� �!�L��@��r>�m��w_�_~��;����c��|߉ðT,W�������\>X��.��&��n���W_�Y �� ���ǉ���Czڻz�9[eW��(�n�U(K���l^.�%�
:�z���$�&�v����f�L �@: �lF���k��H�ʳ��s�g�?���=�N�X(ˢ�l�$
���C�(
3�����i�N�������I M�Y e3"]��@K:�P�{�nUλc���Ў�F��t �e8j�m�:�F��6_gJ�;*Q{J>;�0��)�(�\ǒ$;�l�/��=��/>M�+�%�M�P*���T�8̷V�2;j�������7?p�K># `(3�-�(��o4��������٪.=sql�a�Q�Yd4�ɚ�QsͶ�G��'-��x�|�9 #�M_���=���R�;����=��2�u��� N���B{u��AfG�5���������\�_ �`: ��<�=+]�����t|y�E��z��hz�j�B��97�c�$q�Z���Iƙ�5������~N� 0� ��0��nw�5����=���T�쬍u�����K�R9t�\( ���jkm���s͏4�cԎ��R�^�����wy`�t ��雱�{%��W���]�]���d����v�\.��%��3L��i�T��7g����ܑvX͵��%� � �E�8�`���i���ol��6d�5�g?�45W��:�s�H�f�P,F9��g��	Sj8���ie~:�f�fpGr�X�Yjs��� �d�|%/�z��Ϸ�7��t������٪.:ca�������z껞��P�I��rTR�YbY*V�@�&�o�;�i�ή����H�V>�u/�� @F� 2+�s���d�������;wj?UQ���n?(�-wԳ��KJyw���>�ݱ�\�Xb}:NN�����̐DIK.3�>�����k+�8��Z��&�7_7/���~����o�* �:�LK/����U�׋��7?(�`cǱݷ���?�;�[+c�ꌓ�����lb�>ȸ$���je֙��Q�~��Qr^�����L6��):��p��������>���@������#����svԆg��z3�>=l6�^>�E_Y�t̅f�J"��X����y��7����Gz��z��t� 2�@05jE�z��U7~k�|��Ɔ?ޝZ��ZO~���mՉ�路��yq�X
Q̧�8�o�U����]g�<�}]M��S��~�� �g�^8 �6׶��x�irƖ��L�pcS޻~$��ƃr�is�G��&�Fӵ ��V$�sMs��>�}���\Xi]{��/� d�Խ� �v�κ�c����e�jo����r�rG�q�6u���ĮP�C=���y��F�S�{��ʠם��,Li_wvn�;���� Ȩ�|! �V�Y������V���9(q����k��ǭ����.�!���˄��路�u/_ĲQ�H����ά%�/�v�^�ml�SeaJ��y���хs��	��"�L5���%{e�|I���J�l�c�{�#�z�\�wA}�Y[Ķ�I�z����P,��؜~ �˱m9�nU�����Ç?��P��ǯݳ"�BG���pU��2�W>}:�)03��� ��^�~�g���A�#���M��]�r�R[~�j�|i�CLA���8�����'�#�i����',؅b����w�F����&������$��=�EOg��l�����_���}R  �t 3#��֏]�Sv/�Ӌ����6j����~�>9g{M=�mR)�&�q�Q�-+�甼�֤}�J?JKՁS�Xv�s���sN�=�l��vխ�����M�3[gܲ6j�n����o�� S {�� �AO�Q��,������|k_C6ڮ����@K�>�N{���E=v������ ޶]����F��T�����Q��q��Sw��.8��e[�v�?�����ܫ>�ã�"���ZU�2�~�)A��Iz�곞|��ڜ��o>�)�]���o�ߒ���U=a{U&���RJl	ݳ�R;����o�r�J�<��'2���Ӌ�f�(�4Wt����޺��]�k�s�9O٥��
�צ�<�%��暣������w�K� L�l>#�&ٽP�M�?w.�7�]ݔ�f/�O߼O�׋���m����u*I�eKvU�� .�}�H�8�?�z��O�s[3ȱ-9c�-�=g��h��J���g.ʎ������`3��l������������%� �":���צ���;����h�j�ߔ�{���O?{[U���%ψPO�D�Wrμ%�.��v,�7y�1E<cF�{���Nyw��,���R�t���3����ZOL��s͏e��z������
 L �/��g��޽,_�{e8e}�t������s�#쪫���e��I%��,���=%y��=��,�|�1u�y�:k�)�Yw
UO���q5�$�����N���{W&�F��ή�<+�ˢ���'}J `�� p׶�|�6y����l�?�ܔ�'J��`c�>�){�ԥg.J�s��J�k�EEi���EO��ʽ+i�͛����cY{�n��9���l��K/�w#�Ŷ�VP����c?�mF͵�D��ϸ���� �B: E����s�n�p����lڴw=*��{W��~�rIz�rf]4�O�?kΖs��Eh�r�J_�~,��4�Ϙ��kvq{I���Ƽ�O�X��էnzP��p۴���D]Ti��o��[ �� �����p�[�_�/޹$�&m��?Η�Z���[���>����Q�Dq,E[��[.�R�Ձ���Xl����BO#?��vV�����Q�D����~�����ޑ��>-������ʇ>t�5�@ `��w5 �ql˺d��R��ms�6��X�r���tߪ<q���]����I"uO�>�����-K�Hj���1N��E��Z��Y���*V~� n�֣����$�"�H�C�^�����~4�y�_�ȵ�_. 0�̼
 �i�?y�9�������ou�vd��Qu���OJC]O�sb*�$�5�{jyQ���X�e���e�w}-f��ڲ������l�8�#����	i����P��[�Ϸ>�qTG�M�t�#����[_� 3�@���c�d��8S�_���~@�ۛ�>]��[�_�'��S�.��ZAL�c]�ۖ���Zp䩻�d��ȁv�F{(�����/��4Wtegݓ�UW��]��������,|W�Hݜ�<��A8�=t��۴Lg?���|����g��@���nw�`R��)s�����o�א�ciSG�t�ޱ�5��/���}^X*&���U͉Tl9oKQ,�"M_�j/����`3b:<���9����ֲ-�+9)8�7x�(;'
4������ᬘhD;�O�:�G[�:�9�|Ε/}z_ `F� F��-�s�zP�[��e�2��w��9;��{W���u�页�𶥚n(w�κ�N6֗&��W�JU��/�]�V�Ix���}M?:�
cF�gW����4�Ki�W\)�,�����D2�^�R����p̃�ݑ�w>�a���Apn�{�u/}�� �!���;��b���������P��k���c[O;{�<qϼ��]�r�k�>j����[�w�ǿɓ�[��I��]���r뮸��ϟ�)��j_��z*\����V�t�(KY��sr���m՜,�4�]����2��D���F����|���6~�t��Og�fE�������k^��C��w��W�����g|}����U��瞒�Z���ƺ���ƽ+�v4�:�������M���ޭyʞyٳX2~���$Ib��ϙˉ3W��=gU�=%�'v�$�r_��A�ԉ�^�S)��X>��E[��{[%G�IK����������M�9?Ҭ���O�#�Zo�������
 ̠��H`���7�/y���km���[��m5|���X?t�6����a�����:r�^jo�bn8�~�isR�g��]���~����I.��Λs������h_�+��k�(i"&�@�5TK��K��
���v���$9"\�X2��Cz����D����h�F�R�k������׼��W�� ����U�Lz��W��K�������_��TG������n�ou$��5��|��C�廖�������˙U4=���4Q�4����(���8��V��N��V �j/J�0�EI���P��w��Fx-����zd��G��z�x�k�z�\����Z#�>Ҭ���X]Zi��C�\�_ f�`��w���������}�Y��=�����:�/ٻ���w�8rI�~�������>�͗�2Mt��ǧ�^��-�%�-/e�n��^T��$�P⶟�M?�w_��^��~��~���Ǔwm�])�l�x��=+��4��8�sl�Jb��?�^��r灖ܶ�)�ڃ��YsM��_u��^��� �q:��x�^���Ho��n�F�k�������E��PS}��k��y��3�����ێzQ�KC���5������pC;��t��W9}�rZ�[\e��怕�#I#^E:�{���A�:i�u�X���r޵-����;�~��ǚ�]!�i��ӿ��mq��S��'�׏�t��Dݳ������]�	��+���8�����^}��	 �@09:�/�/�z{�#˛�!#׶�ǳ]���Yj7�{`�;�ϧ�����sPN�R�sw��̭Uɹ���>�w� ��#�zNA>'�|����5KY�+��W�m�8�=�*	�� �� Vj���a"���(Vi�+�>����輓�~ӧ�Yv��$��uޱ�k��ip���o����֧���&mɱ柧>k��>����-��@{�S�׭���b�k��ɥ��knx�eLk��� &�W_�������u���?C#���e�Y۪��Rk _�gy	���S��蠾����Z�s�X߻����������������C�ER�&�w棾;uTY���C�p�ZJ���X�)�:����~zu�G��X��X���Q|���s,K�ß[?��v�[9g8�m����_בm��m�i���,����e���{F=|����z�6<l=�u�ߵ�������u���Y�I�\Z]{�oz�	 �:���k�/{����v��:V1'3j[� Ϲh�<��Pn�wE���1�u��t������<��垰�*�/Vfjd�T� �a������!� oG���w����f�Y��#�&a�Q>��ˏ�Si����8��8�G!�ᆫ���K�O~���\KJ��0}\�>K���m������F:�]�#�z�^��Ⱥ>W��m��{��٥�E{`�{x�ȡ�pY�8����)H_\[�"��? �cp���}���eoy�%����5T� 3εm9wg}x����o��>�QuM���O�כ��/��-���Be�v��t����7�����W{���qc�cU�g��V�?��7]�� 8*�Qn��ۮ|���~}�q��dnN0������.?x�ֱ��kz���4p��_�X���p��^(GہI�S�4�r�3q���H�I��h��-���9������n �1� �s�U/\zŻ>�3p����݂G9��׎�E��DZ�p�怾���-ռ�Y,o�͗Ķ	�G���]��Joxڸv^?F����v�t/��+
 �q� ���W�{}8��?����pۥB�=F����@�Gf�جѣ�z�y}��=+������4��{��c3u�H��v��9��f?���3�G���=��3�g��/��0 �����/{����'��V��	�~T��j�mR�����v�=�iEϑsE�9W�]���z�v�0������F_V��D�����O����y��W���/� �0��>�����_���?������v)����X��x�S���w�^�lN˻N�:�J���4ؽ��O���P˗�;Ho�(��`|G�=����>�������[.�Y �@&|��^u�o��s���?��.���a���k��j�C�z��˝����'2W��u}�b5/���-�\����#6����>���#蟝�7�pr
&��~�C�^�f �4@f���+������_[�&R�
Nؑ#�&ĺ�?�Zj�v۾��ל���˞ښ���j�h�\FڳH�����4��a�/w���?�ݎe=�YW~�j��Ri���]�1j p�t ���+_�oW^��]���~��x��z�+�db��ӣ���mr8�u+U9�7�ӷE}_���]��v��f/�F/��a���F7n&h*��o��n������]}Ū  N� s����� �=�kn���=�?��[��Std�Lr��ǣ�N�o���u:�ki�ϥ�^/y2_��\)���K�������&Qᡬu�������ޛ4E��������Z_��k�� �a:����\��������_{�?���v;9FS7��̭�2tTY�����mu�����B��S�M���}��>���9B�=V��~3���"�~��� 2�͛�����$N.*���O�y�U �:�L����/z�{>w�W[���'�[^({\�o�#�F;2֕2�T�殯o?;�w+�U����0�K�+��+��^��o�4䳾Ӽ^>����"����hx��#���]��8{~4�1���ѩ[}�ɕ�����}R  ��@�y��e7���]����-g�s�ygm�d:�L����cݴ��'J���Az"Gy9���i�ӛ��[<��m����N��>JN�z���=<�]�?�����������ֱ�>m���w'`v�����I&�	!KX* ���j�Z�\�Jݪr+�,"Q�6�9g&��a��L�9�<�jY�����E�׺[[����[Y�,Yg;s���4�FdI`�y�9�����7	��?���_sh�7�F<in�V��C=�'�<~,kFx�]��o~�9o~��&��D��B�*�-���]��~�����I `F	t�-\�bE�>�S����m?a�sN8��E�S?@�2�H��z�?�f$��s��4�������Ծ�?�ɵg� 8 :�V�}�ك��Ư<����g��������Un�']�!Oá���g�n�ݏ�=�� �@���#����<_xۥ��u�1�|�)G/�]�A��g[�vf� OK�F��=�~��?��W���v (����,k�k��s>p��_~h��_>�����쫕=��G"]�w��oSw�zz憩���=|���[�� �� Ё�v��s.}O��o��w�I����^��GB�������w|�2��(����y;^�����F ��@��p��;�p�Y�\���G<��pDf��<�T��:\o}]y=?i���o����b �`�@Ǹ��V���͛����/����`�zhO�M��/��G�[��sxq��c����K��� ���@G�r��Ⱘ���>sג�o��ˊuъ�6�G<�{G��G�c�����}�< 0�:Бn��������s��ŷ<뤓������/Q�X���=oe�^���<K۷߳�����A�������p��?p�Uw.<���?kY��XP*b��ѱ�dW�g:���s���ٞ�;���Sz��O����/ R!Ё�w��s�{�~l�׿���N|�3�u�<���xt�
aZQs̣�������\����1 ��}�����q8�̵-���K�{��=�s��6�󱩓�?\�n��� $I�����r���W���՜�N���r�a��R)�ºB��0w�m�,�_����o $K�<ʕ+VL��e�^w��������O\t��"h9ˊ[8�w��W_|�W �� ��#�Ͻ5K����w.8�}�}�qs��vu y��D���;>r�ڳW Z�@x׎���o�<�����#O|���]���@�z�t�Ĺ۾�lQ���<��� -F��=���꿯����r�-�y�I'�0�["̲b���Ň�ZZ�v��#� hI`?|h��w��w��ᴯ��{���OX|��ӁY����Q�m[NX0u�GW��W��&�����>�/���K�z�=?\\}�3N�_�?G�͢|�؉�v^r�%�W mA�<W_|����G���_p���'3gA����/LL��7��O]|�9_ ��0�>���y�����s��Ɠ�;�k^OQ�3fw�����%�.}ˇV�i" �v:�ɲF�C���?���a��3N^���oN�P���0^_>w�[t��9@{� 3lO����o<�_�s�ǲC�x�P�W_>V_޻kO��Y�t �p��t���q8��͛W���{?ӽp�i'/?R�O�?�O-����M�u�+�� ����4o}��ˮ���eo=��es���L������;>���ۄ9@g� ɞ[��kg]z�%Y���sT���@�ZT�u��Y���w��� J�̂�.>�J���[���۾Y82,Zv\8ni(����7²�m�.�|�5��ݯK>; ��:�,ZX����w���4�,9>�xԒХԡ-��z��m?8b���W��ܯ ؋@H@oq:<#���?��-�B8ty8��¼�b Z_�������c�����~ �1t���<_| �m���7gYX���p���5uh-���f[��;�����]��r ��@H���x��a�;ÿ���-<&,_�8��vUR6/L֏���/�u7�u��y_���K� ��t��5o_�	���	wo��{��#�:&d�S�dB+�x訹��c��U7�~�t ��$�ZD�Ǐ��B�����?j,
��a[�5m0[v_-��q���>��� x:@��M����������ug�c�0
8��C�qd������Ͼس� ����v������_	?	�LΏ�>/��~H���̘�o�;�1w�����}χ�v��O�=' �L� m������@�cl^������|apy�_�f�Ǝ�3��%}�=-��� @�u�zxf����ƃ�{��;&�����ǿ�ǖſ�v�޽�����5׌���  �@hs�S�9}�>&����]=�]���#�<cc���������֜��  �@�t�9a<�2�yl����c���Ï����:�+�����mK�ƾ�p^�Е��v[ �Y&�:Ts'�S�m�}Lg�p���p�Xo�Q�?ƻ�h?��חf�<�wꖅs��h�{ $�w` �b>���}����L�۽�܏&煇���c.��zvߺ^�5��k��K�柞�wX�C+�6  Q��RȲ�xu[�Xx~x L��*����v��M����� ����K�;\�5v�9S_����y��!�xB=���z8��y������p�xo�gr^����0�̖��vl_�3�O�t����Ϲ) @�� 업ŉ�p�D�����}{#��DO�wj~�/ゝhn����ᰞ��b���O:����_; �t �������X:��3|ض;ط�`�obn<z��ag�rϰ�d��Wc�kW8�g<1g,����ݥRim �6"��1�`?4���_��k��Ĝp�T���ީ��{��Y!�(s�FXT�w���{&b�����% @�� Ps�z8nn��ټ���\.�=��ͯ�5U<sk������e[C����(�;ȜB)����aI<�ca,�E @'� tW^��q��#��o�������ɼ�5;�S�׻��ј3o,��ʃ��[Y���DXP����#ė�L����  �4����r�/5,�v��.���z��[��9~}�t׉�݋v�=�q��3�ZSҼ��/��Cb�/,N�E�Saaw=,��CW�� ��� $��w��Gq��=�:k���=݅��Yo��X#;5�����˻�L��E�~`t�e���м>���1��1�'C6�,  O�@��\7r��q�z��S��y��{�y��dx�����'B�1�ӅE�yW�x�8g2�[��=��X��|�k̚�W���]�q>�{�?g� ��� ����_�3��xL+.���;'^Zo��M��gL���Syq�d#�?��z롻g"/vM���tV(��k⚯)���a=�P��t�Bo���#��Kzo����w;��l� t����84������[{����P��g���؉ɩc�y8�>�L�aa#����=�Ѩ�L�����{Yw�>=ݝ����TW�
�������Bs̳�Ѝ<�P���'�Ph4�wnz*ϊ��BV�y}:���#�B}��X�^��=���Ү���1������b�
]y}�&m @k� �.?��cq�}ϑ�6�h4^�3�� �R:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @: �r�<?4 @�� @�ɲlQ�R�_.�w h hI�B��8|# @�� @Kj4��6"����e���pI �6!��V��j���R���  m@� -+��8t ڂ@ ZV�e��š��o hq Z\�^��B�P�K/l����1��  -L�@���>���:U��j�3�� Z�@��`���������<�bÆ_\�jս Z�@��e˖񾾾<�B��_�����b���[�hU Z���H�Z�>������q.��M Z�@�6������{l����F�	t h1��óB���Н����������? @� ������~T�^����ᗍ���
 �": �����s{���E���7�H}��  -@�@�q~{��N��~u\����@+� ����n�����3���q\  q ���5k�T*?̲��O�krq��{K��G $L�@����8;�3�<�P�V�����M %��MdY�� �S\�b���T�Z�)�J� � � ��x4�Q��f��y~]�R)��� $F�@�(�J?�V�ߎ��ӞH��V�e� H�@�6���1B��s���1҃H % ��'���z�Jz�R)���k $@�@������'�|V���juq�T� �e �L��W�}�)�C%F�����5�4 0K: ��y��}jlllC�;����jG�722R 0: ��/�pG�R��������h�ƍg�\�r" �A&����j��x{�N���;SSS������� D �ЪU�n�V������ׯONN~itt������	 p�t hS���(
�ݳ�!.�/��X�~�i����	 pt hSCCCߪT*7��OŲB��j���R�ts �L�@˲�� П��x�Y��sc�" �$���Ũ�5����OUO��7T*�g���K   �\�^oWW�+�t^�)���p�Z=���E4 `�	t hs�W��+�e5N���s�m�v�ƍ��5l �4�  ˲u�����������SSS_]�n�i�W��; �� ��*�J9No
̄�tuu}-�����w � � "��W������	�eY�����-�J_ �4	t �,+�<����f¡q=��R����  �� �T*��Z����̈,���H�t�V�````s ��H�@����g1�o��33"Fz1F�G�.��: �S ����ߛ����8=60��*�Jߎ;~odd� `?t �@]t�õZ�͍F�+�[�3&���������ό�^ ��: t����oT*�R�~(0�~7Fz!F�[E: �J�@+�˛�������ӛ��y��3V�X1 �It �py��;˲���3�M۷o�ݸq�W�\9 �	t �p�ryg�Z}c���P_�i�MMM�#��"�'"������R��!No�GO`��frr�����7z&��#������b��'˲�3.��k�������v�`�t �?�H�x��gǘ\�qq]����?���;�< �� ��;v�cD�����j��q�( �^: �S��_W*��fYvK<}Q�@xo�Z�R*��0 � �͝�k��o�y��x�s�ვJ���� : �8}e�X�Z<]86�_������� :�@ ����=1 _^(��~D`FeYV��'+��o��� t4� <�����U��W�y���3m^\�?����_t�E� �X xR�R�ۣ����X,�u<=40ӎ���y�e��ʚ5k
 t$� 쓡��o�_���B�ps<�̨,�N����Ӎ7�b�ʕ��#��}688��j���8�|��K'''���Y��#���R*�n]�~�oeY��x�fT\ӷW*��/�� t� ��������<�?'��+FGGo�j �ct �))��_j�,Fz�J�������](n�V��/�J? t� <e1��!F��b�!F�����yx\���ddddW ��	t �ii���V��f�Ѹ���������Ϣ� h{ x�n��=�I?:0�ΪT*_-�� �5� ̈����!��,˚�I?)0c�nZ�~�?�S �m	t `Ɣ��;k�ڋ�Fsw�f�ܸ��~���ڗ@ f������J�qzS<~+0#b�����E�� hK �q�ry����������a���Lyg�Z�r�T�D ��t ��������?���20#�<������npp�{��"��&Fz#�V�?�ayy�,��%\�n���_=��ӧ mC� \�T�X�����|U��?���y��c- �6�	 �W*����3Y����nذ��V��= �: pД����j����������S�eٜF�q��͛_�bŊ� @�� �A500�w6l���O�<��}��r�0 ��: p�5o�}q�XlF�sOY��kk���n �4� ̊���{6m�����㟎������������_�g�| Z�@ fͅ^���o|�]wݵ)��+�T=������ -K� �jϻ��]�V�ջҟ��l�*��g��� -I� I��]�ͫ�=��}Q\��8=' В: ��=�J�;N�g΅��uV�V�>��� Z�@ �R.���aÆ�4������Y��<�7m޼��ލ�z: ���k�j�ڋ��J���_���[�n� �W Z�@ �400�7�tjj�x���>+
���˯�袋 �� $k�ʕۆ��O���۔eي��Z\����q( �2: �����z�U�T~�˼�m��e���f.��w Z�@ ZB����5_��;�d����qf �%t �e�H�n�����@��x�xBq���|hh�[��	t ��~�V��,���k��H�X,^�W �'���300���/��W���-Y�x"��V�/.�J� �&���t�E�K�����gW����_ H�@ ZV��;֯_��1�o���	<��>�]�V�W*�� H�@ Z����}�]vٯwuu�e�Ӟ��o
 $K� -o͚5�����P(4#�%����6l8uժU� �$���044�=F��c�>���V���~_� $I� m��7n����ɛ����⚼yݺu��W��; �� ���+Wn��������q��[W�X<?�k �� @�Y�z��鯌1��,�^�ۻ6n����+WN �"����'�_���uK<}~`�,˖NMM5ws�D  ) h[�H��j�������qA� �� @[xp�ƍ�����Z�e�
4�hÆ��jժ $C� mo�ʕ[j��iy��m<=,���ϋ�@H�@ :������_���B�+�����,;}xx��FFF& I� @���Z���F��W1P��vh__�+��� @: �Q��R���c��B�lo  �8�r��1�eY�G��ů�u�֭;���} `�	t �#�H�p�Z=!NB�[,_�� �N� k������'��i�s�%t�$t �c���4FGG�R,o��?:P�e��iӦ�/�pG `V	t ��m�T*���o�X]:O����o���:� t�r���j���8��Й;��V� �N� D�R��J�ri�eá�į�U�Y'� �رc����^�����,=ihh�� �F� ���4n�ƍgNMM}'�.$˲�m�`	t ���\�rK�Z=;��c�f�C
�_���Y#� �T*�R�T>����� �J� <�;v����,NO
 ˲#׭[w��ի� �
� �FFFv�_��1\��)��
���A��� �8��Z�^��`O��I `Vt �'�e�`��xm��6�9t��%� �������j����c��eY���Y#� �ı�{͝w޹*�)��Z��5�P" p�	t �'q��OW*�K��3���y�<`t �}P*�n��jk�����eYvB� 8�: �>��W*�q�>��=W�� `����899Yk��:�,�  �h�ʕ�J�8-�6�
:���  �!˲O�6���-
 �
� ��S����#B{� � `?47��V�_��3B{� �D� �<��>�z[z��� �B�̒���vuu��7���P(�s��pOh_����0KV�^�5�
@�ɲ�m=~ms6o�ܽbŊ� �A%� �S�T�5���y7m�Է}�����������K� ��/�p���y֬Y 8�:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $���╈�B�    IEND�B`�PK
     t$v[���z"  "  /   images/d4c851cf-9fb5-43cd-809f-e1699313b4d2.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  �IDATx��	��yǿ���sg�ҮVZI�@Q"�����lC�rRA)!l��ep�XX!�2C�p�#�X�P��!�х�՞�;G��_��gFI�����U�_�v�{f{z��}�{�^�
uEJu SH�T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu SH�4,�|页Я4�!m��%c ����b�����=Z��vx��0�Y �<��J�N�A?o�џ@(͸�	@�0.L��r�]/�4����F�nb<\��h��ᅛ��pP�\� L5��3}<�7��?-�<�S�:F�[�X(����A�t����|�|M��;s-�i0{�vH�<�x�IeE
�e�6�xwl�4���6�I��<���T������$����֊�g	`��<�	�),O���L���>E0x��� ����,}�Yk؇��X����|�gʅP�Jni0���|��1� ���tZ�����>�"u�̪�p�ҏ�Z���j�%k�-�1 Kxi�u0��yؒ�_Ja���C9�@$�3�:q��mɺn{���;
c.0ֆ`�O��ϫR��Al{/v\��x�%��5Ky��#���Ϸ=���+�%�
5{C��Iyr�nP�|��.�^�a;E�wU�<<�%S��L춓�-oMq6��}�}�4��j�ek�D���Xa䢊���(��%E��Z��پ��)J&����㉓�uc�g��I���{L���G0��:cګ�ձpŲ������j�2�~��F�'�T��8 '4jڬ	�8�p{m�e�AL\���~��m�9cL,6:�(BJ�`p~��d�5m�om5M� �� e�"���y�WY��8��O�Z�&@�X�|Lk��� �n�1v[��3Zc�n���q%k	+ƅ�A!+���8�{]��C?�-7T���N�%5�_��Pp����m���~L ����J*��Ё����MI �N��j���B9�"�8sl,�Ⲽ�r��ML&^�(��5}_�>>A��]�Ӳ�
��3%�L���#u����C������1���u�	7����G5�@��Ko�w�]��ʸ�}
���͆q��{�Xj�)�+T�/o��MWJv�HO/�u��yފ����i���۽�:>�L�
eax�s�i��/cj�����B2��~�����V��qW�R�椪Κ�W��)�qV�@1�̋��=/�/$m�c���P�� ���6]:/c\�q�����R�@�ˮc1�/ߊ-�Z(�3�������'K��?0�?��-��5����|gA�����L��-�$�R��)�`4������ʾ}v�a�����(�@O�F�q"��k[�]��h#�P���\�{�=�p��AiL
��Oi1�S�DAw��˶W}fY��0YUd%�ti�3П�w�C���[N�Z(4 _��5�d
<��r~��!H� F%�%�����~�����,3p[�����L����FB��blk��-i��Fn-�P�]e>�fC���a�����N�����A���Z)4 IY�~䀵K)LP���h����A/�B������C�A":a$S�P#�$˰W�T`����9�
���9�^��>YG�8�.k¾Q#>�@�F?OC��i(�orG�Z�YW�ފ� !���-�N#%w�j�Ѐ8L�B^�iP��0��OE4�>�1ޣ.[�J1�B��L2�H��V���.	{[l�
�"k��C�,vtU�K�����K��I ���ˣ�e���s��z)d1��:���;��a ]�6�|��s��-�,0U��:�b�g�q�("1�m�u �cY13�5�\/���M��4-��3E�8W���@ �X �/�mL�J�#�Vu�W�ˌ�.�I��׀�"�WD���m�S4�H�0�X��'W��s=#+�eEH v�
a(F܌e��(`���V>a���n�� G*��uÎ5"�}�K���jF��`X� Cӝx�����瘆��l�|w�� @R�gm��N1Rur=�`�i��yp;~��-����y��2�`��9�ˢ�3䙔�	�]�2��T��3�0���N�W�I�g6b��w��1����H)�
�1_����u`p�.���%B�e�{cv��ݕ���[ST��3�?��a���.��R�PW\P41Ȅ*&�jaZeUƫ��t�%�h�$}�#�;O�]�<�H����|�`ڇ[��,xV�{+������͢JST]��%U31P$?Ps�>G8�kZ�AGѳ2hE	�
���P���t�@A"��ܿz��֍���[���ᘦ�x&~� � �+Y�P���޽/���1���)�B�� ڄ�X|�X����������E7AX
�'bŘA֑�j�g,�q�c��OЪ^G�r����7���iA�;#>T �� �:T������"(�!��h��7Yl��N�2�E�GK�Y���s��;mP�I���2/׶v�	��-|�,���s�/���:��H��w��qM���#%�'��T&��_�)s<P^_�ng@|��!������A���E���do�lN/@η�߆tj����;�<t���1���J�g+-�ڑ8Z�]��Zh@<ǆ��3@���5�;��s�n���;ت�#�dR�
�7K�M�A?�ǳ+�C��!,������8��G[���X���*�̟:���8%�7��K4e{便C呮Ύh̄j�sY��btϱ0ߧ�����x�����}�o�5��[�q����G����� 0]�'k�#�Gd�m�h!�4�&�h^���z���s���c�����	F�
�+l,��	�uK�L=��G�@vmZ	�b�\_2��E�M���qt�ze�/�%�()h�;C;�pǲ�4i�*�g�`dL���|��*���T9����0�T���a)\ e��o=�MO۪JK=k7��9ƌ|og�&�Ub�B9ȕ�_�GB�Nt]00��$t�>��a+ĄR`,Q����P��\OG�^��1������Ԙ�k�����B��*��eaDZ����ʍ����Z�k�QmM7���P��\[��v5�7�a�u�A�r�H<Y����K�,��cƀR�)���C�9��1����bq�)ji�ա����++�=r4U3�Msٔ/ u}��5+�d���B�!���'2��u��76�٧��I-i��"����D0�!)�<�uC���μ@��̌�ؾ�#$1��8�b�v�JxN�pGV�^�Ea�����r��	ZȗlB�!t���~��-5��;oj3���S��v�l��s��b���% =g��ؚu��(�಼'���Y倻�Qn�\���3��Z[��Ԥ�tPyxo�-Y�`J)��}�
�^�vĠ�O��|	�Th@t& S��d�"��%ʭ��i-줱X�1��۠�1gLh�F&���I(8>B�S�E_�5}/�Ha)=$�%�����
��P4�h�+0*��Ƙ�H�z�6���[��RZ���O���~��W��D����BB�KsV{��a�܎���O�ЈY��3Ʊ^��w7wó����p¨L�����֖V5�@��}��K�D�₦0N�Tyil�r�lX���:�=k��5�M��k�ܻҖ�6Wr8Q���orCE��5"���a��\:kƷ�ٷ�v��`K�Qg�Ǡ1"e�YG��9Ț����{[z �)�!��2	�%�pT����X�Eۃ��B��`��B�Ɋ�������W�q=�f�_��� �	Z~q�W�
Ȓo� �/|�̦�_�	7^z撞lnU&��wl����+��9=W�R%�<�ߕw�#���vO�����i�Al@+Qh�-a�/XC�We��;O����?nn��s��=�C�j���;�<޾�7p畧���~���<v���\ws�п�s}":����R���Q��W�c���|mӬ��Y�D����kPK�d�܏��"��}&�p�z����K>����IZϯ��x.�r�gAK�Q�I�@�c��1�d}c���;E����5�.�^5�J������y�
��>����ݻ:L��21�b�`�������A�0���XV�g�0�v�z��Ǚ�U��R��izz�s�����S�'[�w�p���؃�j0�z�fB�V���!'4�`e�_َ��4�~]�t�':YRZqGLp��A���Ն&ն����ͦv8qp1�\�� ��q0&���߹>���`�9��T�3o�&2���_í��.��O�ͅ�'�����j�k�KF�l�l���l��\/���__e~� ?�3A۰���kZϡ*�@�E����Y�.�pc0f�3��u+�Zf:��d7GK
<M�򫢎�
����a8(�@������w=��~�Ec��Qа��Au ���\Y�ݧLn��u/@$|��V��9��ic8@9^�Э�iި^��,�IQ�2�kM�� ^��]����ǡ�ˠ�A;��i0o�<���=���}�a��ˁ&���|�
���E{ �E+?XYЎ�,/����b��h#��k��?~i,�����H�����b��/�ȨA�@HT�UP�CiA��-²��5��� �
�r�JV@�|��1P�_�e&�\���B�
��K���q��~��Ҭ{��*��+ �}��j,�byJ�Q��w^� {.\w�q�Z��>P�c�"�Wa�E)�\,OD�J�d�a�C^۾�5X��Ox+Y�E-U���]��~�&w8���n�1�����gbq��W���6��"���)ݿ��i��	;�V(x|Z}��U9>?�cEH��>֕��\"�H 9�}��5<r EH]{T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu ��=P��&q    IEND�B`�PK
     t$v[�e�e�  �  /   images/3d0a314b-f708-4b2c-819f-35c414b123ec.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx���	���}����tH��$s�F��`.� �v�aBf'�O��ēd���`q��$��Ɍ3;;�M2�0�F�@�!��!�9BWKBg�������[���V���<�t!d�<���[����l    �8�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   � ��c����Je^�V�ӨՎ�4�����T�ޓN����I�j�S�F����T�֛�Z��ߓK�7��r#�*'�k��p�K!��6����!�5�H5��S�dv�����J��յ��5k� h �Fޙr��|�~b�RY��V��V*s2���T���fh�����K/����sJ�L�X�fG>2��J.����n)�ӯ׳ٗ�s漺�O�� ��	t :ֳ7��[ڿ��B�zN�Z=&W��k~����{饾�oI�ȥ��B�s.�Ri����E?�6m�|��C�|~o9�����R:�������G�ԉ_�B)  G�@�#<�|�	S��s2��ݥ�)�Ri~����
�z&��z=���<zBX�#o�������W*�����\������N?����7� 0a: m��U�Nɕ�Ww����/4?�޼��nE�V3�������3����/�x���7.�x`,��B���t��K���  ��@K[��O��;w~�06vy��؇zFFNȽ�ڔ����V�z�����~e����=wd����������7uw?|��5�  ���ʧ?]|��k�1~y��ة]O>yt�V��]�\�\.�9y��d����fK�]r�c����r_�����`��N��o\{��Ӫ��=�×�=��IS��hq���I��'%�Y!|��c.��������e�k.��W p�: �y��??::�dR���gt���M��j4�OT�tɶ�du=y��S[�;o�p_�����{�;�.���� Da�7����w㤑�kz^y�t���m�@+zk���k���֭���|�������}�-# ��#fݒ%��J�>>ytt��_<��G9������}�$�����f�%�l�2宝���X��b �@`�={㍽�={�?�;v�e�[�i�7����<�d��y��˞�鹧�����֬) �P�qw[���0ix����?�J9?��VS��]�<j�쯿r���4c��E��� ��t ���˗�0�R��i7.ΕJ�&�J��Oݳ�����~w�ԩ_ߗ��ɥk�n �: ����򱱏Oڿ���[����t�w)W,N�],^?+����K/�ށ�So9�C�J��� ڔ@�xbժ{GG�ɴ���J���T��y��?ع�7^���
�岻�� ��t ޗ�+V��>8����^;����*g���iɪ��t��^v�3{�L�O���_3 @�� �k�6�����h����[��M�L�z=��`���ƅn�3u������w Z�@��=��?�wh�fn���p�#�gx���㦭{����.^|gc֬�x�-��W��$����q���*?3mÆ�ɤ� �)��Ξ;:�����7�x�U�N����c{ �"�xG�\��ģ��~{���%ۊD.S.��ܹse}Ϟ��P�oߤI�w�w� �t ~��Wϟ28����L��~V�r��j���Mߵk�����o�N���B��y��=�������}v�o,M'@�K����v-n~]_��UWݿ���sW�y�  � �V��1wt��gnذ�� m&���l}��o�5/\s�ݛ���[v�}C ""�:س7�؛۹���6]+���r�{����O��=�d�-/M����׬� ��@�PO/]��_~���ccSt�\��7g۶_��ۻ��e���u� �� �ѥK�������l�z\��522縑��{�%�|j�QG}���o. �"�:D2 n��=�?}۶�B��
����{��/]qŷ��:���z��  L���W>�����/����w�~�z=3}׮�'>��ŋ������|: I����˗��>�Ŀ�Z,N�!ɖ�}s>5upp��U�~}ѝw> `t�6���ճg����Ӷl��a;;�'�##8f�����+�x�4oޯ�}�-# Ƒ@h3�t�9�7�j2�����^O�صkqyh�ѧ�/���s�W ���&Y�jἽ{��o��3pX�K���m���W.��cCs��+C� ��5n�)���O~f֦M��T�]�q��{�\4���o<�t��s��- �a$�Z�c+W����_��9CC�`Bd���l���.�l����i�wl pt�������͛?�qu�Sj֬L������k�;j�Z5��L޻������^���<wݺ�
 �>	t����fN��S6o>7��0:Z�_tQWH�R�^o4����|���ju`��ؽ����d��c�n��KW\q�L�_,~���x�:@y|ٲ��6l������ �Icd�����LɄt:��>=�m>��'���o(��P��7o�V7n�&�7�C����v]������U���{�x�:@x��?�޷��3�n�.�לq����@;������|�?���8p�Vk���b��zSatt�����s�\s�^xS�曽���"�"���ۺ���>:�8�o�V���?�ߛ�4)�=��QH���w�U7l�T_y�Ҍ����t����}�Ͽ���|k��z�=�� �	t��%���l��+�Z-`�����N��s�f����K�{��*�X���r��gO��z���	�ſ~rŊ����k� p:@���S���d�-�4lig���7FG멞�����$���睗	��U߽�V{��r��;re=W.��e�~�k�r�׾��  ?�@���Wϟ���e���B{�H�;��i���HϜ�i>�s\Еl��|���ꫯVB��9_��zz���׿z�e�=��Y3 �t��<�bŕ�l��Rir�	���/Xp����T*=~��|�?�Fm��J���M���r}۔�{?�56���?��_<��۟ �6:@$�[��Wfo��ϓ!S���֭�����*RٓO�'�ܞ=���ϗ*/�P	�jۗzat��y��~���K?���{� ��xp�={㍽}[����[�p��|�֨T�\nB��g���/��'w�E��K/�+�ח����L��u̶m������Щ]�YW���	t�#���L۸��CC�8����ع���?BoH��ܙgrg��OΪ��}�\{�J�no4R�v��Ć�:iݒ%?���� �p�<�r���7m��\�8=@$�C��@���Ϊw5�]�j���;8T�MC}���g�V����+n�t�����'���Ǘ-[~�֭�W�\���{��0KϚ�),[֛�S�|�;����_NV��M�����V���+~��k�
 t4�0��]����l��k���d�P�7B:=!����z��{�\PHΨW_x�ܨ�B;ɗJSl��W�W��7�֮�3 б�8�@�]s���ٺ����(�~B�ܨ��]KϞ�k�ԤI��G?ړ[��P~��R�����=w��-��;�����O���_�v�B>�{��O۾�� ��m�]��@�W��=�P~≱��/WB�H�뙣�o��/^u��S���_ t�(������Sz�o�J���	Z@2I=�uV!D,5}z��tio�3*�G�������Fj�Ν+_��)']z���6��"���߬\9u����CC��Z�-����O~2[}�����ط�-�v��]�ox��5/���p��5� @G� ���իg�߱���������H�18XKM��	� �Je.�g�;.Wy��R����a�ܔ�{�
a�+����'~�� @�� ���eˎ=f`����QZP2�=�*���L*w�]�Nȕ~�X}����	�N&��{ցg���go��cg�r�H ��	t���[˗/8n��/7�|V�u��)��CJM��)\w]_�7*�*6��Zz������ү�~��V}��;�� h[�0z���N�?0���^� -�>0���ɖ����|���c��|�����{8�F�GW����w��f �-	t����+>|��m�+�����޽���h=�ӓ-,�˥�_ܝ=��|�k_���ٲ��3<|�����z����Y�- �v:�a���U��ݶ�ϲ�6�܇�]�����3fd�����Շ�u���=z��>�߿��5kv ڊ@x��X���9[�~)[*M�F�۷W���.�"�9������7�l�JO�O6��|����.Z�fo �mt���[+V3o`��\�4%t�Tww�Q,6m��B����33]��d_r6���S�Po�r���s�<{�י��>:�{��s~������d����rg�](�}�H��7�2��;�y�F��H�q�v���_xaw��>v｣�Z��{���7޸����^���D:@� ���n�9k��;�FF����s��.�NM�t�<ra�Ҟ���<���z=4v��o�m�?&=o^���þ���X{�Jh1���'|0�/������׬) Z�@x����O��i���##�B�K�<������@+�]+V�6#=�J������@-�Ɓ~Pww���Sy��r��(�� �I���׳��y[�?�~͚�����]���{g|����cC�˞tR�Ќ�$���罹O�t7��x�#�x��CS߼�-j�t�����}�T*w晅��ٙ�u�FCC-�E=eϞ��J�Y��? �,�p�7ݔ����y��gK����W^ٓ]��g����>:��䒮�7�9hK��[���r���K�OM��	m,=gN���~�o���Zj���ݻ/�k����}���$��K�>�'3��]�X�Sr��/�I
��Z��Ї��{�ԫ����m*�V~�R��̛�͞yf>{�	�d�ZhG����{���O��F��8jǎ��.]��{�����#��w/�쌁�e�]5���teO;����W\���'����V�&��7��ʝqF>{��l+�T*�]�Y�ҥ��/�r�%*��h����'W�x���k� ���3<�t�����Ц2��e
K���&O~�[�3�Taٲ�◾4�jgwyo����+��ח2'��ϟ{n!�K�Lv��|���̌�u�H�|m�����۶}����.�瞧 -C����Xq�1۶���|��M*r�ߕ?��� ���Iw]{mo1��^���j#�_2�<9�P}��r��=�hQ!={v[��HϘ��ᆾ�=����.�L��ưo�ك˖��rݺM���V?@�GV�Z�`۶���V�Ӷ��S�%Kz��{X��JϚ�I�H/�];�J�v9������R���j%���r���f؆6�J�b[�����C�V�����p߾�z����}�-#��	t����u>k˖�j����LfΜLa��ԤI�Oمs�f�U��m��;Q��H�n�PɞrJ>ᅅ��Z�p�Q����N��W�%��{����n�t�m���ݑ?��c���^����=22/���9�
�\�5�ӷ�m�={jɊj�3%������/��g�]H�S���֟����Ԕ)����z���'����]]����3��	t���#������CIe2!�U��SN����͈)\sMOchh��c�U���Q�<�t���˕��w�N>9�|}��;�|�Cyݺ���1v3w�X��O��v�_ �%����˖]?g��O�6���I�/��|��=?�=��������;��p�|����^�毸��Χ'�9���}'������ڶ�X������� @�:�[�^��y[����_������W��M���{����]�?�+_n�UF�_m۶���x {�y]�E�
�}�b�����v}�}c_��p�oDe��¼;�t}�Ջ֬ DG�4={㍽�6l��L���Dr�Ua��d%�H~�s�����)�w�h��ֶ�o{,&׽xqwj֬�~=r��f���~�H�S D�0::{ڮ]�|�� @tZ�"��ҷm۟��P�ܹ����~��!{�����ݵ���� oi4�&Fo�u8��r���ʫ�i�2=�_�W������`ԑ>iϞ=w�5�s�׾�� @T:��x�oM� ��t:�/��;w���ݞ�aP߷�^{�5���;�z(?�D��ys��dIOjʔ�=���<9���O�׬iE�sv����W�xn�ڵw �!Ё��|�z͜-[~!����ڗ-��.\�1J&�/^�ӌ��Ʈ]��#j۷�F����WvgO<1ί�C�������WLΤ��o����۷�ރ˖=s�u� Q�@����+�6_��A�^o����S]�^ۓ>��\�Xr-U�u���!�S��h�R��n�h}`������V��G�������pĈ�����㇆���M7-N�|s��'@'�@��������C�Kuw�����7�Z@��ص|yO�_I�7Ï�<�l�鵃7L�|Dn x�F�'>�;��/G=8�op������j>u -�b�p{f��_��u������%+u����[j@z��\rV���C� o��曵⭷(,_ޛ�?�%_���z��^3񎑣v��_֯Z�Т;�|$ pD��<���K��8gǎ_-�+t�:T+d�ػ����xIԖ�c8����N�n��H�`�Z������r9�HO���}�x��/?��[F G�@:�m�����K�Z�
-�Ӣ�[2� 9g|p���M� o#�3�����޽��%�t%�C�Iϙ�M��$o6$�>1*���*l���ͧ� 8b:�QNٿ��{���v0���{���e2��%KzFo�-��q���.���z���zZqx\�M?�|yoi��hg/�x�ͫ�����Ϲ��� G�@:ƣK�^q��@hao���%��C���Nw�X�[lFz2�;�;�|������Hr.=� �����G?�]~��Xg/���#���G/Z�f[ `�	t�#��ս�������W��zzRݫV��T�&9�[X���t�]#&���$�!J_��pr�;ys'���g���*�חB���r߬;����k N�a~����bqFhQ�R����ZmZ���=��\㢋�ʏ<2২��Q����dBz����"=��]I�W_}�"4e��3��.ι��� �Ph{�W��d�ƍKC�Juu��>���d�9��ܹ�{�Ԓ��~���ݵ�d%�������T*��暞���pm��(���y���<����k�� L���dj���[��U���2�еbEOz֬���ߵ$\����>88\�2\�G}Ϟ��HOv����T��r�T��z�_��p3ԣ;ב)�{�����O. 0a:��N޿�s����C+J�B~ٲ������I2�T!w�Í��Dz�;Fz>���;����'ׯ������h������gM `Bt�m=~�u��޼��Т�_ޝ]�0:P�����b�V���ص�6v�]#�d�{�MwOϜ�)\uUwiݺ��F����k�o<{��ξ喑 ���@�:j������Zr�9����YgBK������t｣�R��$��J��3����j��gO<1_߾�Vy��&����;����_ Ɲ@�ҳK��Z�m'��|���]pAW�`�$C��O<]���W�=��ha��d�Ah!�K.���U�m�Z���k��G�.���{�}( 0�:�v_�z�Qo��OB�uT&��-�)y�������&��3U_z���4i,��ݡ�$��,�)�z���H\[F����}�~���K�_���F�q$Ё�3m��?�T����ח.\{mo2�9�wޚ�^ۻw89k�g�<�T)=uj:{�i-uL$�|X��w��ۇ�Qb�=22嵐�_i>�| `�t��<�bŅӶl�(��l6սreo�=��7-�������/h��Ƶ�H��=TLO��Iϛ�2�u����R#3kV&���g�����^���qǛ�q�2?� ż}�~7َZL��+�;���(5yr���c_��p�]���kd��G�o�aR�bR�7�����wגG�3$	�F���O�r�g����6��� ���@���ҥ��o����;�B�S:�:�w+=wn6w�U=����J*�oi�ڑ���Kv��O�Vk4�7߬%C��;v��V�>pƞ=W=�bŇ.Z��;��N�m����6mj�k�2��e��́C����h�N�WR�$�ˏ<R�_~y�x�Y����޽�Z�Ɋ��=���v|��9CC�k>[ 8�:�&�����i���z{S���{Z����/������qctWR�ʳϖ�s�d�'�|�v�$��k?�E��k����w�S˖���u�n Vhy.[v����W�V�J��%Kz�����V�N�����/����(��)=�P13wn&5eʻ��P�7##�ڞ=�z�M=yT;}X�={~�����O_�� 8l:����t��R�)��?�+}�ѹ�{W(�˗�o��@htt+q(��F��{G�����q�J��O��љ����6��^ ��@K{|��s�n�z~h!������k�7b��1#�=���Z3��O=U�_pAWG�g�w�a}��Y3 8,:��f�N+]����>�5;٢x_���ʓO�U7m���_3/�X����)S.������� 8,:в�\��ɯ�~fh!�+��N����
Q�V��~�T~��R(�l=�ݩ׃8?|f�޽�U�>��w�	 �ohY3�����-��=��|���w�^5���/WJ�<2��D S�v�IV�- �	t�%=�bŕ�6o>�U�OS�&��]�����uk��������Cdf��}�W���w��f �}�@K����7��X=O�T[��;�:xwJ�z��G�*/�P6��ܢ1����l>�� ��"Ё��~Ŋk&m�|B��Z����]��.U�x�R~��b����!r���Y�~�깋�c{ �=�@˙�o_묞���s^�8d���z��(V_y�������8��ͧ�< �	t��<�|�u��7/-��Lm/Z�̈́T_z�\���)���g���W?�z���ck �=�@K�58�2�3ٓO�e,���PT���=Vy��R ZR�V�MN��& �t�e<�bŇ{7m:)��TWW*�����~�w�J��;R߳�Yshq���fݒ%���w�P �]�@˘=:��C��{��袮TO���?��-�_�z1YA@��T*=h4�e�� �kh	.[v�m��- 3{v&w����;jT*����g�}������_�� xW:��˿�������J��e�u�t�%V���dJ{��Gj;vx�m(W,N_02��ͧ�= ���b�x�y�i�v]Z@��S�|���w�ص�:z�]�ax�yshc3����A��k^Dћ�h�r�\��Z6��_pAW�mU_{�R���Q�͡��8p�˖-9ݺ� �L�Qk�tSz۽��
- w�y�ԤIý��sϕ����m�b���?k~� �@���SO��c��!v}}��9�?��h����b�g��(���?��+N�x�ڗ �D�Q�64�B�_|qW*�3�����*V_xA�C'����J�_j>�L ��t Z��Z�p�ƍ'�ȥf���N:)�;I�?�`����s�`S��r��>�[���JE�C ЁhM���
L����p�U�;�Z�t���8B�\��ٶ����� ��:����3��x��̜9�����@���7Z}�Uq4���䨒@8^TQZ0<����ؔ��v�T��y�^o��[7Z{�5q�P���iɑ�K�� �O%Ё(M�!D.3o^6{�Ξ'��g��9�������O5��z ��@t�q���m�|Z�\���]����㏏�����/n�t�o�n�� xG�Όb�b��=;�=��C�*�?_*?�D) ��|�4��'�\�|z{ �yq	Dg����!r�.(8{B��W��*��a���?��@T�X���ܦM�C��3f�����g�k۶U���7� �L<sݒ%���w�P �m	t *�GG���.Z�������=��4j� p(ҵZnn*����� x[�ʤ���C�R==�܉'v��yr�����6FG-��ʤ��A��#�D�U��ɿ������gB&�ѫ��o~��lo �R߁���ʕS?z�]� ?A���9p�?D,�Ʉ���C���R����NxOҵZv����5��� �O�@7ݔ�瞨��gN>9�������T߽�V���Mlޗ��� �ޖ@���SO-]P*M˝uVǮ�7�����w��jչs�}�<u�7�\t뭻 ?B�Q�:6�����ٙ����=��o��� �>���L~p0��? ~DǾ��qp{�ڵ煈e�<�cW��[�T*/���9p��8�ls� ?F�GܓO?������|>�9�Ď�F����׊�ag;p��8p�7��{�-�� ~H�G\_��4D,w�)�T3�C�<��h��[ہ�*��^ٻ����[ ?$Ё#�wx8���'�ܑ����^�T���J ��Ʈ
�Gt��zt���=��>?D*5mZ:=gN&t�dk{��G�8�>; �#:pD����z�w�gO9%R����^y���訃���)�3[����� �A8�zFF.˝tR.t��޽��sϕ�8�[�� ��"Ё#���N��̛�MM��q��K��F�Q���6it�� �	t��y���?rR�׫e:p����k�ڦM� 0��������<�5� Ё#hZ��,�*�
�:+Ы�F�� $]�����U�_	 t���97D*3wn&5iR����C��gJ��!w���T�"t��:pD��ߟ�~��cB��'��Qw�'תU����	�S,F;�`�	t��)/�]�E��<��v����sϕŢkՀ	�5<<�9t���Q/@�x��˗�H�f�J��w���F�l�8bR�zfZ����{@����],�"�=�����X��w��GTo�|i� 82�GG�He�=6ڭ����s �ccg :0���Ss7Fy�y��+��3�c��W�="�}����M7�S7��&	��	t`��T�W�He�9&2�T��Z���3Vρ#.S�v���n>�N �`�p�b��!R�CT_{���zD��ZM�C�@G��@<���B�2G�1���=W ��;7 t��y!
�!����7g����SS�t����޽�ڶm� ��bqA �p�P}����^O�e�=�c�'V��v��ȏ��|�ӟ.���/��t��y1
ġ���P�Tz������\�Vy��J �H�^ϼ�qc�3���CuċQ ݕ�I!R�y�:b{{�WʡT�|D��VKΡt�c	t`B��ƎJuw�R�'G���p�����s J]�ʩ��	t`Bu���Jϛ��T���������aP��:0a��b�1�M�zB�2s�v�����P���#}`�t`���R�He���@�����@����GW��}�w� :�@&L�T:+�(�
�Y��>�mob�h4R�r9y3��@����*�?"��4)
��g{;�
�����\�t$�L�\�2'D(={vۯ�'j��f{;�|�r\ �P�0ٱ�!B��j��u���@����Q�C	t`B<��ߝ{����m���۫�Z- �.[.� J�"S.����=㙙3���y��9�"�Ҵ С:0!ҕ�)!B�L�o�ĵ�ږ-h	�j��5�S	t`B�k��C��M˄t:ʕ�åQ.7�;w����t�|j�@:�@&D3��e�Mk����ρ��U�����p �0��ryn�P���m���@K�T���$Ё	��Tf��;!�w�|��|��� Ё:0!��r�Sy�0 ��{�@ZJ�\� :�@��m�����/�����Ɓ�F�� -$[�N H��nA�:;4�MJO�B������g��s���j�(��ow�J%�q==�������a԰�hA�j�; t ���t�e�;�f����h͚b � w�o4QNp}}��v	t�%�FG�7w_ D��.[��Juu����P�7���@*d��$w�t���\�>=D(���ց�m4jЁU��j�8w�z}j�Qww[oqo��s�e����t`�e��(=����+�����t����q$Ёq���'�����Ȉt�ee#=0�:0�R�zW�P:�o�@�@�J7�B:�@�_��1���=�mqZW�� F��.�hdB�R�Bhg���,뛻 �H���q~��f�z=�JVЁ����!Ё��f���#�T�oq��ha�:�q�|���t�[�C&�O�)���-+�u*Ё|��]�g�S����+�Z�@�r�D�zt��J�C۳�ha�Dw�����J�
:в��/O���.�@o����z�ahai�t �����~���^w:���6'�'	t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@ xc�z��h����N��t� h{ ���̮ry֑��q>6�P� h{ ��f2��lv�`�:5 �8�  ?Ŵ\n�Z�gF��I Ƒ@ �f
���R�T�w ' �gH��8�P�5P,U! `t �C��>��k���؜z�  ��@ 8D�T�zT����RiN8�� ��@hc�f@��j��\W:]ʤR�����;�g����k ��ЦJ�z~W�4�B.@�I�Gz�щ�3]��x� m�X.wm/��[pis]�tqv���H�ٮ_�p� m�V��GJ��Z�b�m��N�%�Տ����5 '��&��jn��:@>�.%q�:8j��q� ��@hq�F#526�]�ם5�#4_�T���w%מ��~��E���J����Usg�����)vN���C��5 �ТFK��r�jK-�q�M����HVғ�Ut �+��b��Z&Y5o4� "��d�:�NWB��Q��Y*�� �����˅�JŴh:M2���B:]J���!q�@ �t�P����cc=�F����1;��ՕN�B�!�v�J�Mp�p� �s}�lf.��'�)�%q��T�U�� �)ק���r{�����7K��c�zw ��D�D��it�������p�ԮRiF�^����J�D��it�f�N��B��T*�F���  ��@���� ��t���\n���Je�jur �q �"��4�;��U(���T&U�S ��p�>�V!�����w'Pr�����޺u���־"6!�@�ق��8�$�U,���L��=g�9�%3��ɛ����x&�M���l��xc1#��lf�@hi��[�w���/T�,KH���ߪ��{�$Cw�������C�ðk$ �"��Ev��w�f#8t��mW�zސU;��<�0��Vg
  F�@�q|�;�eUM��Rf�� �&!���8>���&��qn�Db�ry۪����+ �It h�O~'��pn&3�XV(�DQz[�B� ��@���4�������m)�
�@~�t����  4� ��i���yڶ}1PE��JeN$��
 ��#��A�R����ߣf���=ۮ���(�u��� Z�@ � Sځ=��<�8e1���-��@�7�  -C� ��tݝ9�)������R��+�&� ��"� @C��R#��T^T��J�W ��t  �0}��h�뎋��*���(�
   � @Ct��Ā뎉�vT�3JQ�  A� �i�y~���C��@>�  ��  `Zem����j���&��W  0�  ��g��ٞ�C5��=cA�/  �@  �"mە��7d�6G7O>�F�`P  0�  �,���M��bfwT�3  ��  `J�`^&����@�0�U��  ��  ���Q���m�e�b�ry���  G� �Co4��\��@�(r�U*�U�}  �G� �C�t�{�]�Q��Z��!� IB� ��R����ۮ��B��Qmy<  �A� �I��N��9NIG���\�r� H ~x ��6��]�S�8�\*�	D\  �t  pP�S���T*/R"ֶJeV�i  �t  p@q�������(�  	F� �wԝJM��j{�2�EY  �t  �_9�.�tݝb�8��Q�%  �  �SƶK�<oX����Q�#  �	  ���mW�x�v����<#��7} @!� ��o�s=o��8���� �  ��  v�o�y�̐];V�<A�5� @"� @M���r,+�0;��3 �6E�  �D����͵�@T
��P�:Kj_*  �@ ����<m۾�Ei� �	t  :����=ۮ���(Jm�Tf��|  �� @�R����ۮ���(r�T*s#G  � :  j����$
�r�V*s�s @'!� �@��ΞT� ��܎�|v �
  �@ ����R�}�;!R"��s_��  �at  :HO*5>�cb ��*�Y�(� �D� �!�l;?�uG�PC���re �E� ���]��y�b��ʌR� �F� ��<�.���b�a�(DQ�  ��t  �Xڶ+s=oȪ-�6�N���^  :  �*�!_59��|�g<�  ��  �!G$���ٵc��3]#A0(  `7 �6Gy8��9���
a����  ~� @�D"�mb�Rf�W��9  �@� �>T�mA�"�rl˒�R��W�y+��ry۪��R{  �@ �=�l��q���ݶm�+�ű�(��S�]�[#��J��U*�9  �@ �d�h,�T�@�\EV�+���r�ߧG�u�����r��Q��q����  ���  $���q�W��c)�� ��)ǩE�mw��!�o/T��Z�̉j� �wB� �`^M��*5����n�W�������1��1�r{K�<'�~ ���L  *E��*���^���G�-�*��@hY�  ��B� �@n�^�@*��e�G�9  �B� �0)�ʙ(�C�l�/��  �I!� H'�*z�v1T�q�B��  L� @B�QT�EѨ�d۽�ee   �p���yٶ{��
  8d:  ���
rQ4"����S��.߶s  ��@ �`�Ra-Ε22Ϋ����v�  �)#� 0�R���8�#1�oۙ�m�
  �:  R��8�m�B1P`�^ɲ�,  Ӆ@ �0:��ȹ�T 
,+]�qn��  L'  ��8M)勁�8w���oQ�  L;  �d�h<��(��T�8 �at  �ḫTYY�S���,[  @C�  �����R%1����8 ��t  Z̍�B:��b�H�.�qG�#  ��t  Z(E�L��@J�*;NdY�/  ��� �ERJ��Q4.�һ��q�
  h
 ��������綝  �4:  Mǹ��:C��/�,O  @S�  4��T���U[�m������  �t:  Mb)���[VV  @K�  4�RQW�#=Ul�ˏ/  -C� �h��yղ�U��  �R:  �bq���J�b ߶3��  �r:  ��\���(����J��g	  0� @��K)U��.�6q �At   Ec�(����8w����9} �At  �Y:'\��b�вR%�1  F!� �F�(�{J�@�e9E�˲  �@ `��QT��� Rq��  ��@ `�J�2Q4!R"���8�  �"� �"'�*q����t��g �,~� `8~X@�ahEJ�	W�����:C����8w�������D hk: L#��AP���=G)?kz��vZ�h�ue�XLg���� �- ��5��8W��w��:Ȇ�U�En�����	�F�ZM�a�t{��h: �' ������wK�0E��y�qz��ڎ~#P��g=/ȥӌ�@�!�`
��Ӫ�;Q1j�)��jq?��ʶ��[VV��J�JJ�)؝���e�F `�t 8DLi�<���<�C�@e���m�K���M�S��T��7�  �C��!`J{��q�G����V\����8݂��gJLy�6A��$0��c�8M)勁|��Tl�Wб��w=�ޓ�2� �@��Ĕ�Ε���8Ϋb�����m�	:��գ���d2�� 	E��A�@ǹ#�8^��q^��-��w�P�g��H�#=�F�  �? ���+�i�Jb�вRE��b�P.�a�]�Ǻt H ����-EyO��(�,�8ǁ����Ql�K�� �`Xo���q�{QT)˲u�K�(��ץ�f�UǶ�t 0� {�q�G�)�T��	1���mƏ���A��Kכ�q^: ��@�=�͉��ޱ]�D��m��8z6�>/=I��ccG�s���;��� @� �`6��lvU�Y�b ��8�#�r��y\�z.�6�(r<��������o��� � : H{ĹU���퍠�e���߀"�o��(2rZ��[Vƶ��V�,0J��H*���3	;�{A`-ܰ���>��n�� m�@���i���mWu���ʶU6����W;�-�<��M�R�tM�𮧽wg2���T�z�'߸��%_��w�
 �1@�R���U��_�z�w1܌��t��G_���+g�������CE��H���8���q�z���\��H��ysߋ?����e m�@�qt��K%��8��g�'!����ү�}����B �� :���8��t:���tJJ��wU?������.�����
 �@Ǩǹ�e� ~_=���t�2�U2֜���?�ɇ�r�M�	 �@G�q>^*��04�� ZLG�~�4}$��Xt�O?��{��r��h':���wk�Mk'����n���s�l�y��{���$ �&t mo�\N�N ��{�\vM?'}�sϝx�y������� � ����L}�) �I��[���<��)�Nɜ����q�����A  �t mKǹ�� �!)W�)�a\.�66һK%g���7�O� �@Ж��M%q SW�TR�e���b�y�7�\���{�y� @�� �N9s}C) �iQ(�]'�t7���P�=��}���W����� H(n`����� ����_[��k�m+1P*������{���&�^�T:����:� ��!�ۯ��l��ץ�h������>?=Y  �t mC�uE��w� ��0�E��g�/|�ٕ�|��]q�-� H@[�;�s�9 4�>�Ro�i���nI�#�|㟯���/]sME  At �ǎ� �\���>ct4=����OW	 $� ��H;�@��9]ǉL�4n�sϭ��������w
 $7� Ko
��T� Z$�kgw1��V�s��#� �@�X�ƐM� �u�����;���@�6o����>t�_�uק �@�H�j���� �Rz�t*ŗ����>��Ǯ�����k��, `8@���"S���J%�r�Ho'��.���/�p_�t� ��t �����r�8 ���F��������Q�x���ꭷ�% `0@�*֝��j��=�C�{����3 F�H}��y� `.}쥗J�&�6��7����/�{�M �P:��`j; ��ԣ�����O?}U�@�0� ��I�����l���;�5nW������?��5}�]	 �@`<}���M
  ��k�>z��]�g<��'���K��Uƭ� nx�@�@�(�,=ս7�5n�����������~Z �0��0��&�G� �(~��rS�H3���?v�W^�(: �� �)e��U^�  ��;�JU�0���_?����' / c�q�1 $�~7vø��� �at F
�M�� �x�n�Gѯ��?��w��9 Cp��H�J�3�����+9]�g�z��������: ��7 @[�3��4wǶ�E��}{���;����m��� �t �)2� ڎ��ޓ��b���^�j�@�07� ��G�9V �O5���a�q�:vmΦM�x���ꭷ�% �b: �0z �K���mX�;Q$=o����� -ƍ0 c0z �z6��[��������]_]��  �B: c0z ���wg2F�E�V*vjh����O	 �7� ���9 t=�����s��6n�3�#�����@��;��6�>{h���.8�+���) �"�h�0�,�=��a�(���x�6���)��et -�w� @G���q�P2c�Fvr�R:���g�
 �����L��b���y�}�on��j� ���=��� @G�v-orS)��E�n�����@�:���0� :V%�}��7	 ���e��j� �����K%�k�����g�&#���� �H���Qk�3[�|.~ �4��e|F����BM���[�	 � ��%��@l �K����c��LsH}������  �D:���p� `�3!�Nb��qj���?� ��@�Lo ��YU�N�I��m;^ ��t M��v ���4�H)ˤ��������/�����# MB�h�*�� �������V��7���~Y �It MWe�9 `/&���� @� �J����v ���4w��X�9?"r۷/ h"@S�9 `t���T$��߹3��W\�}�k* M@�h��N�  �E�+bL����Ro����� h@S�͗  �&����� ��@�4�ctX ��[ˌ�! �$:��	�s ��ah٩�9�>:�# �$:��a�9 �@L[�ޛϻ��zu�W׮- 4��iX 8����>RQ$n�pq��� F�h
}�-�� ����s!�4��)BF� A���7���cc�
 4��)�  p��Fqb�t�0  �:��	t �A���k��c���3 M@�h
�6� ���,�q�]��� �� Ma�zB ����+ˠ@�|����|�]_Z��y�"�4;� �~Sל<�*΍t E�h8F� ����5-�S��) F�h8F� �e�ώRi� @�� �t �d����*� �@�p� �$���$��� F�h�0	t �����S.g �@�p�b 09ƍ�W�i�#�  `�ݭV]�#�4\|��: `RL���\@� δQ  &ˊ82@��   0�io�::�& �4\��pW H2F�4�   �E �F�@�8�DJ���|VmO% ͔��R�?��T HČ�h@��x;�&e۾ hk�(4D��M{��`t��1 �G�h8}�e�] �x�&Ёt ��M `Rt ��@�p��a��� `��g�Q�nY�_ ��t �( `����� ��, �!�g��C�h8�v� �Oq�8�D�h�0�t ���o�_b֠h@��7Y�pc ���7wt @�: `��04*�A�:�����tZ  8Xq�S� :���|�FA  ��Ȩ@g@3� �M�  �p�
�C���ᘦ ��H��0��t Mዸn� �wV	CWC�h@S�J�]�"� �!�� :/~ ����k܀ �@��g���s �bԋ��U��"� ����@�,:���;� (qL<bM	 4��)�Nm�6� `ߪQ��� ��@�4z�8ϲ� �~�?+�[�w �B�h�J�=�!� �U�V�?бx�4�M�ۛ�
  �cZ�3z���z���.Ge��V��| �?P�2�G���t M�o�|�tZ�"  ����ƶ9�@�� ���^�qt �(��h:��*V�i֡ �E/��� ��@�T�j�f: `o��?7�kОt M�op*Je2�U  v)�~F���sF�4�����j&�y: `�|���� ��@�t�rٝ�yLs ��>� 0���s �@�h:�� �T�}�v%����%�� �3qz;�h@K�i�3=O  ����q��5F����%�4��RY��@g+A"��s��f ���D��e�; t��r9��Q�:��ɗJ���c+
 �㔢(��q���s �B�h�|t�:θ  :�x���0R��t -5V,z�== �,A|Z�T1�� Z�@�Rzj#��@���~��@�J:���S3�� d�T2ns8��h5@��e'�fݔR�  �^!���(2��g�3�9f@3� �0Z.w��� ���Rɸ��5F��������y�Tm�  @�*FQ����-�>��s�f@�� �1����;* ��5Z*w���N��5��q ��@`��b1�����J� h;�(ʚ8z~0S�#��h�1�<��jw��	 �팖�F�v�����h�QF�E���߶�� �6*Je�ժq���������% G�0�E�V{Y� �eg��-�rmy�N� �@`��B!�30��� �&��禎����X�J�?
��#�ig��3;��) �DS"��B�ȝ����̞N�1��#��P.�*���,�, ����� ���`Gϵ�u+ F�0�p��=���@��
�)3b {��G�̸ @�� �������l�  ���Tz��&���zˮ 4��h��|.��W��5 H���7Q*�b�Ɏ�ka&�U ��t F��.��fzވ  cG��#�:�@�L�e�#�O�����l 	1���z��HǹeM~�:;��_ ��t ���P�Y��SS3 j|�ԍ�ɮ=ע8�+��� �@�~X#�j߀�
 �X;��>S�K=���J.~�[�*
 4� 1F�t����*�Y� `��0�)W�FNm�e�\+wuU ��@�(C�|��������3 С�����|Vu�q�����)t �R�}k���� �1yj���P��k~O�F�& �$������e-��� `���oǩ�uaOϣ M@�H�����E}}[�P  -S���~�T�G��X�=E��- M@�H�(�d[�00/��! ��E���|�l����l6���� h@b��c�t__*5& ���Q*��Q4����q>�����`^�xC �t ��3��f~������%d�; 4�X�+��O7�T7���Θ� @�� -�h�Ȋ]9����[ @Õ���7H�`S��^����A��!�$Z�)��>�'8�؞��hX~�ɪ  F�w�m|��u�z�|�S�5�7��Z �It ��J��GמGQd٧������x��� � Qܾ���~S�;�t�O��y���z�w�� @�� �������!� ����g���׏D##�  ��P�4�����i��ZqΜ-��K �B�H$'������߯�v*w�y����Ǣ|��! H���j�R���k4]S��*3f�' �D:�D�]�R�tz�wae���;�{�[�R�� 0E�a�3V,��`�9�]�������* �D:�ı����Nz���ݝ���GT�{��+� ��)DQ���DV7�q�+�^w�� MD�H��w�KR==��X���>[ K�`�*Je��ǻ�p:Χsj�V�;w���� @3� �ժ���R��hQW�>���  ZU��2>�+�����5ݪ3f�- �d:�D�-Y"ޜ9=L��_�.]���z��+ 8 }��汱>��SӦ{�y]�J���� 4� Q�O9e�������c{��ձ�/Y �~E��l�7=εFĹ6�`�ȧ��z� @�� #=c��8��� l���ra8V�կ�t ؇ �7�:11���g�k�Xw^W^��'��c �F�H=znM�n��};u�I}�(+=�4[��j#�q��A`|�7jݹ����{{�V �t ���r�s�qS�8z$=�jU_�q� P�Gη��'b�Q����,�5o	 � � �N:Ilם�G�re_��$ ��j����DĹ�J5����p�ϙ��Ut Ƴ⛱��+��c�H/s��\Q �C��ڷNL��oGE��_ h��z�/�TW״�<������l�dY����4
,�ջ�')��)\�؂c�^wݛ -B�0[|3ֿjU�>��H���re۲"�PQ*�el�7	G�i�ܱ}O�E�n�� h����^q�9�9��B&��cۡ @+)��6>ޝ�8o��{*�r��+V���v� @�� �揍ɖ�fi�y�)�q6|ߨ��]]��m mh<{�'&���ޱ}O#G�_uUY ��t W��}�x��e���\���9���ם�Y��pN:���yo�I���.�?Wy��/ ����j�a(S�N��%�����s�mx���t.��<׭
 $\��kW*���+	��8�F.�˛n�G ��t M�o�� �Z����l�?Μ��^,�� �L�� +�,g[�0P�V��{53ε�ᇯ�'� h5@�LG�O<��D������Pv*��H���G�>+�c� $�oY����ޤ�V��8/wwK�/���V�V#�4���#}*jkҿ��ښt�uz�wx+��� I
QԵ}b�+);��5��uԯ������t MU_W8�H�Uټ~����ǔ�N7�n���{.��Y��tcAз3��$aZ���ܹ� A�h����o��[n�yq�;�L������0���.�q"{�T,U*�Zo��"ε�c�y���A �:����HߴI6�]+�?�q���6��R��֥wg�e۲��8 �F�2C�|O�֛k���(�R�/ 0��e�+ҫ;vȦ5kd�(oΜ�����X>���媜��Ւv���Z�ڎ��~���L � :����H�yy��k�ݳ6�nO����S���>Bm�XH�v��q9�-�L �0:���7h��N���\��n�If�}��]��)w}zʻz�;��h��R٭cc=Iۥ���q�y��׭�O �0: cL�9�*����y����f������w��(6vy��5��}��BZ��q�l[£���<�� �it F��H��eٰA��Q�s�9?+�N����y���3��Z �U���^?��V_��jÇ����~�N ��U �2-�˿��2�#Q�������o��~��t �E����~�H������L��0�RGu�l�  `�ֿR�>��0���)}��[oɛ�]'s�H�.XдQ'=�^�+��p�C�[��mb"���)q��8�g�r��{ eƫ% ��8�ǩFzm��u�d�=�Q���ִ�� l}�� &�F�5۶w���Z%��Gq� ��t F�7vz�E��O��#���j�����?�f�K�M0U���B�����5���tS�Xq����� �� ��o�t�O��tm��g��}��=�<�h�hz���l:͹� �@7�H��;Q*��p�����`e�I'}T~�C �� ���Q��Ou�ʶm�u�����c�m�U�Rq*�j�+��]�� bQ�3<1�M��{j�1j�2z�	_��UWM�]^ h0@b�#}:vx�*�z��RڸQ���?;�j��d��[�b1�n*�yL{:�>:mG��S�}s���I���id��Kׯ�� 	`ޫ( ��t$�Vkg�O��SOIy�V�{�*=8��!}$ۘ�g��L�q݊ ��eզ�����ή��ܞ�TJ�-]z�<�� @� ��Y�#[�Cɿ�Ҕ>V%�7���d�{߫�W�j���R���Sߙ��CfYV�Je���ߨ�������YM�aw�Lg�L[o���+V<p��7�H  !t ��x�5����·������~�������\
��������jj�ק��7��>��P�d�#��t�W:I���l!��0�ah��)0q�y���Y�E����ɏ, �:�D�o�g�!���Ֆ�n��X���+����q�2��V]G����(�v�O�ǲ�_ �Ӂ��(��ü�֙��(��i�(���+W^q>�H@[�Z��Z��Ϫ-����7o���
ټ~�t/[�f�}�8�L��@���Q��z�>�����\X����.{���y�������{Z���׭�V  at m#��g-^�Zm��Od�駧���/�(�M�d�?���.m�0Q�Z�˖v�0��TQ���;R.��K����2yJ{]a`��-]z���� I�v?8 t6+���s�tq���.	�S[����{ߓ�NP3?�����kU�w�+K��j�07}J{]};W����o~3/ �@m� ��c����-?����xc�o��g���2���W�˗����L}̡���,���r[�W%aJ{����ͥ7���	 $T[�  ���}�3j���d�=��
�)}<�6}�w��j֟���}}-���w�t�j[#�@3��jqD&Z��{�}���iGI��^71kV�O<I�W  �t mM��>p�)�Y�Pm��v�w���,��7n��SOU���.��:Գ��F�8�۞ڻ ޑ��>��:���=0P;�{���J�8�a���:Γ"p]U8唏�񵯕 ,9�� 0�y�%����~｢GԧJ�������K2�O�De-j����=�2�㨬���HU L;��d��9�،������e�����Oҳf��?��D�d���춝�����[.��w� H8@ǰ]ך��J���P|�7����Аl���Y����\������a�u˲��y��^�(��J !���p��I���?ܵ�אw�g{�;��fϮ�8�u�-i��u;�>���o��S m y�� 0E=�c�,Q��[��qlj�������/H��Wj��N;M�T�������ܹi5oތ�Yg�W��'�,Gccl*�A>��u�q9k�<��堿��Y���_���uW�ƤH⨹V����?���_	 �@Gr<Ϛ��K���j�~4-�]�i��='3��^�}�1�5��Bq�KU�-[֛:�؞��7%��o��Mj�oL'���FFrf�t�ҥ��ҥi�d�Vm����F�͓�_�BTd��I5�B�Q;���/~~ݺ- m"��� 0Mr��֦���/e��G��F�����&���|�>����u�R�,\(�ŋ�L�(᫯J���%��Y�aEQ����,�稣�q�Oz��?�ޠ��S%3��z��Ӳ�f�%uԼn��U?��7�� @!�t<�6}�> =K��Fӫ;vL��-o�R[���z��3B=�$�dD�;N��6���kRٴI��twѢ���]]�a����R�ͩߠ[t�%J�iW��cHҹ��3t�1/��	 � v�.\h-��R5�a��|�ڔ�)SJ��M�h���W�g�����T�:n�"I-^,^�b���-[�S��Fr��={�Ҝ,]�Q}}�{�f�-Ouw[>�鷏b{��}o���:̓r����͝[�,Y.<  �nt ؃�JY3�菤oŊڑl�>;-W��;��S2��sҿr�8�tq��M��k�=����$}���J��z-փ�+��RG��������)բ:���͝��~�������Z��;Y����׬) �! �����{�N8A����6�]�ʏ<�Hm���U����S���������,[&��k|���_���u���,ϳ����%K�j�|7.Sc��Y���fά�Vn��k�0�B�U#���Wq�?# Цt x]K��6�}�	�q��U*��q������2��c���o�z6+�	���]]"˗K��Dv�h�f�n�(A�yF��{zj#�jѢ��Q�G�M]���9�Zx���5kv^z�Lg�-�����S��o�� @#�� ,Ǳ��^�L��g�z�q-���Z�����POuw��j#냃�+�v�,і-���T�x�6�h�8����۲xqV-��̙��I���O��/��C5,Γ�;��l]��ы���� �� IO{_�яJi�f���{�G�t��Qu���}+V�F�ݾ>1Um'�t��f=u��QJB�6I巿���Q�~�牷h�8��y�J�R����0�T�����96�ȵv�ξ��#��z��~v� @ �`����[�W���믫�w�-���i��z�z-ԟxB��K�>Gy�1����vWs�_ݧ�&jxX�8փ�[ŏ/��m8D��I�(_�@��{!����>�\��@X*�����KX.7�s�0�W�Lg��آEc�O?�HٰA �� nb����7��6�u��V�s�S��>+;�wZG�t�N<�|��.\X���;��D܀A�Nz�?���/���##m�.�okG7N�vhKvW����+�q�*���2P��-���ܩ�mzԼQ��n��^�g�.�����ϸ�j�� �:��[��h��7�o��%m&�1����Y�L�<�h�����H���i�����ś=[�N:Iz�;Nlו$�M��Ov{�cr���ھݷ�z�Rݸ1�n��zt�Toomd\_�������愱�ߝ��שX��Wk�`�76�ko�0�JՑO<������#4  !t w�w�����.;v��_�ٱì3ŦI�֌3ΐ�OT�zӷ'���Q3=�~��?�����+�o�Jq��%Itx��g�࠾���*�Td����m���P��ysML$��p��L��C|�,q�G�yoo@(��<L�f�Q����k}��m��� �Ogog����+��ºu� �0:���������K/=���/΍���k���Y����eƙg�����y>�#�z����裏֦���t�d�,I�hZfVe�̜����|y��J)�R	Վ�54T��m�-[�(�'�&��#�ٳŞ1C��3Ŏ�<�㲾�[-��?Ae۶��o�=7���{�0ׂL&�8����v�} �mo����k�}��V�>�~��f
���jxN6k�<�,X��a��ש^~�v�t=���jKu%w%An���o����n|��NP��(�\~;ڷo�:ڷo���q%l@�zzd<�;��!?�ˎ�\��I^r���Y�h�>jq쩧��ysC?W'�����z�_��ڵ7	 t(@S�7^?�#�������L��֑��C��䓕��ڈP���Q��/d�HבGJ�'J��å֨�F��Kǖ9s���E{ZG�����P����h����
v�؈�1��q��Ċ/[_��qGd�Ǜ%�gm��Im���gd��g:Z�uZ�k:·�:�?}����. ��t MG�m�^x��f���g; ҵT.����)�(�z�F���P�/�T�����˥7��3fH;��"�tw��˓��Q�8�=ێ�|>��x���@FG}dD���ؘ�j5�øf{^mD\o�f��j׮ W��{���{d<j��A����?/z}�t��?�暎�g��w�|� �p:������oב>+��L�D��d2����Gf�q���󡇬��lRLL��Cծ�������Ү����pwݔ�i����Y�ʉȍ� ��P�T>X�bǼ��]�s�������J�Ƿ_V:-V6+v�ˉ��8���R�?�#��������@^y�6R^|��R�F�]��g������? �@�::ү��g.���_^�J5d�R�x6}��У�����a�O��՗>�]O}�9�X�:�(��H��F��N�o���A_���q�t �z>~.q�I�Y�J���ڣT*�}W�R�J�W�\�JEſV���M��\W�L�rzzlg`@?��^���{���G[�1�+������G��I�Jg�G�'^x��S�����Z�y�����+�p��`@K]�nݍ��zuiƃ����3����8��U޺Uvơ�#�Q�v�����r:��z��w�KrG!v��$��v���jI����71tTբ>~n����~{����h�CO_:�j��a�k;~�G�k��a�DGZ:]�������q�ڙ���?������G���8����n�5��v]u���}�����_��o~#a�дϭ�\��w2?�����%7�� ���wc ��פ��g>�'�6l�I���+*3w��?�\���^y�Q晆�S��qX����k�u�wsLm���F���y��_���^C�Z_���\ϲ}���4������d�2�;u}���8����7�H��^t F�|ݺ���袳Ԇ�w��tt�}}��R����I��e��':�]ӣ�zzo|��ܒ%ҽtim��+2�$�Ǣ����\_a�����������˅Cg�y��7�p�  � ����Y�ȿ^x�J��c����Ѿ;�$���^+�����#���Xo䨺�G�wO��m�,\X]���Y�0]�ϫz�7n�Vl��4�?T���G�8��?�f�O �O: �\~��/���a���#/��f��F�6���}T[�F�5�����K6���c�+���a�Im}4�bz������Rx�U}fyKv�g�|�
�f��O:��ϭY�  ��@`�������W�����/���B�n{��O���l����L�F���d�'j�]OϞ]����Eb1b�&�GG��T���:̛����0Z���-Y��]��]�M  �@`�_s���^|�?���'�<��?���T��#��&o�G�+[�֮�j��Qu}�/����ǁ���gs�(ׁ�J�~D���v��o�/?����G �A �풟�����gw�~��?�رz���j�ժX���x�3��4'��̂�+�p�d��c���6I)���[oIuǎ�L[�;�OB��jۊ�����N�_�J  �@`��w����?�ڰ�
�Ze����a6u
���n����4}��uo�<��?_��d2�yB� ��А�u��*���b�|���g�)��~�� L
� .���/�ӟ���o�v�Y铡�BO���ꪅ#�z����K_��@I��8�k���T�hoc��?<,�-[���H�A^��\���B������T��h�������|� ��� ��n�ޚ�����<�xN�Gp��4!�k�ϯ������]�-=>=c���̑�5wn�h7��������Q�U��}{-���Vn�?�(g]��+VFW���Ϯ[�1j p�t �r�7��ʚի�o޶�Ł-[x��q'=IF��.z�q�%��]�����*��>n��8sf����@o�7m�w�J��8�+q��_+���`����y�[�-Z~��u; p�t �s�ڵ��aњl��eo����Vi�h�8i�s�HO��]�W^����p��S�࠸z����To�>���,,�����W���^{�Ϥ)���ק���[��X��'~���e� L� �.��ι�3�����z��g:��S��s�`7et��pף��8nK���=�קGߥ�_:���~q����_���E���z3����s��S�'��h�i�}�����
 `Z� ��u���������g}�]�܁O�=�F�3֍�=(��y���}���_q��Tw�8��=����l�vD������Ӽ^��G��|^�BA��һ�����;��_Gժ��z�3u�q�z�U�>��u�� ��!�$��֮}�_��/�O=�̱��u�щ*�u=֣(�g��u�:H�(/�q��X���qqv:��c���_����ka���z���?���>^=j�8ֱ�{��^z���{:�����֣�ah��"\�o��jA��9ߗv��9�䍥ߞ�y�1o�-Z������ ��"�����[�B�]����#{�+�O>���T��G{҃�����Qg�a��ۼy�tZ�X���շ��i 4�����喿��'?y���w�sĪU�n?w�M��`Oʔx��5�f(̜Y=�O^�n� �0:��s�M7=������'���1����;�x��lﵿI[Î�!���,[������]uUQ  E�hK�UW�֧}���������y�c'|��$�{{=҉�ζ�4u������Fç��O�_���� ��t m��o�/k/�t��l8fٲ9م) �Cl�h��B{�3�O��E���˗��%k�<" ��!�����^�1~�w]_߿,ݺ��9'��P���7�J�'#����9�ğ|�G?��<�  ��@�1.Y����r�%��v�=�8f��~o��!�)ܵ����{s��,��3�p���ҥ���7�' �� �t��_wݯ���]]7����u�)��8�E�k�|]=������o�
�=���F͟|R  �C��H����O��E�0p�}?;v��Y�E���6r0Q�������~�d{����#:������˖�Ǩ9 ��@б._���a�����^��k��;��r]J�CL6N�����Ow�����������6F�NG�W���;�8O�~Z  f �t�o���5���?�x����>��YFӱ{�/!�D��qĶ��G����_��  �B�@��|��a�.�ે���Y|���TO�m����+����JΪ@����:{w !�@� ��sʨ��TTF8#;�g�IUu'3�m�򠻪9�9Td�ħ��qDf�����:.@P���;�T�[�փʖ�Iߪ��ι�ޯ�!��!!�|_}������<�v[  =�1.\�������Æ:*�{���(d��P�V�������>�`�+�y��[ �� �e�W���5מwމ|�Y�d�ܙ�.ҁ�������g��n�r  y�	�s�շ�i�U����E����>���:f��@򆺺F}�����O}jY��7 �A�<�w�[�7k/����6|����_;��uv:���i�j��7�8�ug{���t��a����]w��6�v�-K������;Ϋ��$�����G���E�\|� MI�솳?��{�t�u�{��/}��#=�G!ҁ��86��~�s�;��k�) ��:�8��k�1N�?z�2�k_���gwM;�@��3�<pp��ǿ��O|��� @�� ���7��8}���O��E��_���?�c���:��Ξ=���n8�3�9?l�4;@+� �u��[��}ߵ��~��o[p�1�Y��:0a�b�o>���{�ao?�� h9`�d}}�8�=�z�;������3:��)��B�c;f��|�1_�w��o;K��4�0��C��u��v�}w����ccg.��nzl��#�ڂ@�KN_�~,N�X{�K����?�(�S�:�T�ۯ�(�M;,8s��G ڄ@�������ƣ����+�rgt��:f����m�3gx�s�s���g	s��$����G�/h��N;��j����wN?�� ���c��G��N����' hS`��~�����'��÷/�ַ����:�,��:��Z>=��?���}��m�v֧> ho`Λ~�϶o�#����
Y�ߞ��L�V{�#~6�x�;ξ�����n �+����Y���O8!�7:���'���p�a��|�:��g��r��_�-��3���  �C�$���~y���q=����4>gN��hQ �K-��.ܼ�#n<���.��r ��@H����Gq�d��p�~s�,	�3������MK��9|�A�������O~2 �S� �k<����c��Z-�w�]a�#���1ܳ\. i��_�[-ڴ��C?6#�_~���c v�@h1 6qĮ�;¼��$�j<��iS &��Y�F7/Y�!�x�Eo���[÷� `O	t�&4<sf��B�c�}������0��?��� �]cS�ֶz�C�]s�1���ϖ0Q:@��~����'���+������4dc����2�˅mlٹx��p���~�54�~N ��#�ZD-���,�5��?�a�ڰ!�ݸ1�C7�`�eY�6o���!�|;7oޟ���>���� �[:@�:5<z�	��/�l	]w��k�/~B��'�|�ܹC�/�04g��w�[��!���}A����ٳ��/}�1}ǎ0#�z�����C��:�z#���ܱp������Y7�pS�� �k��͜�����)�_�X�2�G?
��󐍎h������ڲ㠃���?�笫��ݝr &�@hS�7�?��1�g����������)��Zͮ��|�#;.�%?wn錫��/ @B: a��#l>�]��Z-t>�@��яBW��·
u��ӄ�]ڱ`�O�x����˧�;�7�  E�ߐ�r�>���zU�24�6n3~��0;�ԭ[�jdƌ��<�}��[k�g���7�{t�&!�xR#ӧ�G�����y����C���u�ݡ��?��;L��ԩ����oZ��?��s?p�7��� �	t v��y��C/yɮG�gn��� ���8�}~��h�ap���}��)S�\��ғ/��t ���k<?x��F����`����a�ƍaz���fl���^gdY��?l[�0�8䐰c��3^���X,�/ @� L�F��?�/x���Mٱ#L���03�Y7��|�|~t4�[ƦO�<0�xֳ�ТE��|l֬  �B��W�̜F�:*l��^�_V*����s�9)�u���M�^<�G���ó:��E{������A�zd}(�;��i�6 Ю: ���^��8}�W�ߺ��)�o�|f��Л:6o>nʣ�.���3����<��OUuu���s�Ё�
�F�Ϟ ��$��t/��ʑ8]=>~�K�.|xӦ�;�m{Un˖%Ӷn�;m˖S�o�Ȅ{Z��0��~���cx��0�x���9�>eJ  ��@ YoZ��q��ߌ�_�詧��������m�߱�)[�ԱeKW�iS��}�wt����a��ٻ���!�3��P��F� {N��tο�G�t���7�u֬Cxmmh����O�28�8F��8��ǀ�>4��FF|��q4�t͚����{��q�Zϙ��3���G��RN��Ƕ����������ux���Ν/��G憆���?�s笸��1<<5?4�1m��\nt4׬��5�)�M��bX�Μ�k�� ���a4εF�7��Qt �T���k��+N�q�S��[O;m�]�����gg��!c�Ë���룣󲑑��cc����N���2�)cc����)Sj�ldl�#�=S��~}�9��ƗBG�Z-�?��,�5�6����\-�kYVi\g�X.���8������)�cC��S����cӦ�<�SkӦ����?���xI �: <�ׯ�ӆ�U�VT��N��{ ��@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@ �N�^� ��t ��dY6�\.�*�J� �� 4�\.w\�� �Et �)�j�7�@� @Sʲ��8�? @�� @�z^�Ryy�X�j � ���U��q� �� 4�,����������� hr ����h=�˅6����z�����  ML�@���>2u��Юb���Z���� hb ���ٳw�vV�ׯX�j��/_~ �&%���=���C����,
m*~�����>C��u�Y	t hr}}}��J�Ѹ��X�7�}�(.� hB Z@�^0j[��U1ҿ�lt ��@����8�\܇)�z��+����y�{~ ��t hw��@#����~����5}}}; 4	� - F���w�=�˺����H���g� 4� - ����o;%F�Uqo��fw ��@�022�aʔ)��qv�R�+�� �8� -`�ʕ�����,�~Cܓ���~�X��  	� �:�%����^��Z�>T(� H�@��e��@\qo�Z��Jej�X�> @�: ��[�ő��F����k��r�T*]  1 ZD�X|�R��G\�0��#���j5+
� H�@����1B������A��� ��8�"�~u'�\.�K��G $@�@��yG���b��4�T���H�R9�X,V L2� -�^�_%П��OY��1��
��� `�t h13g������������Z�.�����o4 �$� �b.���m�r������ܮh���g,[�lg �}L�@���Z�vNp&��z�����c��#}K �}H�@Z�|��J��ٸ<5��^5<<�����7���� `� Т����*�˽y�Eh솸e�����8����� �� -����;�r��|]`O���\�TN+�7 ��: ��,��:�g�+���HG��� �E ZX��[c\~:.��SS���u�r�٥R�� �� -ntt�='�����o�R9���ki4 `�	t hq+V��'�e%.�x��߲eˢիW��c� �h �@�e�5�E��a�g$��kGFF�r�e���bŊ{ L� m�P(���R\�L��vtt|5��J�� &�@�6C�J�Sq���D84˲��=}s�X�j �gH�@{YZ��/��aN��.��g5�$ �3 ����Ň*�ʅqyS`BdY6-F���j��B��6 �� �fb�&F�uqyv`B�H��H�������] `t hC�|��ccc���&RO�\�ܶmۻ���j v�@�6t�%�<Z�VO��j_n<��0q?/���:������ �&� m�P(|�\.������1�s1��� <] �X�TZS�T^|}o8��k׮=c�ҥ# ��@�6W���4˲�屁��G[�n��z��-[�lg �'!��͕J��J�m1ԿC}��D;eddd}���D: OF� ���~P.���7�150��4<<�����m>��� �.�R�K1��,˲&\��7wvv^#�G��x: �k1�?#����.��]]]��z��q] � �۶m+ň\��������8_ �1: ��_���3�,�%^�,�7��R�<X,�w �q ��7�W��7���������-�ˏĽ��  A� O�P(<���r>��j�<<�7������� @�� ����/�ks�\#�&T�e�8n(�˯.�J� hk xR���?�T*o���_�1�`�͌���_~��.�䒻 mK� O�X,�G������/�&ڂ����]z饿�r��M��$�������;��r���eW`BeYv̔)S�a���'-[�lg ��t �i����z�Ry]\~>�������W��� @�� �n)���>˲����PqO�)���^*�> h+ �m���_���z��Y��W\���{OO�W mC� {�T*}�q<X��Ɲ���	�sJ.�[_�T^\,7 ڂ@ �X��oƈ|M��/Ĩ��0q?������ޗ���� �<� <#�#ت��k��-��L�������j|�� @�� �3V(n������s�&ҹ�r�+�R�#��&��	������/ϲ�qN�с	�t����7����3 в: 0aJ����j��Z��x�����2=�����/�yt��%��	U()��'���8^�1Џ���"./ �$� L�R������;;;��a���D��J��o�b�� @�� �^���7#��鿌��,0!���n����I ��t `���^��{*���bX^C=<#qg�qݺu�^q�駏 Z�@ ��b���Z�n���8*̟?����}���s5 �2� �'
�µ�ryS\~"˲�g�oW�Z���˗o �� �3�R��j���z����{,˲i�Z�ڵk׾t�ҥ#��'��}�P(ܶjժߏq������3�[����� MO� �\�������|#ҟ�c�z�}�j���B�� @S� �����o͚5��1^��#�G�/����}��[�hR �4_|�u�֝z�=�����
�Ϛ5�q�P �i	t `R������J��J�sq�.+��7�J�_ ��@ ���w��vK��q����� @S� @2��J�7.�o�����j�zm�� 4� $�T*}qժU/��j�������������k�>��� �G� �i�V�VOl����vǱ�7o�(�W ��@ �T(~�z��W������'��\.���/���K.��� @�� @��-[���������5Y�-<]�����sO �it  i}}}�qzW�\�Y�/u�����q�>X*�� 4� 4���18h��sJ�L��o�8; �: �4b�_300p�O�ˮ����tF��===�	 $O� M�����j�5�z�q��'������� @�: �t
��7.���W���ޒe����9�R��X,o $M� M�K.�3F���#������7��) �4� 4��w�"������獕J��b���d	t ��uww?p饗�����s1D_x\�w��( �,� 4��+Wn���?)��5"�����-�V�:n��� I� @K����#�1�?c���oˍ���E�� $I� -��W�~�����w�]qON��˺W�Xqo  9 h)˖-�#�u�����cu������ @r: �rV�X�9F��1F��e�K���իW��e�v �"���4�'utt�/_�%˲�###���_ H�@ ZV#ҫ����������~� ��#���V(Y�z�I���_Ͳ�@��V�Z���˗+ �� ��e˖=X�VO���_������q� 	� @[(
?xm.��r��/��,�N���}w__�p  	 h����Y�V�R���)����tvv��� � ���R(��\.���%i����  h;�R���s�,�?�������.�l���� �N� m)F�+��qY�kz>���8_ �t h[[�n����zN\���ۃ@H�@ �V___������|��xy|hCY����5k:/���m�I%�����ӳ�\.�9.�cu^h?S� xY��� @�+�J?�T*g���B{����A�L:� �ś���_gY��L��_ �t `ܶm������1XO�������{zz~ �4 `\�q�W�>{dd�����F�,k<�.�&�@ x�e˖=X�TΫ��7�h�B���r����I#� ~K�X��\.0./
m�^��$ 0�: ��ضm[wWW�k�����,;��.[�bŊ{ �B� <��������vy�=�˽8N`�t �'�����J�rU\�3���@�t `Rt �'�eYw�V{s���s� �K� <�B��H�R���PhqY��  0i: �S8�C>z��w/�{Lhms�����_J �9� �N?���r�����Dhq�z��8	t�I � ��b���Z������e�q�v `��  OC�z�\^�kC���$�  O�ԩS�W[���`�t ��iٲe;���5qY-�t��#� vC�e7����� L
� �
��w���q� ��Y�I!� vC�eq�J�qyFhM`�t ��T���=�zKz�޺ �B�L�����-��'����5�Z�;� �D�L�+Vl����t�,k�@��۴�k�NY�t�H `��  ��X,��l_��k֬�ܺu딽��\xᅣ1� ��@ h_|�}��\�2 ��	t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H��@\��@PD    IEND�B`�PK
     t$v[�kZ��  �  /   images/6608fa58-7afa-4488-b64c-2b761d69d6bd.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  �IDATx��	�U�ǿ��ʪ>�/�FA��V�i<vD@YqWCא��Y�q�Й1�u��	cw5vv����@Ggt=wW�G%D9�� ���>��:�z�}�UM�4ts��������ʪ�z����/*%��@$S�d*�LE ��D2�H�"�T"��@$S�d*�LE ��D2�H�"�T"��@$S�d@v,X ������u�a�y�3!��sp����C�\��0�$-�P�������	���ǡ��2�YV0V�JqS�-��;]���jl���i��l:�L���*8g�z�����A8�pǁj�PUu��
���bg��Q���ld&.6S8NW˅~�p>ö��5�̄L��i�S^6n�%���f��ɓ!���0����_�����\|���wr����(AQT>��G���H"���5l/ۺޮ �C]�ee0���@FI��W_�h	.��:aiZ=��?������'�
��+�m(�(
�;�<�V��<��7��{��&���`綾��@6Ȏy󠼵���cS}���m߇o�`�b���Ex�+'��)��{��8�@:m��Zfs�����5�~����?{6�ߴ	dRA��x�����t�������=-ŷ2^C��\&5�lV���!jn{�koݚ�7o6E"a���h-W���OWQ~�ZW�~g]|��;["(�u�"(9xЃa�j9�U�a�R�x�C(�Q!	�!8����J�WTp��!��Յ̵k���m�/�4Y���b��?�ٽ�Ν%��
���҆*��Yy�ʤI�~商��Y��O�L�Nl*dI�	�G��ٳ�|�X�
�����Q>n\�\��a�D0%��>�Pno>��MQ��_uL��(�
����]���R۟#�� ö�6kVH�??���,W܎��� �A!k۾ݴw�/Եy�f��M��0/)�w�I"p��2���Sn��`�2(p ��.�ҝ;�MA��d��� �A�K/#Ë�7B���̫�&�x�����;PUF�%�rZZ��u�EYY��R�?_�%堘Hw"Ɣ�Fm���0��ud̡C��؀���џB��@7�Μ�!�L��n�P%�dI4��	�J�A=��к������o'�˖���C����Q\��%�ֹ������l�5�NC�8�/�L��E��{�3&�*�t>f��/X`x�a�u2��L��f^��&'���	�k1��LF���ffv?ʆ����v���.�Ik�B�(���c�u���Ơ���:���+�x����qج?�)c�Y�F+�=)aǻ�9���yO�)�i.C0/�`^H
����\�Xk`'���ۧMө�;
����}Xy�4���;����4~�����(���D��;�d�=��"�Ǥ�!*�����k������I�� ��c�?����5k�
Ⱥ%K@mj�[�yf���)v��(��*��h	��ۡ�"ﶾeѾ#h%�s��|4&�R`@�����t�������UaFt����[��.�A�3'O����WWC��DY�w�I06��r��=��+��lֵw�0���\�9�55L8RP $��*Z���x A�-}����wWT�S;� ~jr�B*�6�����  ���6fL%�7�#*Ԏ�����r�P����D�ߝ�)0 X	��f�4�[���A�+��m������:P����)/�*|�^�	�c��}�uM�چAz*�T�K�A��)<E>ӓLR����~&�+��<�:�qL�87��E�!�uZ��X�ǣ���\���7�.K���0�
<S�Ϥ��1�pg:j����)���jBUU��� �Ud	���*'9�0����T6q8W���)�ӾaT�z���t)Ĳ��Bb �� B�����8
���4�,��n*U�F�㔠�U��%�� ҫ�Lw	��ya�Q��oK8N$n�U0L$����1
ap�:=$1^��f�;�*�$�
���鵴ㄆ҈ p��Lg2�S.˹w�k���4�`���������EuSҊR���p�A�@Y�"�EnK0�3��i8a��R�0�𣆖C��o��9���B���s\�H�=���}-�K"���	��ؐ.��{c�LF-	�L�/�k�bY��1e
���W�
<ǎT�BP�T�u�s]��{���ڜ�����k�
2�Rð�
����o��f궽�v�xv�,�~c#���33m���,�5�4���I�	&9�>�Љoy�FxӜ�;�G���w2t�RzY$b�"z����0�����[*��U �CI��J�ٱ���;u2�y(����e"��
�m�뎋:�ӟ�xc�w��G���3a��_BP
���?�MP'��Y�����1�h)d�]�۵L�u�]����y����x�3w{�x�Π3n�ݧR��a�Ŷ��]W���{�Z��ر
�#�sf���ꄂNj�/ʼ���=G0�̜�c�\�k�}�l�+�CB�J=�N*9�rA^��]�q�R-k͝㮀�#0 6����g6P(2�H���3M	�cfc�uu [�@
q��(�e^ַ�A�{'���Ye�f.�H�������E�t�.��P8'_f3E���!N����I,ӹ�W�q��w]�9�Ht�tP
H<��V� �g�:�Y�ug�;�[�D����"�p}�����bY4�A)0 =�ࡇ ��Sj)�u��x/ZB��P(��#���}��Gi�;�%�δe�Wsy~�>�U�io�]w�h-kۚ�(4(rUx��{:�sΦ��� �S	�6Z�)e��l4l=��@K�٬�����^J�!Ť5�����@�(�y�)ӄ]���Bt<��(�����h~��ؾ��2�KK;��IOԆ�R�L�̿�� ƒ[����R�4I/;
��*��H� �	��Exh,-��3��r[�2:�pVd4#�aP0��h�0�fiG��w�~J��cG �UU��^S^���,����%m���i��Y�Q[�ɲ�mCɥ�?�7�o�W�\ ����uYc�Q�����}�Z�::��E�X*Y�2�P�T��"pr��'�Ώ�>G7DIE�#�.�j�ca�u�h��][Z*�r��BD}�:u��ܷ��Z%F-\�J�;O�3%����_�����������pnG��ŪT��ٶC+	��h�e��H��)T�7f�>��P�'������K��w킠�T=���a�;[��bU@ۚ5��[o	�t��3Q[��	J�%K"��_���2��Np����c-�!�*�����KU�����	a>u�a�b���{�ݸQh�*%��?JWQ6���>d��C)���<�$��w���������D��d�5�l���]+�^~��&b�fqc�d�>ܞ--%X�"�EO-�*h)A�q�������%:���~��jZG�)��1�`��A����=��E��
 W��WV4zS��9M��<k�HB�E�0�:w���TV�H���p7�%���.]��x:6n���^;42iD�9Bc�j�	u"so�9ArmD�4N+C@n���Hߗ��K��%2MM��k
&�v̀Ch[�R5�ٯ�&��+�@�
H�5�@����)S��k��Ic{�l����ara�1��3��7���م�;T�D��g��3��L--e
Z�7I�������$�]]`b݀	8�8/��m�p��a�7������;�D"N0�'O��?�
���,�Yx�?��իa�����{�Y���7E�����\/&�AA�
>��9�N��--`�Ҳ�U�c}��Wn�k*��c!x�y�a<:������:Yta,��.�h�u�ʕ��'w��y�>��g/��g�����w��c��s<���{��π|X���z�6�_�=={>�:�2��n���*�Ĩy�����	gc�Xtｎ�l߾���ӧ�_0�V���)�ӹ�з�#S�9?��'Zi��[)�-A��5
��J|�^(�
6S�W_�?���5����:5qH�ZU�#�[o���;�t�c,�9�޲~��{�:4�E�E�ob�~/��҆n
Z������믇�o����S�\�
�x�	hŴX�ʙ�#y�Y�8�l��tҕ_|���u�c�!�����She!�|���Ucq���b6�����A�׎jl��"T1M���`�����u�OkS��$
���,��ĈŋW����aG.�L�/�8����$������[�lT�����̯�us�Y���zOj�88��� ��W<����m�@FI	�W9�%�����8x�F zg'�,B��CsC���"13'%��䢮�Ј��Hn �t㧟����G�+d�&|�V@�?�D2�t �ʼO��< �k� 0��!l�`�9�1�� ��Z��$���(��*Q١{ 4����Z����lB.�E��g�����a����l�@�U�
���j،~�o����O�7FB{ ބ6�������6r�?�?���!���@V�X�ulN�`�۪|��Ѥ�_H٠{ $��>P��?-&(��}��m3ZWa/~������/�o��؜���fc��JFR?(侮��_��`s�ӀҬ_0��VQ@H���F~�����b{�?������B�5‐�A�3����!�(E^��%Y�D6 �F?���|���=7��dA/�$�ݦD�D��k4���K�����
�ŧc3��Uh�kH$)��0=�;����@���ө~w
󗏽[i��� �]\}%�>����C�&�� �m� < ��ȉ$����D2�H�"�T"��@$S�d*�LE ��D2�H�"�T"��@$S�d*�L�I�����\�    IEND�B`�PK
     t$v[9&��ސ ސ /   images/b01488b3-8551-4b4c-b09f-2812c4acc168.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  ��IDATx��y�m�Y��=�s����n�$�I��� �1���0(. U�D�	W���T��
�+�JR�#�B�Bʩr*�+�	6�6�hh���o���{�=��o\{�s�{��H�}��^����a���^��}���p8��N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p��h=��?���0>"�����0<�޿T�fS���bߔC�S��)�P��� ����e�C����0x`(gu��]� �(�X�_��y�����<�����:�=B�6�n���7�k���S�#�F�����S�1-0��!$�n<���!��`(���x~��'�����'�G�iX�s�q�8����:��q)v$7���GY4��1@�a�נ��?`�3��`�G1���3�����|��(��P�����ʢ⯥�(e#�]����eXq���8�W��&��n��g�^6���"t�����fq}�4��/������;�M8ٟ�瞀����O�(��p�$���yL��&�PA���-BꊠDO
����La(Z��g<�0Ȝ������I}"ţM-�I���\�C��x1D<���ؾ�,�"���U��_����>��W�7O��'��W�c7��－�y�������� R����g�H�7B$֌���fd�I���*��@�7%t2�}��|�W&��:	"!j�X�c$~���(�#l�bn:n��kuh�$���y,g~Y�����?o��oCc�F���YBY���c��pp��5�[Bo�^��|�vs'Oު7�/��>������?�R�UH�oA*|��Ȉ��;��0G��HDM��3	'}T�v:�lRO /o�g���q"�ٕ7���Zk��'�]�z�����>�=u�*Y���(��TAQ�ş�Y��+�>9����x��py�W���~z�Əݽ����!v_��Ư��T�8��:�e�����P��'mQfDr�^��L�l��0�Kll@��,�&���Mu�1$��َ'R��ь��ND[&�k_�Ch���{=m
��a�X>���D�.�-*Mź(ʋ0;x�<{aYՇЬϡ]�C}p"���w��.^䟛faqt\��_X޹���߆��N4���؟�l��)�u����	=z���S�(�a��<�ؓ	�I=�p{�|�\�b����d�X�]#y_¦_�r��
ϵCR�c�z��MQ�]�i�Ԋ�ҡ��B�d���U������>��!��������~���~i�6_��)��;��.�K��O"W�����ߌ���)��}w#v-���]�$oB!�3� �g]�0���zg�"Z�� +*�&�_
���D�7E,���dGeO>�<{�˘�b@��|�Z�->�	���2���3h��iQ�!��$��ֳ�����_����� ycI�8�u�X�7�N���g?K����N��=��au��hѾ?��si�n�^X��"7�B�L�=��T�t�2�ĉt�
�&�υ�)�moz�G�'���}�B�Y�MS��-��;G}	�8�[\�C? Q� ��hU�P��]ࢤ+ ����:̠�j<���&4q��0o�;��{����W~����?����O���_���p�Ʊ�l�B^-�����G��}ٛ�z�����}�M���[#-���S�dN2eM��@Y��q�o�U��	�D�!LB�&����׳+s*/�GCf"/���*���ҔD/(8�4�ʲck�,��>��~����
��?E�����^���������_trl/��ާ�Y��)Q�=�������8��Cw���+=� ;&Q
��ԍy��.T7�2�q͚�LD��1�<yF7�����~6�ϳw�>Ç�cH����Bo���*{�$�t}M۲�>�WpPԜ�W��y��Zz���",XC���� �1�z��_~���������o|ӗ���_ï�*@�� ���|�����c��ɧ��}�bx��x�[/����E���4ϴ�͢�܁�d>��B���OT��s�|������T{yޡ�� I=Q��š8LeQd<��s��)M��v`�<���Y��c��kfܐ�-J1�3=Z&(�Bq���1��W���Q��A�gB���a�������������z�w�m�\܆fyN�z���n	}u�.�G7`}����3T[ᤆ�����G���}�Z�5S�ؔ���i�T�2�坑�w�'#�4e��N�d�����Q���s:�l�����A��c��(���s�G�������5�����=���-|\C�⍞�u�x�u��妄��jg�c��?���4|?.�_/����o�\U�G��ߋo���!�m�bq�&8��?./ɥ8}xx���bh\��{��~�����v}�n�7�A���j������	�4x2RzT���e���8T�Q�D�/�EٱZCs8��CR��A1G%H��rb;��l�d	[ϛL�OL���А���E���/�}�(
s�� m��#��b�F$��*�j���gc,�������^J��1�Q�'/��Q?I���g f�NN��}��Ї����'��_V�_xk�^�N��}kHm�3�'�h�B��$nN�	�svy�y;2��K[�r������F�<�t��B�� l_�&��ߨ��]��ʱ�4��;�i�Z|o�E��P���z*_KhŇ�-��H�ҕP�ڢa�K���b����g��{CQ�VY��)��o�bY-u��Q8�AY�9�@�7����ڥ� 	7�>����n6'i迹o7�o��˴z[��<�6�e�������	z^)���G�60l6h��Tw��xǖ8���F?�Y�%�n�A�$�Y��s��4|���i4L�dː7b�g�C ��Kz_�qx�z�� �TbB9E5C%�������v��墨>Z��C��̓�%~�N�i뻟���m����S��$��K����@<8^\���7�����o}s�̆�eDm�Yr�h�V��G���K�ʄ5�dYm��YcM����!�v7M�8M��ɀ/�y
�&|O��k�U�Q�je��"f&U	��r�kv�G=�.UH��hS͵�TO�%��~#�E���))Ѯ/C�>���7T��+c5��b���P����Z�Z]U/���;�=��Ւ�+�����.U�5���
{���E1G���gp�[����a�~6���0���$^�+$�5��Hͮ�'�S\����f��ް�=�h��:4С�,��Sw��s�2�
K�� �x�2����4c���ו-{���L,�P�����Q~����N�1�8����$��
�����TTo��_L}�eU}b�����8T���'O\l���3Y�A؃d���_� �,��&4��A��g!��*RW�0�Q�S�Z�du)��u�gk��S�q)M����m��+�l���
$�d�v�ZP6�'V|B�.���Z���J�8U����)X����.�"zVf�R�D"�Ԅ��ǥ�0P(fhЮGB_�tX�(V]�Gl�B[?W_�ٷB��nS�ˡ]��jV}�(��P�m.���%
�ri����r8�]�..�Cc�������e��ě�Q`<>��������ƾY>74�[�YU�6�@"�e[��_Ė��+�=Z�d t��54���{�k��}�V�F���뇒������5k(�K��U�q��'Ƥ\<&��Ul"W/F�}�O^�Tc�e7K��*s���à�����!s��9�/�e��{YY*��G�}kY�~��_[����Vy��G�7�������?�g����˟�xYΟ���c�o2u�[ 6���:��Բ�(RBG�fR��g��6��h+OB�2��Ěφ�Y��^׺�ǔ�L�di��4���L�$|Mnw*���D�F���E�"'�pգG���"��H��S7������c��E�`SA[́lzS<VE㊦|�T�SE��[U�R=�J��M���P��7�v�X����r�D�s�������X8_�`9�K��-���m����OR�^?�L�>�$�o����Ϧ�����9.�%�힓l{%�8l�:O\���wQ���m��(�sȑ��{������oт/��·��K�P����#^!�%O2��v$�6�[y����^N��CN�R�~�=���
�gCk�X;�zM�KB�C�R�}a�8��q�}E,���B�+G��_��x�O���J���߇/��y�ʬ�����	QǊ�T׮~��6-���&���)W���Q�b	���q�	��p��P]�{+ήnQA�N���dr�4UR����̭��&�WRIZQ
i#Y�r=��]at�U 瘞C���v��.���E��GQ (�G��0��.�es���^��t=��~��$�7AW�	������������hj��)��Op!�A�	����⳱�s�֗\N����1G�5�hL��m/��"\\�`6;�cjGIM9�)��NZS�Ã�r*���5
D�o��G��J.iLI2x#E���H=��Fi�"SG�rhg�'b!U��"{)�K��(�|K��<���*���Z'
}	%h��%T�+��J!�!��KK�Z�75)Ih��4]`F*$��>pl�M3���1� ��nA���ֽ�3�:��v�SCGCU�ۋ{Э.��7Mz:����ͧ���w#�7����U���,���q�yG��� �w/G��m�����^�=y�^�	�������.=�A$s�)u����~J���.�%�'�P�D��c||�7$�')Yk�7��ŉ��ҵ�U�+�x�HO\�(M��>Q�ܩ�m��B���Oԭ���j�]�Q_�_�V��b�}�ŋ�?.Nn��o���]� �W�.}y���Ot��?Em�CH�i��^<�nٔAK4̪6�[<F������;1e8�~鉻
s&{&�4#}�b�*��	lY�y��j�LT��Ob�at3��9穓`\CC�*��Nϑb�%�コM#[�ȝhus�	+ 2�;�̡���Հ¹9�*q+�������f�~>���jTZ ���{|��Me��T���^@��Xӭ>����������"�#���>��~���o�!^`���?/�"h��N��-h%�o���p�f����};��ia�p�!A7����T��,J,����8���������3��JiV�+��j(b���yR�xW���*<Ӫ$������ U�D���Vt��X�&8�(�K��	L�ہ��}4eT���� E�Aˋ��S��L�'�n
�q M>���}@8�%4�X��8�ė1Ц�������!K�8�����#�@�%#�p�b��CH�Z���[�D��Et������OǛ_���m��%8΄�������
m�F)���(���X��e;	Ք�Q�����y6Yش6HK�y��vu�2hv�Ϋ�(��?��|G��Սjv����Ko��zG��[`�<�Fǭa�c��s)J���*���"�@�5$�~#�nlq��C74���$ �+�*P=���\�K�i%lG�[P�-*���ch0�([P|���l�	�4b�Qz{�;<�2OM�mgeU]�v����L�����0Ns������
c�R49B�U7<XI�2�4��������x������/7����۟��7�^ox���hKU}p��\�5��?����C�.�A\O�ՙTlEP�S&�MD^�,���gU��L��q�#���u��|�Ŵ)ô=�	b�;%i��x(��z��'V�P����WE9M�R��9��Pc	J$�|�K0�ǊZ�ThTs�[�V*L�����S��'7`�EBm���p��[�(����CYm����(6w�P�����S�� �t���(=5?8Y��@�n�$�i�:P�O.I���@{�T����gI���+��^vE������t��~��3����|3/�^�u3���F*��0�fժ�JT_�<8���}y������Ev�HA-K��Ʃ��yE�j��!�4�5��B�d��%]���i �<��YJdr	����F�sx��-I�Q �E���j}F�ވ�2����.=��.��=N)���+���ŀ����ZS�d��P}�Cw��g��l��lx�?��Ռl�A�][�����csA��k0y���{.m���E�0L-�c�ln��uwq����@B��r�Z�7qt���i�c$��YH}U��H�MV�X��!b�M�"o��K-y۰E^�0�͆Ƥ����mN�|O�z�r�<{sHq�{N��z���<���th�]���b���J��Ē���s�˱u��EӺu�-o�O�{���4d%+�B�%�E��vgҤ�|ҿU�/V����-4qP�B"7e��!?���U��74է._�$?�fx=�5K�tcW�}HV�Yt�����8C߀��,����5�g�O #tB��'V�ul掹jLf��>���.E�>��t�M�&�������QH���ļe��r�6�
�Q[>D">��9#�flٍ�;�%�v�,j��1�GKl)8��-�9����dk��Q��l������([3�W������v=J���k���`���;*!)��)2��Z%�u�h䆢���] ��~��ۣ5CjyOk�%�p��ف����ʒCd̗����"�Ч�bٔ�.6Ų�l���k˾k��l�ȁ6d�H�&Uz��"�21�j���z��I��J�t���xYx���w��x�B�4��l���ob�?�d3�?�<4����s}����(��'ǹx��5yTe��R��s.�K(.聆9#�;[^�ǁ�5ȓӓM%͐X��yE���Ef�ܴ�<=����0Q2%:j��s�A��@�'T�-B�J~��N��ZU���J�ޢ^�Rg�70�ȑ/-g�8$�\�x�^W��ѲB�'jr�5(p�0�RoFT�bI���X�{����(�ltD�W�V�W͠���kMu�%-��#B_�E���]���g�ZVG��X�ְF�=���C�A�_�Vܧ��,}���9��H�u͊� .�S�t>��}]��NaDjޠ�49�Fu2���&��4�Iq6Y��ibq���ۖ�p��gV����s�$���-��2~�䉪>�ţ�����۟�q���o��^��~�����p���?�ͱo~.��/A���Nz�v���g0�1h�7+	��;������?u�g��>:���6�uu_7k}"6���|��C��,a/���F�Q��g�`���:	�����2Ֆ�G�u�J�2d%s8U2�q�R}z��Y��G6�uZº?��>�cΔ� @��)ǥHj����\Z�P���λ/�%�$E�=�Fu����b�V�*��`=����B�r/ǛJ"v�[�Ҭ:8�����{�Xb�s\?�h�[�鉧C�FAn�U���8�7��"eU5̩�.�nG�pX6<�7�5{�c���`R��G%1O33�A����{LЎm�E�~d������Lb�8����\B����v�g�i2�3�HF$}����1e_Ǎx���	I�<���k�y�(g8��8<"��<�y�1 �I܂v.��c"�w����KRmjua�d)����L�)�6�ԇ��ј��A�I�.����������V=��q-�R��zb�ʥ�jΉ�I���y{r���GŊ��΁C�(�ig>-y���]��;e��\�:�~p�fu�2�����i�DR���
�x�2�*y�E��bY�t�87��jr@�l��"��UPi`v5���x2�M�=~%*�ܶ�G��,�8��ʃ��u��CC(���?�w�N҇/�K8��'�����k�YB?��8{����L]��C�|'��L�"(8�&%jZ�6�Z�I	r��u��f��<�B�j�$�C��]w�|턩sm�������7����ط6�2�(�L�L.qd���:�*�P��d˛�v�GV�y'���=�2%������hL��!��(#�f)� �N�0E�6�,o�&`�{�W��G�����x�D�J]&l�d[ઔM<%��� ɉ}�*���� �h�������8�'NR�y�)o�	d� �h��o襱�0��)q�
���0��f�r��Ǆ\%�����vϓv�ں��oד�u�J�L�{g>�Jҕ#Q~�6��X����y �q�BB.`J�L�ڈ�:�u�ذZP3�R"!k��p��Ť�1�2�#��<~�bmr�&��8�e;�n�+�ΪL�ۆ�*d��*�kR�C�
�������Z�c�N�?)�9��>������	b�2M���i�6�߆L�����$I�a��A����;�CCV���%,p<o�AlDAExݒ��Ĺ�"���&��h���y�D��d�o��ɍQ�]ޯ-����0����Q�C��U&�.��Iw��-dW9I��_yi�e#��0Gq��������+��#��C��?Ã?7�y���$���6\����=�u��5t���~�+����nZ��y����!7]fi����u��!+����ֻ>l�),aG�ؙ`�<oBhT.$l]�8)IB��9�}� �������vr�L���g�8	���X�d�r����Nr��Җ�k|�vu�mZ˨J���lM���}��vT� �$&�tY`�.zV���UL�)1+@�!��Uכ�|�����|)$5��0h<�h��!������Ȥ�K̙ȹl��9�n���:��,��+A�0�2�HH��P�<�u��<)��nv2a��3ӕ�9�.�_}�x�т��)�۱F��.��Iց(�EI7�7Z��
u�KTA�6�UC�=��� �y��Y�cR���2�6��7�f��%�ާ���9.u$J؜@�
�h�$>>%0����ш�5mLĥ���L�ٚv�?��37�ƍ!���5��O��}�9{?)�z�$L1���B�A�Y�Y�4�1�5)U�;0���\o�
E��>�آDc¢��������̲mQY��@e�I�^>�y��QǮ���#������&H[�����<�V��g��D�b��0=W>Q�#~��C�����-";�Θz�UF�KF�!��ή���s�O�{p����~�f��{�����=88}^�x�:�(��w�C���ط5vm�xs��\�����Iv����4G1���mR����#׶j��aO?��8Q�h�{����p�b9���W���fVi0˗��Iɐ��%���Y�|�<N��PE�s�Rd_�T���-WH�����K�����P`��	���/ �4ٶK�H�E�{�QY�1�@Vq �HQj���+��� �|�t(m��k^֯_H�v�����
�yݣ$���:�wڵq��,IXr��ĻSq}o�jr�Ib�t�d�(<gh�6�@���*H'%,��%]c�O��qlǡ	ݬ��3��ᔼ��:���f�lW��9�M��ǆ{T:��+J$�}䡠d#$�yGLJ`�~��$v�:Eb*��(�q]s~G�]��2�{$�~]�d�n��/D�`y�doX&����׷eM���"0�$m2���a�l.�4~?���]	Ƶ�Q� ��Х�T<@��`
}��<����2��Η�}��#��u���z�U�=�K$���ƷCI��0����`���q��YwR�T	�J�I�@9�����DCi:�Lw���ԟ4Z�F���`��'�w���?��(�ā����4E�����<0F�9��e�)o �9��bhP��,����N�������S�-\�{�_�h^s�~��'䗪|��=��FR���9���K�XdWyT!i�y�u���}��'�իߝL�f������P���t�B�d�T�C~�]C~~!���S���ݎ���=�ɽ{��c�x�cB�7P�%;p��ě����k�E����s<�,����I��}�ǭ���6��|-�`�VJQU��r^B)K� ��qU�`u�I�ˋP�n�D�Z0z��0�:+�]?�}� ���]l��͠��������.��;AÀ��J�`�I�pE�>�"�{{�ٮ`�lН�����;�V��Im���y�7ޜ�i�ز�NpK�n��晓�se~eRR�@���&B�F)�� �p��F��T)����LHj����x��B��ۥ*�B8�^ݓ�D�³�A�`���{$�ް`'��f|�d�R�!�.�/�Jr*f8�G|CJ�)Q.T�F�0��q�ړ�7{�tM�ˣ���[G�*#9��ǁJjTdC#��$f�\�Z���n��%��>*	��wI#oܜ�Y� jؑ��*�EI�B�����~]!7�\m�K�-����oI��кR��G!wAE���ْ���e/�$Ĩ�y|�
�K���$1EP�sZ^�Ī.t���JGCP���Vu�����`
��+�,s0�m�\��s��c��3ߏ�NGd/N���P�)����,�_�����?�6��x��5E�ͽ�x��>׵���������Nd�Tj2��%id���T1J5~���
F�hIJ�����,[J��Z�8
L����M6�r"��%��k޲��T( 'k���#Yδ�6)]+�})*�x��+=_�Z��,x]l��IL#�r�_@�c��ڈ�����ńD@��d��b&��"lT�l5�R�/���c����T��O��d4��c�(��Y36x�{R�B=	�_1��!˞c���7�&�Q>=���f�ӸQ)$�"h�����ɅD�Q]�����Ċ!9���R��f�U�T�;���z�Y��;{��Ė�iĪ�R4�%_�xL�{=G�b4�F6��*�T�T���D�;ϱA�օPeO��X ��G�b��B٢`�)y����-TցK�&L��57[@���0�D��I>��N�Y����4��n;�q��_�,k[yT$�l����MB�1�_?M�5�a:m�&:�������R�d]!+���Fj�ˊwQ;;;��2ޣS]��^�ry�M����1��������m�u�� E���7
+u�(�h���9j�<+w,K��8?�B[�Oy�<s�^ks�5>yЕ8'cc�%������a/�:���<`	���l�S�����t��i��-����q.�7���u'��2�'_{���f�nD{�e�f��zy�7�n��}Sp�����c�w�z��MsY��MH��hxbL,��X�8fB�>'G�J�c�2�V�D��1̮��v��Ӟ�q��4u��B m���^k� �[r��SsM�E�D ��z�->�	-�ܩ|"���8�nJS���,��{N�+E�%�fn9I���P�`v���s����������I������4�Z)��M���}�������tTW/)7d��TaP-s�,sj��콒$"���(�%O�E�DN�&�����%Jee�x'�|ÄP'�G�U�{����X�%K����O���)����tUm% �͓����=�<_�$9����=�2@B)��0���m��n���B�����Q�M���$e�v��4��C��^�($a�/vyvY֮ t�lO���{�	�#�&I�N	����z��k�pDi����.�CMbp�+~����I!-�8�k;RH�H�TvF�c�a�4�|R~����@�����8�/��]�?kT.���v�H��������۬��S�zY��^��&����DS���|�܃�(&.x́���)��c���C�=7@��c�8�01�tE�Q^�g�r ��is�K�Gp��������b�����^��zp�f���o���� �͇n���l�Z�nȚr��e���(���M��Td빘X��\��DI;�6�ѻ#�sc��l>=�}����������Y��.+U�j��s�09�-�(d��(�rW<�a���@��VzB!Q��~�%5����s����V1(~�wgܣ��ϵ�!7�$���4�萳�U�N�����o0m];ř�`2�\�+{O	1G���H�G��a���$@Tb��J�8���bΨMb�Df� DRP��Vt-�?ML�R#�O��j!��-�o�����t��U1�٠36k��r�10�%�`����kdKx�8�(㼘(SI�N�:�dd��#�LÐO��f���Wa�?�4��#�QY�<�()	���ce�TE��5���d������\��!�I�l��%�I~�����X�۩I��\�@�_1Fr�!Q�>�����\S~y�����*[W'&�җ���6��#�w�����j.�a1�s��r����c���]=���Է�($�Y���mzQ�Ed<���`�J�G;��4giz,;�Ȍ�呻�}<���J���HBoAs�ݖ�)1��`�n��R�F�5�h��#�!\���ǎ�^���p�����ٷ�k�:���w��\܇/������Y�x�g(�F��ҌAk�q�s�{!�s���X� �$�]�*��t���D����^����f�I�qb�G��t�Ԯ$t���&��������[=�vۇ4�,`V�udbˍ]TI[В˽�ul�Ak��]-�k)�T�f-�,�I��� ��X�n6Ht�l�*ۻ��a��X�`��Ⓡ�'j)bN��C�R;kA� �5[#�5j�^�GU��yǥ)m��
Y�I��iY8[7<NG�^tb�S���%����(�@�f+%p5mtC�XQ��`�QJX6?�߶��D��57�LR!mϡ�0h9
S���jc!�dR`'
���S~g&�a!W�tb1S,���Cz��Ф�ˬfR[]�|��<����v�N�<!�M�I�6W���Uyͅ��!_��r�ZW��b���I=�)�Y��N�y��:c�rS�t�ɱsK�k�@��g״�W6^�A\�F�D�k$݊���Y��Q{גI�Y�q�%����!�z��BR��з=,GLt]��K<�j�\ӆ.��o6|�y�dx�뮥nN�qx����ֺ�~�I�*Iv<�����!��v^7OȘ�d�J�@T�9d���C�ׂ(�A�6�{Xv^l�g��&ޫ��w�ò�T�x�p�̛ᵀW����/����E�'o���?>��o�\��ɎBd�s�$�q7�(�7qU����Z����	 �I�:�^���0�|��ڼ�xcn�|�te-\�I��+�8�K��
"tr����ރ�8�~��2Liܖ5��!M��T5W��%���h���!�����QM*w�Ӥ;w+��3N����	mbB��]����l��h�Pn��G/~G���[-]c��>���bΖ��:\P�{����4P��>�$��Bզ�1���Y������e;�>�Y���\u'�Q)נ��8��+������ܘ$5U?mNZhŬ�Qh���Y�[����?m}l��f����x*A��!���D�Ĳ�8ւx�U��L�)�1k�@)��FY��j�
Mw3�I��3�j�y�-C5*�3�&��L����`� l��0,��d/���'�S��Q�7��}O����w�LTe��S�y�͎P�#b��K"qT47���T�V��.���	�ᙧ��'��{w���y�՚�?O{�d��B��:�i�z��3���Y���.���d|�qMoW�����7���'�P��jχIb��3��d�e��њt-��dI��/5�81�?Eq�.>�o��2~�����o�O=w��[x��w���W�Щ��ʃ�o��woo���o7({�}&�ȍĥ�V]�Qj����8��,�rm�X
�\����Jj=9d�i2�¨�e�|2�R��_�l��oyH��X�K`�m�N� mX+&s\�x=U�r�<%�����%�e�_���(��L�n�8���5��%�[6j�V�D�ԝE�QR&�1�M��#��"���P�7meK���v-��ɯ�ތ�}�ݖ�7����Ę,f&_3��������"'XQ�{ ��A�=c�-I�q�2@�޷�\I�Z�=
W*]�{��-
�
')�P�6��(�Fʯ�-
ZY1�����3Q~䦎��}�rL��5�ig�yQ�[bʅ�-��5����g/j���9�e��鐅ɒLXN�
<�Dh*��v=��(�$S����[���EU`Ұ��?l��y�Dɥ�1���b�rh�s���g����QT���є�`zOG%i*���J`r���[a�MY����P�fL�D����pr�&Z�K� 97�l��ԭ[h ��Z�=����3���{���.��p�\q%G�JYŜhG����RhF�6Y��ES���>[÷c͇��c�<
���d��=��M16��{�c*��c?���`��Q��Be�$5<l>s� y�Iߧ�L
�7D����������'O��^x-�U#tv�o������m_�5_��RO;�Q�f'�M��7�NpA��<���G��jN�R35�tڈ�Z��L[�����/�V-{\C����[�����ld���Z̠;D��s\"i�����O��UD"/�he�`1H�N���UQ�1�'�&�c�A2ԣ.�a����%Bt�lQ������aɄ^R�
7��x�k�AA���Q�(���ZT7����\qY���e�"@�ՓUGJB�V5�)&������1�3��I����T�D Q-�������J��VT��������ٔ %4od�W�jz��M��,xR��ͥ�~@W�O���x�m�C���%}'=�A�������*ق��mL�]�Ģ+����2��Z)��YK�y�=-��X�h�&��������F\�4	!XPG<�O�X�k��LjB��vO��(�<`�-�9�ӝ����)A�[����\FK��4����� '�qITUq"�Q`	�A��҂��ě�|mZfv�c5���1O����w�2�]fǯi�Q���笔�=�s�5���8V䵛�`�cՓ!T8�y������§>����wh�p��!\\&h.py)�>��q�KN�f�a��=��������~�%嫝3�D9c���O�	J3����M)��@!�v0�WY1���i����@%�*��}���j�76�O�Y�_^<��Η�=�x5�Z�;/�;������b���D���v��`z%���C��'��\���8Y�r��(�f3J�#��Qdd�2Y�-�h;NH�W��f"��=�	�+���6&�lZ4�q_!�N.p�Bk�B�po렞�$q�a����$�ʽ��I��uAP"_�;IR;���%4�x9l���P���v�@��%o�BǓ$2�(H�uM��cCj�e�m��kzKpduJ�a����L���&&�F��%J���-�M���v��ڴ�EU�L&tRU�8[���H������*o()Ǩ����#nI���\$8[Gh��̯�cu��i&�:��X�ZrBT�\��m�e�F�+3FF�ºB�cP�5E�@�Y<�kŕ�'��{v�Ǚ䮔��{����9�y9Ve�=D��7|��E/)Q8��+�y��l�'�QJ�����c���L}f�!L��S���2P'@�܃�ʥ��p-��(�SE 4AQ��wjmZ������$���������td�^�8��
��^�g��R�d�/8�������{د.���I|����x3�Z�4��,�ʻe�cA��HS���:똃���7k�����k�V�֘e�H楄3��Ys��cE�$�a?U��y6Ie����ݑykk#��p��S�Ǔ�\J�Ѐ���*�G��-��O�x�/��w���pt�Yx��zsvNN�~�� N��uH}#��P��h1r}�F���8�}�s`����Q_�w	�Ɠ�'�����p�[JȵưM#4!�b�[�����F�B�R�7� j����L��6)�2y��UKB���5��� �orC?�|-�5�)�v;�C��5[�}�HW5�4�-yG�4"9�5�lr6�kK��H_	a���&�D�a�5,����B�Z��m�v��1}�Ĺ6u<�en@$��ErCJ�m��jVHz.]��I��8��cŊj�_:kᅳ _zZ���E�q�z�t�/�UO��7����2w= 0n���jb\���|DZh��-JAR��֪d��G�G��[�!}"�.���$;���95H�L$|���������k!��S偽7Ɖ�l�p��8�2 g�ш��5��nZ����$�ܒ���~����nP�=7˱n��a>/y�ɻq�8�c��ɫ� ɯ�+���a�����{�����P�A��ީ�%XR�=��R(1fz"�
]I��Gͫ��Z��>okc+7��q]O����ŭs�[�%�Pb������W0S�Q�x���~�o����'�O��77˗�o�1� �^B盱�B�9{��.�o�7c'�9��i)����Jyw���V�FBFw�#0�~�q��ݷ^)B��M�T�Oj�(��7���T �h����Y �WJ��h}�E�Y9���
s�r�`��	��� 	.I�<m�B�z��*�|��`6�Z�Գ�w>��ۈuS��{A�|�E�F7t�^uɤ�4�
&�^]-f$����ȵ'q�f�(j�M���7!��J�B���Υ�!R5�^E'�Uڝ��������iܼ��2�^z�����}�n�"'lKD�g����2���``ۮ�G����5�$����1L��
6�7���8�M����/�t��9���lߛ��R�V�J�R�/����"����(��܈֧ݮ!f��zy��B��غ��eO\�$�Uz>�M����څI�O=OI��^&�����[��N��� JIp�g=���f�
NN��`�d^�ť�w@��е�T�6dE�&��b��_��h`�l��ym��� smnM����d�sK��9�۝���������5����W@KC9	���310���"c̰�r�Ʀ%�E���J}�U�Uku�S�|��?���~�s�j�N���]��>K5̧(x�߬�<�:[���9��d�jKCޓ{�^����7QmL,�.Fbe�MҰ�x�+o`��R��8=�� ?�g�w�W VhT�膤wS�5�$K&I�iސ���9W��.b����ӽZb�e�b˴�e�#Gv'M��K�:ơ��s)��삋��Ye���Y��uÊ��p�tL��J��y���Dr��ܥ��d-��Z�K�;�d��F��j������0�OJ]8E3Yon��q׾P�yW��(\�o��O$fg
�e�@�m��v��~5��h�
�]�`�����&!A����JMi�Z,tS��Q�n[2_C�X��e�=|��4��1����⍽z6L����#Xמɸ�\����Ҵ�_S(&��C>.�<�sV� _��� �W�=�&vlK㧍@�gcYƿ�9���1�
��LZ[k$�7�+�-o
!=��㰘��Y<�ٽ�R�f15�w�`��o>�a�Y絜� ��\P�6<B>JF~�y���^Qv��;߷�I����5z*���VVԜ�2��B,�>I�d�=��Fϱ(�]�C��R?����ֿ���\��=_�M\����߮��ˢ]/x蚿�7���mX���ZXw?b�,��d�=\nA.@�`$B$׹�G�\ՌU�]gAoY1��)��?�zVi`���e����R7��w!���F�t,g�X� �	iyS9�� �z�`�B�]�TW�}�E�������Jv"���8�t���s�%�4He|��D��yC�$�,�Y�W@ز�L��b3����
d��`�2oՆ#�/fg�{�Ƌ��8�4�D����,�l�XJb��Ś�X�i k�K�vڃ��3xжp�V��&�WD���5V�5�xW��Cf���ˎ�%@�H,�ŻA���Nj5�2�˅D-K�d:Sd�e��}[����{�P��M�A�zK�"[^V�8Q�lL���9���Zq��;M��Q1�މ1�vW}�q�5u�5�M�� ��=����=9fP�6D����w�w�	���)�Ԝ�m������'�C��%~��jV��Bߺ����{3,�h �ӎm�Iߴ�����D�Ъ�]��E�:O��t,�*�Y1�fM<��d��f/%+!��^J�r"��� &���5�ZE~S�]��șh.w�o$;���M�cE9�����W��V���?;|A	����7��+a6?��]��Y>N��ҾɺI'[�)�֨bK�BIE� 6���Y�[Hٕ9�Y�	Q�R��mvZA�א����i�^���n�3)с�C����DpqM�$i�媺��ؔ��dRW�-��I�u)[��ЙЭ_�N��]R��.uqXs�$MBt���*ĬJC�w���7�'�\�㉘b ������A�D�f1+� ���Ж���bҽ�)9���&���b�Iw��)f��'*g	��W�]�pѯڄ�v�Ǽ
땐���lܵ��<rz>z�N��e��Io��22�;z�;��=��u3
g���[�׺J�����>�"(9!e.5��q���Q�*��[�f������k���My׫�Z�6'caT&s:�T����7(��|�jS�y2�('.xs[v�g/����
��bG'��#i�~�ʣtB�F<5�[3�..a���=��S\gN��ٽy'�'N��=�,8==�^�FZA���p��1�+��	����d{�\�&��^����Vr�����+%6M����ż�ܹQ����s��8��,T�q�GjPV%{�����>�۱��Aw���܊Ο=�`��>?�A��^��'C�~>D�s1u��7,�j�LV	b�V$�/)j@�.A�����`$�m-������B���y����W������B��ꦁ||�V��GGv��Y��Fi�ܩ�O��2�M��g�'�&)����ִ�]�T�ɼ��7m�J�mM�`�voE)t���D�����nd��5O}M�U��h'�<g�j"|�u��FO��_���Kq�L����ͪ���~"̙��$�
*y����8&��"��Q2� ٤fVע0tH�\Y �O5H�ڑ���6��yr�u�ǧ�E�T��0q7�5��O:)eK]U��9>��޾�z�$.֬�ۢ��k���5��%��!RzO%瘃�:W��k�֯��A�%:$�G�'�v��C��{-+U�,���q�U���my�;��߯S��ؓ�ܾ�w�J�A� "_��>�
�ɯ�s��K �1i�
��25�s�|�V���N�H/���baW|�e�{�̏P� ��/pXpY��l��U\��� �����Pq�Uڿ��R�k���ԃ�L�������mu����2�?���J[1�Za�'��Jr8�\$�p�y���H+�,TN�ᨖy*R�\�;\Փ t�,H3�����ۼ�o�-g?�V��yo~z
_(|A�k��(@������6�ݱojj#)�C�G���	���ٹC\��9�eM%�����ė�T��4�['%��Xr����c���[��M�W�9d�`�����抓�"�Zgk4e��(`P� L�)�ߣ�1��&����d�S��
� Tiꓩ�6�����k��6*�};.$�.¤5�J6��R��JB��5*=�6��v�|�Il�ܠ���}��yF�\$�g��u�㺃YAЈ�*�</Q;k=
�V��ӆ+������Q2��h�T����-슊
)�Qq9�f���D��Z
|��엲���x�"ߚ�6S��+��0��ʓ����
��Ne/}��,Gj�K%e�Pi+YY���d��[�k/��O�[�&�?��i�YҤx���AjV@���E�	�����Ī��xt�,�q��m��.�O���#v~�]��\������"ϋo� ���k=iR�y���pl�ĭ^c!q񪬳\x��Gp��-�=u�\5��ڼ\�f.}+��G��ʧ�D2�����qP'�ڔMf���Q�޿�������k�h,#��lyu����'
jV�B���f�Dm�
�*�*5x��۝;�C<HR���x���>�+*y�0/M�p+�Q&L�~���z�7�����������i�����З�_�yw���OR��t��J����	]���i�&s���?�Ŏ]����.�	�o�g4Ɍ�����N"u���ͳ�29N>^'�Ð�n�ט�	{�)�SD��,K.���hЉ�GڧE������\��r�*y�t��C�lx����zr���U��_����bw��������ըoG���j҇5�:
L�fJ�uϊ�.֔욖x�w�;+��%g�����$q�8.�`����� �^�����>�H�?u��`���h�L.�d�G�,9�}�~[� �[�+��|)�Ňg8.sn�kQ�	����c�,?�L0W�Z�Q��H�5�G���S���G�C�Tyz�enϧ�u_��re.��}-Wb�3� 6B��c��#���� ���|~]����͛�m�۩.Jj庀�>��x�e�g��g�>����Ƃ�"Q�Z��y�PE����5m�u߄�2��M��'�}u<��e�ݞ7�Q׍�f('�'a���޺?I� ��e�
�;%ҽ�R�ް�j0�@U�+jo�BwL�
k�-�&��6�\�[,� U��{�;��o�/߇/>yp6�w����S}���خރ��[�Z�݈Ƹ9g>�eHY�-�=�7�)]�l�&�.!�4ɴ�^d[�G�u!��Ab�����Ʉy���nPS��/��c-9͍����^��kRO-�:��7ߦ�,�YE-�Ӗ�X�%u��������v�c;�)1�'n^!�ȅd��wǥB�\&l���Ucۥ+c&��B�t[���fz�-�v�ޟ1S<�X��M�t�EA�čt8Ӏ,sj&�.*�!��G{r%%���RuA-�QXPc���A?���N@���޷e�?I'�2.�>+Y��w�I=deI�ħd��)E{��Wf=p�y�����1Z���s�Q����i��@7M2덟S�ݒ�)�����~���Rj)AQs�NC�Ӷux}B�u��+�r�q��W��%� 3�ާ��{1Q�g�1�l6���S8����//6��@�s"*�(��n@�@����-$����N��E���1�y���5u>��:ٟ�6	�U����z��l��0�E>�=6~!+}��NtJ�ZJ&�V4�}ˊߞ��S�>M��i�3i�6�(�v:�0�9J����l�I	�)Q,�PH;eRBe��5�3�;�凊�����c�m._�����������4H���tެ����.�J��,b+{�Ԣm1i;2iB[��5��|��F�m?X�%�+Y��D���C��n�V��qn�kH�:�ݴg��191X&1�d
ŤDm��0j��ʠ�\��;$�%���)�Ei=��-��ص�m-So� �~�~�o9k�Hb� j
���]`B�=7[�V�&�3�a�����K|�V�uu�E&W������S����cS�<�<M�A��x�s"ur�i�R�PgŪ{К�pQ���-���a�1e5sC-Q�K� ���G���X��u�3>�p�I*�Fg2=F(]���Bھ��q��9�X?�q��ǿ(�2�ę3�r���&��6��p��v^��a!����g�'W��z��y�by]��nb�+��QK�aHJX�6�)��Vб�(�3T(G5�Pt�>*_�f�!%<v���|
���H%n�wy��3��U04�,����@�P]�}��r*T��v�����{f.E9�+s�����'d�h�)~i*���!�,�Y����c�E1GB�>�A1���o�I�5v�g�G<J�;��εC�a�7e��+����'��v����z��z�\�3?�볗�v�ڿ�oV7c��d�iQ,\݀%��>���F�����Z�$<��c�nJ���Y %\�qڍ���B)�1�ʎQ�u��j���D��:(�O��>*x�#%�¦s�꒝�QM�n`�.�I�Y�gy^��(=�Ţ�ms+�$�`�#W�}ZpB�ԄG%�"9�Js�b�m�9�{ ݞvz�����l�̇[@��:�J'��}�>l_f���y0]�����g�#�j�������}�%NJm39���#�;]].�J��
Y&d�RNӒ�"�>���:�"]���u��ļ4ꉹ����&�8�����G������,`Io����QP[�#�r�r�X�R�'���%�T��)����v��Q�񑐷�aK1���n���&�]"�
��הG҈������V�����T*q���^�Q��I��QJ�+��XN���]]Wp���a����K�Z���vg�
�K�G�5`��1oDĝ���!�~���Z9I��W�"�v݅���V�{-f�|bi�c���� �����x!}�֕ +p�x���mu.�B�&[�Vѡ�
"��̶(
5Ri����V�?���_���~�fu��x��������i87�α��h���з_ie�����s��\wXz�Ķ-W�J��Q�y����}_C�y���Z��H�8Y�6�f&���˙���da�
��s���2��S�`\�I�=��$I(��B밂U���A����3�jId��6R��>hֶ�֔`{��-� �h%��Q��'� G�"\7��)5��M:�!>J L?ÉA�|n�h�.4S�̃!���p��JmH�dT�8�90� �E�V#��ą�(���yAU�7:��I�[ɂ7 ��r�Q+>��Xm�!!��,�_�� ���[�}�C~�k�:K�s�5���CĞ
Ʉ�.M��H���Z�Ie$�[P���;,��T �"�6�&��(k�Qޝ1������:���*���6},�I��c
��\s�#n�[�V����8<>��%	�����/kr��PłyX!��ap����T� �d��|t졛�+VVc'�[�S�MFXZ���m�n�n�C&W�ǳ=/,*����#q��{���D��2U� �*�p�o����HZ��N'y:�U��$�����bQ侢����q㙏w�;/�N�y�g���B��l�8�<j���f�]�݄����n��m[zP�}��2�\����s�JY!�,�HDDL�5�
�1JIb�D_�<��� �)�A0��/�!���*����9���֚�K���k����?�Z{�S�����s����/�����F��V��t��ˋ"�A#�"���鑹,��`�̈́�[���5��������B��x�_�z�Ν���|�	�l��([�"��mܒ�5g&��1�f�S&a����_RQ�<�����l5O��؟;�vW~߇�٣�n�;�)�+� F��^`��T�h�=��Z�&Ώ_M��^�����_Rз8t�G҆*�mc$����&4/����^�eD@�h����.jW����%�	�� �ѺJ"Zsƹ�o��]�4�De��V:݀�-�?Gk�"T����6y͗�`���Gl([���\��*�B����=�����~���:~�P�=��FӨ���V�W�B���ԁCa$e%�aj'XU	��U14D1���7�o�p/���#�%l��Go^��ڝ���F�H��Q���t�TP�O�F��/�"���t���h���F#�J�� ���Wo�p�Z�23ʴ�O���s_U��P,l�$Z=��}�WD�u-���Gn�Mw2��yvs>�mn�"�}���_�_=d7�]�WFțu����ϑ?�^5�d��0_�ޡ�es��)j�3ݨ�>(��K#ǳd�D�3`m>��)$�HT�V��ΒH�-��^�"��~|������������*�]�o�B������]�@�?|�����_���ﱰ4W�� jq׼(N�E�Y���̳*`���*��m1��*:T�
dw��gIQ@����ș�ur��.�"�TK�L�g�^+Y���S�Yy�r��	�!73P��q�o�[�MY�,��N�^�*�8�ŭ�v,@X�c��>�5QAU#�U���Z��ރ���š	j�Q��
�&�tcg�:Z?8j?ۚ�O���M\P���M(4�� )>X�:R�*�ܽ�F_�����c�vV�MiOh���J�v2��q̨���#�246��L&P�����6�$B��a�9�vC��4,e����=[Ӯ�B������|��{on �J����\�2�^�h:�C���Y�綞'+"�����b=9� S�^m!8�,=��� ��ת}Đ5_1�V���L����v���LD��se����^Id��^8�Љ�\��ֺ�y�M�����tu*T�iȑ뱚�x{~�PFQ������Ⱦr�e���ʔy�/
����u��{a�D�ߊ�����f����ve�޾���\<�(G �޾�<�b8==�W/��U�z�F�W���x�z�5-���ES��!��m��|,Z�{�ϛ�����&��!J]e�+y�׈�hx�]��8w��c���
%�\�c��5��]Y���P�����iz5��O_�~�W�?����{���o��SW�K�������/��ߙ/����R���3�7�ޔ 9Zz��zG�ඉ}���?��-�[�p�G�Q�w�& Q��<Y��Xt`F7��z���b (�ZS�@3��j�m�>�/4����ۧ����ůy���A��O���=R��ٵ: ������(.2h[tC���{�gI��X����R�#O���v���?:�.�7:�:��G6zv���E����X��5mg�k�>SV8f��E�=h`x�y�2�	t����vʙldΓd?�#"���z?^�6�Q�эk?&��@�E���Mݷ���;0��~�*�J�%��T���'%
�R�m䳃��d��1M�y:t����~�Zm����O.ج���ѱ�3n�B��k���	UrC}���=J�1�}[E�-���{I�Î�	E���E�V���uAWCx�b��(�o�J���ûw����������׋vYC�1z:�z������|��ƛ���z�����M��n��V����qQ��
;��#X��6��:I�y��B�-K�o1���嫿�k�����߿���@8�SU��E�b��:������r}�̝[��܅�k�}1���ҼUe�F��& �WK��׷�z�2�|�/�����;�ë�)��ټR��x���k��My�R�!6����#ú)Ѫ
~�ho�G�A(�zz�t���$��˸�!� ��Hκ�RC�4ԑ��}Ԯ^��T^�jJ��Ew�w��+(K��kZ��L��*��պ��7�$����@���?l���[��\�^�� �Δ��Z��j�g��^"6}� %��QI��45��}?0���:�1��-�y��d����q�۵�\	���Oϕ��zG��j���uI���^ڌ��Τ���e���A��OƓ�C���Y]u�S;oto*��B��ί1XJg�d���ߎ�����Ɔ�����i�G�KΝ<�11����=r����X3x��:}�x6���u���o�%����(E��(��PN{���=P3{ʾ��Fˣ����ʚF��3ӵx��� ����_��*E�5��,��g��=�*���֢%_�O�����q'��uq���ֶ�A�Q��[�I#�̅F�*̋7p6���	F�$�D&�5���0��y���X���oǽ��:e���)���տ�L�j�>�3؞�����|���eQ�y2��W�����j�ӲP� Ǣ�K�	ia �RʂF��p|�J��3��<�R��Y?_d�슥��D�e�a�bļ��{jA�\7w0���k����s� &�Q��~-�I�C/j�x�E�>�P61�i(q�ﾐ�fDn�^B���E=Kg8�|%�v,�j���^z4�'U {�+����^��N���r?v�|��~�c���"��"�n��]{�k`��!wc/ÞܱEj��[�������g�/�t_�6a'Y1�1����ӱr%ͼ|����qS�^(f/c��hG��U��y�ݼ��a�n��h7��^��n�
��
�j�f�k0"+g�5���xM�%R����y�0��>����_��b�X���k�n��m���x�9�˽��qel�M���wX5Nξ��zd1��q@eBGE�j�B�\ �
��G��OS��4�e-fI�ā������2���y^}V���<͗`,�Z�ʆC��՚^}�u�v�.ݙ�]4��V�	���Q��6��'��%�%�������Dr0�-���4R�`�"���i�?��|��v�ǿ:��/M�~ ��?�S�����~��o�ݛo��e�������4=�}{��������
|[<0�B/
	 ��V�3������;�t�,�l�╏P臷���J�{�M&0���T�%��f���z��az��ɽn�����k-�^��I��[m�m)�ħ{J���f*J��(�L+zW��(�=x����Rf�UE���Q�'Q5 ���Q�6dw��
��>�x�;�A+�cإ���i��S~3�)�~/�#�������/��]���~���gi�`�z��+:5�)���Nb)~�F��cW� j��L��W�Z�0/s*F�j�0Pj�g�yP��y�A�j��`Е���,=�hu���nê��"�� �vh��>B�6{ġ�S�3�Ҷ��e#�:e�yVj���{�V�+�^���7A�o q��v	~B��7���=��Y��s�[���o5r��������xi߱ȴ"�v�����	��ݴ�`0�e�"'�p'<z��PB��2���^�O4���^��q�R�2���Mꮽz?Rׁx�[|�0Ѯ��~o��Z��Z�k_�� F���ϕ���VV
�WC�H�ޟ��Y��,w�X���\�����g����*O����$���)�߲B�^I�w����[����z�3����M�'�Xh/j��f����K8�}1��̛��
��-���H,�76Ў�$j�w�P{�H(�I&� >A��La�ڊ NrJWq"�`�#��/lG��!�������Cs���@�4�@M��|����=��y-�i�g"V�adi8�!4�he����r�����ʹ��Q��=�VkQ�4tƇ�ܳ�uɳ[�7��B�aý�x���Xv�~��[�@���g���ES����]�Mi{��+J' ��\C;�"?�Ctk*�=v�K��f5C~���Q���� |ٓ���5̹a7�Pn@v5�Xg���nAp���:�BGs�?�?�7�ɦ���9�sW��Z6�@:�ixI�ui�yr
Xc�����f87�҇��{x)�ѯ���|��k�z�O�Vv��9[�IG�t1DNU��6�M�GMљѢz(2�un��
�<��1�9�n�F��D%4�gww�{x[��I�����E uw,��`�P��\���R#>Fm,_Zu.rۿ�&�.�w�g~{T��H�&�� _t�m�~��"�%s���v,��]xv�b�5���Z���1�xw�����O����q! �G�|??7]/��\O�X���S`]K�g�kW�jW0�Ek�/��nu���H���T��$��g�B5����T�Ҹ3��Q�	�T���������<�Ӣ��y~g�3ⓖ��v>[*���z2��������NĚ�d��$:AMyy�>����R���R<yx�0��ё�Ex�(o�����X�v(w��G�n���RPϳ���Pc3�|�I\Y�:��g�/��7��nKy��%X��^������s�G6��yR�O�d�˂9t
_�9l�:hy������G{���<�*Dd��Wu��B��(�#�����1#/��KJ��G���*�j@p�Gq=�߶���#�#`��5�[����a����s���oU�Zֆ'W�5����
��@@%�=��iP��h���j���c���/4��X�j�����`�o7"��]�d#01�یZ_OU��� W�E�2�a���rc�^�v߮��#Ǒ���Ԩ]�GN��=����C��g���쳢�Sq¦yV�6@��"��tY�S�-�E�i�(ݛuy��y�u�Y�i�.ku�;��~zA��I-��m�]N5VMRq�6�5+;L�$�x�&�^�s߃Y�����'q\�w��������X�~���:b�����y�\�����?��O������I����r:���;����#C����^��MTDs�)�	�dJ3��-d8x��=��j�pn�gXwP�×�f6Ҳ-�lԖ���#��T@�D�d�T�gm"ϜJ�'��`�	�fq�`�nf�*���)ن�Z���� e*�)�{eIT`h}KWB7���F*��~���BN���I%E�3D���d�|����x]��ˇ��	H������Ť%q���<?E�7a�	��|k������)Ȗ>YjL8w4��l�o`��톻=|�ݩ�`4��|��m5���E��"����Ma^�߆��/4��;��e��t�Eq�ky|(c��F9[s�`����]5>_>��z�^o�|0!��V#�ټ�Z�`LF�\���EԨSwpz4WN����)�1_>���hl�s���ma�c�{�{d� *n���Y8��M1��"�d�31(����JȪ�*��.���OU���;Ԩ@Ȟ&0C�*1�qI�A�
	�X���F&���솲�_�4"G��Vͨ�=���@)�� _PE�.w���Z`��*��R<GI��eY^e��N��mr�|�^I>��V��:O]e������`_�����(6��~N�?��iT܉�0�
��� h�<��z�� QE&�=�!4�����f��ʎ�q�ȏ7�b��s���c<���K��-ʗ���)|{v*<������/?���u>������
}z���;����g�z��G���o\Ϗo��(�f�o�n_k�9�hiUT6=��u���
�M��Wa?�Cnop�Ml�:H]h�V9L�ʏ����?d�S��u��z����_/f�����)s��7��s�}�5LIDds���z󰗻�^r*�bi�y'sQ;����bя� ��:��z)C?�����ߒ���2�{��N�~$�r��nA��z%�����`JX|C�}��C��2�O���>&N���ۼ��|;ߟ>��
P������15t{��RE�&,��8"�l; �]����A��J��& ���=�Z��Z��i�Li�̅�_�?u?�z���ކ�o���Wf��n�m���TC�7�^�lS�Z�f�3Y�,��x�����$���uj���4�^/�k�j��ag�[�}��-�S���%r[bթ�hN�hk>�����f��;^A�������ϋGC�`pg$�	�H��?ʬ���P�����,?S��Md��{�Ҍ���2X��>���]�~�x޻E%t����>��e�fP����nJ�fpVo�0�Cu�܈P%O�!V:�i�#,��e�L�^�-��r�4���\�J���Ff���^.���5�a�%8���5�c)�U���$��_����Z�5�x1"��?�B�ݡ�҃���?���;����r� �j�-$kɎ\�ε,�D3��ܳ���nl�G~�؀3n�s(�k�z�5�����TA���~'�~_��P�����pS̛UG����������<�I`����ьr���-
���܅;PHI�g2����/�,S���{Z~$OO�,ro������^����=�q�N��p���b	k�k�8��7�v�K�*�AC~�4k��7k�!���y��>�����><�~�.��?d��z����ƶ�])�qP�3��M����Q�e0J�P ��΢��40��B�^��؟�[�}��
�l[�7j�'�b3g�!�[�L�<�Q����sg^����W-��Fz2�ޑ5���t�Y%S�p��Y�_7&��6����S7c���Zq%�G�|��1���H��ӏZ����^q��P�5�^�s������
!��x|(:�c����6�"J���W��g�q���g�(F�8��*熕k�
7�mܶw/�6�V�����T��!�������Hw,���
��(�=�[�*�\��4�F1Dfᑣ�eV��:?	*���, F(Y*����=���m6�=�q]��7�s�+{���F�����������G�����_����)�����Nq9?�����/ͧw��KٜW�6S�vX�Y4������>�j1�:Յ���E����6��=��� Z�����ꅺ��+h*��}��·�|��m�^ͯ�3a��Ԭ��1��6
�C�Xl���CQ��������l�}��+
�5=x��\e�'�J 2������[?/_����Y�Կ
�i<�c��S�X�.wd�4:)�0ރn�$�_��M�JáG���`	U��Xނ�^�O��S�Q��>Hj��X�K�ȣ�N]���y~92u��2L4wYv X����xO��ˇ��-�ZL��mpٓU����|�$��.���YM�er;�������]�|��#kh�b4V.��0���Մv�HYt$;�C�0�R"���HY�R�Q2��o���j�U�����ߩg��ٔ��P�^���{��cp����������K������ah�`�'�����Q��=Gy�;$�eg{���9��k�*��2CM���LK����(鬕;���U���m��aE�`.<�a%�����y�-oU����wP��+%�}i���9�7�w"���R'X��*�H�~�>�ax*â\��s�5��<rR�l�)֋���*����=%d�_�9W���(u��)ʟ\b��������w��<=�H��>������|щ<�-�g�\��t~���ǯ�Z�;ԙG(oҼNT��$��y���@��h�Xzu�&��d�.���`qԉwf��
�#ʮ����X�Y�fx��͡},gۉ�vM�b��ڭ��N��=���P�*�VEUlQU�vo�8��v��+�Rm#	l���������}W޾�L��b�;��>�I{G>V|*w��vh�`���R꽭/�=5T�B��z�~
�U�] �����龻v�����dyҒ+��C�Fs��:ۅE�wr�������E��'�;$,YS�g,�R��j���|�|������V5�7��C�*�|M�#Z*�yD��Հ�T�h��: #jpr�s�AHF�*�g�v<gO�ʛ��(�\��p%V.���#'�	��l��>k�q{�.��t<�9�܍C�>o����о({�ES�~���VC�5�Η�pxQ��f �^�7<Lf=Ǯ��p�� ����1����%ˈ�'��G�����zQ��R����ƽېf�9�_�7�S�l���`�AI�X�m�0KG뫆�6�BE։�@C��x�a���gȸ�V��HAʈzP�VR ��4F��K�� ��V�l���;��7�7=�wG@�4�A�p;�FS�
^oE�;{�a�p�2�)#�o����o��O���	w��Ǐ�����&-���r�����_�>�V�� �?+9�D�����Dn���P�ތ�J�<���}���B Q�1z�C�/�v���LD���D]FCZz82y��L�%k���Ѽ��� �k��A�u��9�F�l�+�2?r0[,g����Q�~�/9\�P4j���g����O�$���坻�����x�����>�s��r?����!f��A7��;=f��թ�r����7o���<�	�m��	�7E���j!���N�UE�^0�=�]�0ʎ�xWzp Ѷ�ݩf�+Bc�.mL1Ez�#̡յ�xnU�o�Tz�ln�^��z����.u��v��Ô�y*�w3�=��5u#�͇�0��a�����	r��X�EP�7��4�S9�U;�dݧ,�,��n�WȵwOE�T�\2Дzĝ� w��_B���+bvy�/מ�����i_�V3���9�lQ�\�/n4@bM�Ziٮ(���ӎ���l錸�ދT����C���~�B^�AK�H�؁�x��P������^���A�]O͢�9T�0We��h�H&�<�8�X޳ WCJ��u�_���P�@|_�eO<�G��X�Gp��j�]�G:�����`�y�������ȝ����.���9m��8�}nʹ����z�f*/��#e#�rT�	;��_ᡫ�D�M��~���B8��?��5���p�V~��)�ӻwEYܕ�9a�~�x�n>��篧ޯ��妴-��֯�Sd
�kiU.w�PK	�]�}�]>-�p��<DW�����db�&�ڒlK�hf���D7�O��?ف<ǟ{a�B�.�*,�1��|�<�gR<��X�Dw��jݦ�=��r�E�#<�{���@A���x�&:��C��x�k���*7���{E�iX��Q��r���G������o�#�h���hlT�-U��{� �(z�\eq�H���k>f��?��j��"���c2(N�/g�3�!0�נ[���Ƶ�&wE���p����r��������{ �s^�<g0�0�*;<�1Ve&R+7N�KG��{v��`�Y�֥�^e~����������U��e��W�a���$��^Z-�9b�A���Ú��geAiL�����4Sb6�we�3���_k�;���-�$����]�:�òq�ۯ��$���o=��R�7n<6�C�>v�-O��i�{ Os80����{��Ľ����@�j`��dW���[��As��_?��.���H�w�a�^&�,*Ӯw\ټJǭ君���)w��w�am4bi^jmuٺR�g B�)�"�"���T�����i�/:	e|�����gU=aE���}n�Ý�C�Y�tb�<��JW+m�]n�՛��c�������NW�@�fݪ�oķPw�m�9���YC��Ɯ���ǿY�\R�U���M��U�yz�R!�����ݟ-��_ZO?z��w��IO��fKN�=g״�rP�"���:�ⱆ�����Oͳ��F5�-�����&ر i"�K,���w(�Sq�)p@�;/�G>yY�������Z$uY�b��R�ŰZ��޳�n#X����+��:e�/��-���� ��+�,�c�w�5� ������;I�b�.Y���o�)�2V@ǿ>|F �~X���/ ������읟�����E�5M�	(-xS(dHKk2	X���ee)HP��i��])\���e�]O��VHF	�\P<g����Y]i���n���;֍=�t
Z�X�������#�	���W>E�G�W���2GE��/�\�2v��/㶔�>�c�OlMH�J�-Azu�l�1�F����k�^��pC��4T�J�[.��c[�c�ߣ�j�@���(�в<�j6��!W�&�����|�����W��zY�F�ʚ�F/(u��G%A}��%��ٲ��T��X�W�n3fl�A��V~]��|��\�@{�ym���|��:�v�U�r@�#��6�
v��16 ��<0������y��)G�o^_g|M8���{��@�T����^�N�^�Q2��j7ID4g���I�5�e�6�>I.���0%a�:�M�Ր���~��� �	Q�M<��!x� ���h��u��Ɖ0���i�(�U��p�J�|(J�]��ׁ�]�L]6�Dyٵ�����~��]����`z�S\�=1""�bK��QvEE��%��x�����ͯ�ӣ\���oV�6~U��y�����|�{���ry�3���'�R//`S���^�{vK����ۉ�{ܿo�Ym��|r��������jZ����P&XЁ�D��}C�Z���NoF$ӟ�<��Iw
��T��c��^�]�+s���p�Y�~����s|�#k�A0��I.E8^�<w0�t(J�(��0f��JA���;�k�KV����Px ��(��;ʮ���Kf�����|b��N�/j���roZa^�-�"5���^�OE�(X����dG:K'�(��pZ����֮��Ɯ&��|�B�y_ky�%�s�j��5����H�I�}(61\\���f��24l�7��ml�T0�_��-���kϏ�U<{O���e(�����]_B�����uL
����|�`�+���t�j���G2��	 �aQ� �0�M�#��%��������k�F3��/�H�zu���^��"��ЯG���G����J��(wϻQn�ѽ�u�������)�8����׮u�5��Th,|�M���1�t���`�Q�A��}���!��8���@�3��G���U#�u��
9U�ƣC)/u洚A� e�����@6;(sz�@�f���Q�2	�@RW�h༃�;�sU�����Λr8�Jl��/�?|G�&��J��n�����t�Gv�a�l,}9�3�Ǘ�vr���_�������7���w�vΉ4x���Q�$��տ"ǻ����r�!����|_~�w��w.~����ß��>|��H!�S����	�k�CPC�#7�e5A�7�k�xc�Nw�=��Y�l�ia}Iئvj������
EA{�@]<��K��Of��~���7 �&W�F�ҶP*6��9�����@��(�����;��ϏT�;@��%ɑ)t�Y�XD=����xG3�3�b/J=�1@ɸ��(�VTeƼ(<*�1� c[��B[�d\�
�t|Ey��cic��@�b,(*�8�T�V�<u��aC��������_�9���>m���B��(%�2(�����#�zܰ��Oh�{�k��cUVַhƗP�[��i�/��}����6�'%sx�QwH��[�u����)����Yk����W��ο�_-�bD�ƙ�%�g�_����&D�D�*��9�S��g�0�������K����_���E�0ʳ�~��fS��*W���u-�Bv�o��90!�y�V�}�����'�TY𖵁e@9	0HW#z��ޒ�#Q��ma���f^�T:Aw����Av��F9 'Hڲu@�JC�Q��L�x��]��'���e��7 ���\�SJj5��jm� Wp��,�Ψ���#��b�5
#��li� ���Q��'��7�]���d��e�$��r��xqGE���t��G����FU�Jy���LGd��pE|���~��?���ez�O����cw~�������3ǻ?F�������o,O��}�ˤ?	�������������K�:��ѿ6_>��r�����,��2��B�����(��#C�z�B����.d]�>_��Fl�΅�Y{o�;(�����`ĬV��֖�6��j�Y�͆ͧr��V_7��jt��w>z�t�|�m���P`�V����0T�r�e<�1���/x�j��ɱh���:'-J��<� ژef�|����>�G���ͥ��Aٟ��6Z��A��$�X7�_S�p�V���"S4���깣.tz����<&�����N�p`e�)��z[�|���{p6���<�����Buؙ2���T�����QO>�,h���&"��'2���	ePF5����gZ	Q 8�y�T�=���k	�	����h��B����~�`+�%i����L�ԑ�Ӵ���v����a������������o%|�=	o��^Fxxz�AF8�i�ծ'{�ޒ�S�6ɪrO��&�<qk8�X5�4w��֛����;�:��:��g�M��L
r+z*`o��ͤ����7I�v�ow����Jf�s���� #��a���SLf+�|!4�R�mQ{��U��){РZ}��*�C�s���a	�N��\k�=��(�E#?��rw�A��� 5�+Y�"�(-�bmR���̓M�{�<��k包�s����z���ȍ�����W� 	�X�n����7����������o��Q��Kx���3?.�w��zz��/������E����1�zJ���^}�����b��_^�_�L�~(i�uU�����)�\�0{2�sS�J��)i�o0�S��k������^�M�3f��2��,����]��Y��j�XRi��f�<�`���E�F�Y� f�H٨�q�� w���$��@�X�z���+n(�u_'%��%B�k���|*��*��H�v �����S`�:h-��� �b�6!p�،7D�`D'�i�]���N8�����N;�&'J�"㜨�I�h�6ʺ�TA�%�".4G�ܽ�����}U'O��(�$w���RKn�S̐c.�6Y`?tr� S�y�>�^�b&�x�	��\��\A\���U//(�M�?�� ����s���&�B���f����^W�c7��-a#�
�V�x�5����=H�'�2k�hDyІ�@�Q����[�3��B��p����hshƇ�_h��o�����'?2p>n�N�j��ޠ�#Z���j��dЎ�����o��d�\���2C�l�F��|]ƭ(��q�^aZ�*�s�>C�"�F1��tb4c5cdD
o��l����rN:��#Д����0p�*���)s���aΡ�9��K�b.z���i6�mvc�@p�ph0�|
�Z���&�e�@���J6��=�]��3���1���^��P�U�yv^<R�Z���h5��q �^�kz�'ְ~+��������Ç�����c<��7��.�Yb��e��\߭���^NOO�qH��,oW,��D��JT�U�B�8W��JD�є�hyg�vӺI\��B��J�6*xcguk�d��,��J�7҉꥛'�JK���o+ָ���Nݕ�e�m�l9x&��WE�vޠ�������M��P��=��_�sQ������l �@iڒ�J7�/. ���w)��t9��z�R'q"�@��:� �̆���\b���0��m*�QK��8�k�`"ܰ�$��? ��aEe_5E�C�჆�%���1�"F*C��{܊?C���B/F�Ս��q��s�xkY�D��╧����6H�A~��4[F�?�x� d��HE����?x��y{y�yA���h��Z�����~�=�E�Z�pg�D~D	>�8�}��lmO3�(����%�:G:f�Ww���YY9�G��Ywo��.�E2�K�����@pl�a���<e��Sj���؅��O��kn��κ�9���E��^�6����zѡ���F�2(��30

JvFU�Y�~��B���ܠ���d8�S����Ho����B������T��a�g��7��N���̢eFW�!�2�.��"Vn��R#�ڼ�;M�e��˼�^��3�k;���׌��Z횃��#�H
j�qR?�K��̈]��p��;�u�#N�Aκ*jȽ�_nijX���^�Œ粀�?����,�{w|�_��W��K����o�P&�nW��8�e~?~��0�{w�æ���7��&Xsò��Ր�W�#N�-�.�Ym��o<��+��m���t��z���!��O�X��W�UB������h���ϩ���\-��_b2/]|��í-C�n,����W��w����W�v���P��sD��&4v.4�������X�����^	9��bw��?��r+���A�T����k�"(�E�� �a���F
���cK7A�\ط��G�M�;�"���t���ר��qo���I-x�\L��@���潺���^Wh��@ܫ<u��Aq�,�X��t���Y��}Piy��x����.�]�y��6'����R �W���B�\^𸫡ZݠfH޶��7I�t���<l�zC!7Ӭy�����ׄr6�Bx��i��Iz0����#a�;3������*���*=i5�Cv���bƚg��0���;2�4(�f�u��s�Tai{С�U�(��@Xwz�96�	��p��C�l�.K8�f`k��/�_�����W��ْ�)�x'/����t���8 pV�夥���;**�ʜ�0n�FUi��}4åS U�6��
�ZD���ٕWVO��1j8z�^8�/h����ɼ��O�欶�:����c$�Jb=�����!zS�t�I�l{�y�?���� �G.�a;r�����$A<�n�C3��N�ةde��:�Hw��`�����ͿYd�����ey�_N��<}�5ٽjy�1_�O% ����b�}��_�����|�����vd�P���G��X��f��h8!�����n�m�	d�w�j�I�-#nl�B	.�sd^kf�C�D#!w�aRe�,�b�b�?�!9�a��1�6���S+��.=�nl�f�TO��C��+0I�
�<�FI�h�K}��+�B8�X��R,עG�j��J�p���V��{� ����?�.��yf��$�)�;B�#����
*ǫ�㡚���k��-q����͑-Z���"wAv�9�l�Rjq�j8 �ʜ�*^ h��fDqj�ddC�M�	��?���LP�n���Z��	x�����4���TҰ�z�D�fF��e"o��!��}�E��[w#�H&���uvZ�;���u���˕D��A�{9̛r�q|�y�;�W�7�y7q�[p��1�
�P�F}��0��憊ԥ�	���TƦ(��Pq w��5]N���Za�@����'�>�8��K	�*>�*������%kŬC��
a{&70k�q���p��,-]�m]��*���G��"Ζz0#2�yp����� *P���}"�YPB�n5��3����Q)�I;�r���)΋�����2��X�h��j�RW`[�F]Ng�=�d\��Ԩ�<:\�i4��H�Ȍ�[��`qs��	�R�m����
 ��e��F���e�,C����m|e!������fBS�`|d)�j�;k�8$u�$
��R��k��7D[&Ϟ?�LsFkHD}5:�&1�3k�K 8���g��g�����H���S3��,�拲��鼻�}�l�m����U���!��_�K�]���˸N_r�W���EeMO����d���伝γ.w�hO�pe5p�{_m+�{g��C]���6�79��Mx�ˬ��[�+��5�g�{)*1��P�@ќ�#3�.e�3��Z�֬��^T���{C���vv�\=�g�K*|�N�{-��Z�
�s�k����X^/
�28.x��lp���9��a�����bq�z�j��5�I��Z(ڽ�Uw��V9�:Ҕ��\���R58"m\k^��`�	���x�a��1Rټ�D���H ��頣���'��t��{x�QK���+S�k��=�1D���ܤo�4u�0�,{;�A�s(FJ�*�3Il�{�U�^����ж�K��c�O����F�˖��"K~�~m��:=�J����X`�i�d�� ���׳�X8Y-�X#.`B�関p���	4��K�?烬��A��3dނLF��-�P�O�u�s�;���-�"-7C񩣗o�xĔY_� �{n7/^���\���/��K��R��` d%�B�G3�c7��Xj EO���Z�b@�y1,&x�Eֳ��jT�Ҝ��2'�E��4ן�>�zյk[݇Nڢ���,��f�mx���|J+2Lm�G���cr��1jU���eF�y^x�+��"����l����]��~_�5�-%%'̘��J~�٢7�����ڵ�8}�ݘ���/��B��e�v�_,��/��t<��Ӕ����G�Я7�����ӍW�勁 ��b��Y���CUw�A�
]������f�5G�7���T!�usl�)s������7���H��,�����묗����Vt��x� >v�F��v���ϴ��ȊBNū�3s�$��!�0�arS!�[6-�o*�3-t|�aa���f�żj�!0co���	I9�~�Z�fz>l�������
�-{�o���]�E���@V�VU�/��5�l�R�.���8E�ࡺ��z�NAE�ymC������i�2Ӓ>�LG[��:��M,I��iTH4� C	��\�j��<�:c!�����n'��I��GcV���TI��](�5�T�F��-W�^T�P�R\�@�X��M0xN5��k�^)l�R�"�;�S�t� ����+J����e\��I+�ɈA�]�^ۚ/E�.\�2�|Y�I<<H��R����JP�"��t���/5�����9Ϲʯ�7M������;�=�a3HhU��0T�orHr��N�rrh�W�o�ߒ�z�����e��@��vy������Ϣ��e���AT�]Ǌ�մ)��ޒ�0e� O���҃��ү���j��L����X�f�Væ�5צ]eJ�� ����ݞ0B+`����l�25<?�F1U�N!�wa��c(�2n������*�o���&g�Ôٚcjs�Ϸꊬ�<d��p���Y�_��Af�0��N������(��?���!��5��z��@��}ݓ�_.�~x%��t���H�g�s�Y"�<#n�κj�\��j��Z}Zk�y���ÿ���s_�b����b�Hj����p:�a�[����b��l�+]�|7m�Iܣϝww n�$6���Þ1�.�_{\P]P炞j�,����}�
�j�-�= ���"~HT1cf&x�˩x�g�ۓ�,� ���_�lQ�FMT�(�������4Dsa�)�f�;f�R����U)ЋAsj����٪$�Z��Pj�ˌ9_5�5���U�5Pb�^����[�LYU���;�ژ�7ڔ�-3He((��S���|\��zb��z���j,rL��H�c�e�>�fr�{�.r��|I��5�5��r�H[�Y�����f��8��FSp����;����`G��QK�`
0m2g��!ܑ0FZ�;��OD$���`|���aZ=��dB�8�����Sj��������ӕ�2U��Y��ۜiV�R4�w�F;��hF��ٔ�a%˥v�\�eK �^KKP���)��A��r��(��#�qnTc
f�	���:q\w�}U(|�S�e^�G�
�_k��t~z���|v�]Ĕ[�*4��N��Q��$w���=4�&]5���'���9+(5ƀtƃ���(mV�/j��?Z�T����DC,Z«F�쾴[�r�h=�b���2��A�����^,ؼ<i��Ų{�|�?��b ������/RH������rxuW�O��p�6X���n0o&�J9h�`4��6ܢ�;�E�T����$7�i�z�b�s��C����d�~ּY�YoQ��;���� η ��>�ռ�zn���_��$�%�Nj�lY�`���(�q����ղ���ٰ6�8]�����_ɫ�D�k<���<�u=ɮ̻#�;�6�A]����q<)S�7�q��`�W{>�<�^_]�b���F��9.�[�S���kٻW)󟗵4���j�\�,�5���ê����Sÿxл�!Q����Q��a#v#W<��<��,ݲ�0�ؙ�z�ȓ"����F8*VܰA�f,K������ �^k�PG��j�V���Z��k�~�)��G�p��h���H/d�AO��ֻ@��Þ�º&����j�!_8	j(�t(+�)_��>�$���`�,{K��^�>-����y�����)�l�@�*n<t��k�p���w��\W4�{�;jgyoW��N��bH|��f�>(�J��#E(t'a-�{��x���c�̇2�����2�߳�C�=��_�8�\.EV\�ф(�x��[h#խ�>�A�s����^gk P��#Qcx,�O�14J��I�����:C�FK}�hA2'�S�T��,JlFͨ|�]���T�����/��Y������6*:fz��y���>�(�N����r�2;�7�C���d��Ǹ��dr��d:�dBn� ��-H?4>�
ָ�k�]�݄�{в�T,d�5�ja�P����^�:k�-�TE{��u5x{V�f�J����[E�pc@����/yX���zo!KO������wEi(���c�2(����/:_���e�����<�X>��7��}���?��˗r����H��x�[k/rL-��FmF�]x+3CX\��BL6�5��C0�}�J�j�n�[�U�Ì��E��\��z��/j�2�s�2!�˓�	6���  ��(�	�rMG��쵁�iJu� 2�({������LN�'|�!�J!�0k��܋��M]�zO���-B��^,���H*Ą���hB1�wW���~�t��=n'Dhj��H��ܯ�e�~P�c��!�ދ�P /�׈�l�j����TJ(�J�{Y���ԕ��h�l0�H	���F��8YjE�EANq^ߌ�'����?���d#Ϝ��	����u���[�n��O���uͲ���酘�x�^��T��h��S��H_15�ߧ��O_�r~'+�9�1��YRԸ�M�/�{+i�[���S�mܺ�Q���a��"Ug�v��ji����1K�{��C��T�u��'�*I;?�"�CB6��+t�1�^�@�0����Π�"�:�W*T\��%�2~Wˊ���S�6E�
�F3<E��e���;a2� �f����b�9M��ray*�x�{F��#�t�-�+��_2�u��W�fZ�8�?�2W��� �]U��Ԉ	��������A=�Z��r������O��lR���Dj�X��^6�q��u%�߫�s+�ţ��f����G#���_Ex�7�y�B�zF��F���l�f��`��V���
S�e|1��ꗴ�T�M^C.�@�`M��t�K:˵x�;z�څ	`%ҷ��l�_W�k`��0�+�D��Us5��ZUw���ɐ�bv��5̮�E�tRj3_I%\9�E�!+�y�Y�A�Ϻpԇ/:�Oҁd�m�'���%m0Z���9;Qs�S9�u���	�cC����|-�P���,ic�-#|�;`Q�����͍d�Q�5���D�N�g| �}���T�\�����%�^�E�o����S�A�US�̎a-�IM�hx���=�f
 9�.RG��|���LX��yR��e��	�Zd��9�e����<��K��)��,�B���d�Ժjz �fT����x��OGvΆ|s=Ίh
m>��I*7��܊���^$�B1��ӏ�B/��I��;&�~��>X�ԓ������si��s/��m�#�{UIg���4�<�5��q�5:��W��D7R�F�S��⍲D��B44+��:_�5������ƃ;�v�xR�ol|�ը��!�ֵ�K�(���U_��)�Ք���$�������1���[�q��:f��&^�o��e\���ڴ,6��Yǔ�K86d�7h^���YrUug��EZYWP+?c�&��'�jq���6�D-:��m���s��DVj'�mj�����m"�-M�D5�j��;@�7P}�O��n�v�7��(Fs�s�4q8�p�Ѯ��9��L��;pYhZy���4/^>�T�2��M�ZԣKy�۵Eu�1R�g֍5�Bnat��l�'"r�F����K��^�ΤOP�%=D���׉��m�l��mfX�sX6�Z��zs��9\�/��Bw4�S�s��Ra�Z�3���2(P�Q��շbp��]�EC�;4	v��Rk�1�E=v������H�k�>E=�$-�Y�Y�=t�Udu�ʗ:b;�ڣ��x�Rt9�Z����cɏ�� �O�殏�-{�@yG�R� �[�rH��2%b�kxD������qB|��U��%w{_�
�4:Ae�-:j�����U����0D�QC�.�U�j6Fd�ޡ�/�+%ș�[���H(Q?�T���1ƫM�c\�%=���jy�{� o�-G���ʉ��D������x���Te*t���*V���б��l��u�>��1����K�������+]ĕK���,5luJ]��T�k��D}3��1�!-4X�{�Zme�N����Q����~�y�P�����\qЛ:���a{S[�f�����)3x�9I�b�Cgr�#�pP��8	qG �A�%��dT3I1p	�v�Qe�=���bI�GQO&���^ƽ2�h��);Z�^��� �$����e�ު��o�+sg���i9fiHy�4�'�����Ud�1r�-�;��>�	�g��9�]k�]�)6O?�S f{�+�>�_8�4� B�)*�o͚'�.B��a�'�ZiT����kFY�P"�l^�������Z�w>�{h.�]_�sQR��v��M��`����s�G�~�U>6$�2GG-��$H*�n�O��j���rϹy��[d�om�U�W��e*[�4���#䦠0�Z�_�˜����h��O4�P�^���y���e�x���T�Us���g�u:X����n��u�y"������lF���ڢ3��{&U��KD�P���F�0��j�v��,�*�I������bYҵD�\�8��W� .����x�.2�B��K�'-=Pm~�+a�c���N�8nkIjtI�8��=��"iN��yP�i�����|4�1�M�w�W^���Tʀj\+��2��!<E�W��,�>(ۜ5�5��|��ӓuTZ�L�uVC� ��'�2!Xʴ�u}9��۷��o�][��H���t�xj�J�5�orP�����~H��y����������J[�	t���9�����T螇�]֠!��Lup�"��b���`����9K#4[�@*��`Z��Z�c��1���w�t�if�&.���ھ��4���	>[��֐OX�D9ٞh^�vÈx,.����-��{�m/��K(t ������ÑN!l'����$�K�e�����_oy�f����E���u�,�r�,�|fDdUJ&��&�8�Z~�� [nz� Թ�3�c_����{�ˇ���]�-o.��4!�~P�=�U�h�og�XH3%��Q��HqF����7c��{T:���һ7�a��а:Wm.�3�T<�� �������/J�м(��uR�
Q�{4����= �g��%3�@PT\�W��8�d��F�qԖ�=p��2��j=����d��+����[��{��ކYuL�+��
G-�A;߻�.ʚ�S�P�>� %H��A�������1��ԹGid@��9��-E�C��(��o��<�/y��(���Y+]X6������TCY��q�A2V��bڿ��]�j'5
��fP�Z{��[����Z��+����j���a��.ZX�5���an���z9�8�}�5���|p�b_��A}:�Gft�5�:Q['�)��c�Ot�MQ�x(t���5��3k�n�B�^�����4��7Mf��
dd̖re��3�U��;uF���S�7 u�4���wv jߝ=��u[7Ր��Em���X��j�:���L��i7��N�3xogL�*����, Ve�̄5U+�X>1��Ͳ	ղ�&p�y�=��ج�ؽ)�d�bo¯�-;#�sM����oW�z{!:)!wO����J�S
]ﱻyq#�3���o��S���N�u�j�QsE�����Dm4��|[���TVS�k]��pV0�\X���/ ��2�ҟ�����O�G.�����ox�����ɭ��Ɖy�®�\���B�h��y��Us��B�����љҎN"�=���l2�+�vQ�1޼��@���I�hHvd��a�SK��������nH�%;����Y�:�Y�ͨm��V�����O��u��$��/:T�\'/� pѽ��@Kւ�!^�!���ѭ��� �8_����MQiL-�I5��'�,'�����F#=&rVG���޲{��>zy[�3�O�p_{o����)�*�BS��2Ou��=�Z$�ys��>sтqT�cP�~9�.�������|6�G���{y����vd&�Z�tU�;�ᄓy�����F���(5���������{�7U9^���9>�h;R�J�D�����S�!v c����GH����W[��h���-f2�uh��K��/lݔǮ�a�����t��M��%*k�����X$:�,	Z~�����������4%��A��?qD�兼!�ߴ�+���ArM�6ewd�5o� @�e�?�k����u��n�u�&��1ED�mg����ք�ǎO��)���\��V�􎓆m��Z4����»�}�>[��� H��Fp��.Ys�:��	AX��H���9'5�ZAdN��p;���\}��u2��4�:�`�*`-nV�N�kf{�ME�k��ec���.�W-d�ls��>��\H�JO*4��Ž�' �,���;t�4(���,2b$E��dB�Ě��|ءMk��!�u-��Z�?|M4�����s�o�"*D� /C=깷X;���-KW�z����ޅ��bWe�J���3�m00	[U�.��+y���~u������b(ܽ"�BXic�F��O����@��1�8t/�M�on���C��\����h����ޜں�{��ޔ��1���UDIt���ǫ(��b�u���):�_/W9O�XT�|���������P@a���[��c����ɯS�ٍ��1k`����椦�����"�	���|�n�<p:��dS�jWx�7|q|t��'�<�փ�+MK��������p�%Ǫ�=�Ө�?&���tG.�9�b��:�t�rOM��T�����b�FPY��B��e�P�;�<����5��rR��$+uj)$�7�M���ɸ�T�5?%n��{����Yn��d�mYN���o�u-��,�q���@�k��I��j���b���d��5��i�
2 �Cq��`�,e�f#Fl��� Osy�Z�n"�.�թ������7�W��7를��`t���6���NĐ��Z�ǋ��S�P!^T@w�첵�$��)�K��t�vmv���s�C�u�:�ʎu�L�X��yV�e*m4�*����U��!�O�?�yN�7�ej�Lq��&��#����x��qhy�m(>Kjv��ﯼY�7k�ז�:N��9�u�Ϫ0�s�8��(%?�¨Mfg:5&�5�����؃g�Δ	�8h�U�+K����hS
��cq͐�0ߤ*nU�ye�BW���D�f.t웧�&�z�=B�wl�	��@������.܌�.�Շq��ȸQ��\�yY�3x��c�s��B�tr���i*��|�ӗ_J.?������#�]#{+^�ݣ*Tx��v5t�����<�͑�_|�Zt�sp�$�x�7o�U+���Q�s�fD��إ�q�'=�g�q�̽dN��E'����Lu�J��5��l��|Tm~�^$�q���t�ь��YBL��1A����o��.�r}z����s���ւzk��<n���1�������&T�Z[բ�������gC
�pb�u�s���iH��s�m�N�Я�Թ;���䣇O[�yօ���BK��?zv�hc��)[��>9�cQ�.U�^�'�f�u��:@P"o~�>3DO�T���� HaR��*>���A���Q��	���z��d�P�ZZ��^��H�bV O��k��S֒W�L��>6����`
ٵU�� �X�	.�k���T����D��@Y�H��s�S�gۯYs�@�/��uT��}�o�2[<��h��^�	��c+���E�!���-g��x���Bl{D^<����3H=O�)�A��).v&-c%���S���Y�8_AJ�P��!�>�.Zb
Q):��WOO��){K�V-QL.���SJݘl�����g.��q�ѧ�i��-#K���[:��L=E�e���v'P�Kf�K/Yˠ��9o�����F[��lNZƷNgF㰗�W��1D0�2�^)��O���"��x$�/OOdSŜX��л�]s��alo�^���؅~MuQ��}�f�\����a�x�4S�����Y�7j`[�����1���`kC/'��7'��B5���P��?��C����d\V��Z6-�#T%wZ���:��Е`6�ࣩ�c�ܢʧ	:(��$�|-F%B=g9��i��~�xSɄdp�!6!Ѽ�ҾT��/�`��!�=㩛�I^�Zۘޜ�n��p�M�&�:�F�J�dl �`�V�<yp�g��6��ã��}������n*�ȸ����V0e���	9��+����}�e_��+zI�*�Es��*�Ȗ�'6���NP��8/sA�q�.Ve���'礬M�se�^��jW/�}�.�a��:˪�W_T�F���.Q���5`sXC~m�5�csB�.G�i�K��tm-?W۰�jȬ�w���0`�T�sE) b ~�ݛ�L��6��!��fy��$)BXؕ�ꛒ�j��J5Y�k�)�X݆@�OlB�a}�ƨ��F�Q݆�v��s�Bq��wķ�r/�e�O|_NE��"�V��e4�����k���@���l\�B����YEpk>1�=g/uꗈ�닥�1�C�76��e~�QŮH��F��y����vņy-��r�F,(��XΤLV$�������|jb��"�o-���ZU�'��YB9����;�o�;��9?��L�H4��e�����\�����d�Ie=���yk��2jȇ����\/�H����q������j��>W�Q��J�}��j�;cb�r3���9�UYVI5:C��U��6�^��;��Jι!��Sg�(�Zw����ӥ?a��V���^�V�H�"�a�`����R�&\�ʈ�sq_�g�Q(��	�TF(t�8��Ud�z�]TZ�ƌd��x��F��M�ӻ��EK�Ue��=�mq���t�=����{��S��C�i����5Ёoܺk�h�Xd��8���">���٨�"c�˥�+j�͆A3�(�e�,eU�d5|��mDb�D6n��	�Us��J�C�0{NT	�1c`���A��=dޕ.�X�"��3u��Ϳ��0up+���i��l@6����k2wF*
,?J"���b���F{4쌶��ߕ�q�#��7
�f7{@�v���zdqnJ�[��������r�T_˭�OoU�**����`�&�TЈET���=m��5f�J���Ns�'�aqlJ�[��f4��k�zn}4��ހ7{��ą�&B�c���W%����hBY��A����^�t�̧"S�.�r(�X�A,DB�l�>ur�NV�J��RP��|.�j��"����͞�3�g��z!qr����k�����;��? �}��]��:�w�K����}���G����B�n4��W�i��ϛG5����S`&V��й��c��&��YGH��a3�ӎM�d3��V`�<�k+(�w���b6jZ�_HC��;zd�`�F������:�9��kx��e�\߈R�9�' �4x�B�5��ቻ��=Z�=9����s�����t���s�P}�ze�^�NG���~{�\���=�ݤy���_c�p$C��m������<��,r9'|R6$ ����n��d���m��R]-̥u�qc/������|�ڂ�\�y��m̭���Bwo��G���6v/�7���Q���T�,����H��#�U����(�~@/o�%�JAp��,����J��}��C����<�~GR�f/_�O���j%Gv����L�?��-���V���=�����/|���&�������N?����6˯�6���Ssw6�*'+u3*MOC��<�>T�J�����u7�>ro�w��Y?����.g4���)���#Zs�����._���\�/ܘ_�aKm~~{M����u(�y^h� ��B��f�@�����'t�f@!R� ���q��}�B�`Z�k J���O^2���P������J���s��Moϫ�j���jx��KV���[��,f!��}_�D<��/�/g�>q]��C��i획�0l��#Z��E6",���6�QJ쵞,�JE�2�)fӬ�ͤg<��(�l�9j�=��?>���s^ܟőϣ囌|$/��P����IjzU�a�5�7�_'����Q����0|��7��	�ȿ�������]����E���K�D�د��@♋��N �q�snJeET.F���o�Z��DJ�hD�TV��w	�AS�h�{�aC|��7�\O�m!JEs�u����e�q�yގe#q�Ǻ���戊|U�R�����.֒4g C�c�qI����1�^^Gg�W{��wk���ft�<S��~b�ޚ�'
j/I��9�����^Z��k��Y���sG���܌�d�
��IN������+�w`�u]�� ���y2�l���W3��Iޘ�U��d }�=�����V`h�E�Qۛ�J�`�t���C9_��LG�f�"OW���漸�S�,����k������ X�q
�d����E��	�LO��q5,��)����s� =�����W��I�q�ˌ~�De^�q�(l��d����V���\��mc��f��jP�h�D������T�������m�}Иs��9�}����q�Ĥ	�*��"Tj�����_��T(�*�TI�6UUTR����
A!iS�$�$`'q�q|�N��{�}��{�9Y��c̵�>�~�{Ϸ_�1�c��c�>/�1t�B�q�u�=�]x�Ơ_"X�Ew�f�g-#(Icǚ(�j�B�D��c�'��Tv���O�b�9쵵!GAc�b"���u4�����%#��Q\-�B�y����4L.ׅO7��^�
�B;��w�.��+c�M��������1�tḖ��(4����h���'-wt3���F$7��I�#�-�HL�fF�N?5]ł���7[j�T�0��#� � r��q��e���ۢQ�Y3�&�33������y1K1;����Ɣ��\6#� U�[C��T��HQ�@����\w;n��趚Y�r�ɯ���ū1�{g�I��6�u���J?8�]x�}�\ô�]�馝W��YQ��>�f��YX�<�YE�dAZ�k�:��d|�+%�{O�U>������J��,~���ٽ4�a|��>.&ĵ<*�����\��X�2�-��e��51��v�����+�na'1�?]P�H������ح ��N!���Q�s�`�I{�}�X�[�Z��t��3�b��d>�q�>_[��T�[�F��?��5�����/ҭ��ug\Q׮���
NâpW���h�Z��Y6�@I�퓺�80�lq|��\p�i�
�#J�դ�g�h\+��Y���!����mĚ�N���IK s��u��}�Ќ�%�
��ڔP?HEYj-Z�Brs��%�V�n2s��e�_����Q��h ���V�]�6�%e7���� CFٓF���iY�I*�OU�	��
j_�����"`Ò�{*1�=������]�9d|�nbT���h�p�#�i�&�x�c�X����?���0���ŝ_�ĹK����<G*8un�Q��s�}�Y�/ִF�n�axO��vX�;�փ��tӻ�7J���CȠ)Ow��ΩT�5؄08�Yc�۰:��{�A�����fD_�i��2v��U��0�6ޙE~�n�Z'Ԉ�o��7�����`��( #�=��q1Â�|��<�4�[l
{Ũ+5#�}x�X����qL���}qa4Ɓ_\֕�ĭ~rGJ��&��V'.�49���r3 ��v;y�,Ϝ�Z��޵�]ځ̜a69윀7�˝F|��4B_`"n�V�9#�tC�@�[~o���z �����i�=`^G|������\QK�P�CI�*����Q�f��]8�8����j]���^+����!u������%����V�(��r�0�E�0�i�b*��[K���63j��Z�����f�q�dj���#�)ƓX�3���������:7���R6p��G�(�NC��wT��R�u'�Q]L�3Ўj�ڔ��]�^&�ɻ���{�~��ǫ�ۈ���Ns4׉��lD��q��_"��T�j�\���#�������ALk�����Ê
,��̚�!#�2ݎ�W�\ڵhz*`�U�%d���?# ��E�kc0�⸎��ÞfC1�-�H�ܥĈ��.񹷑0��-��dk����]�/��8L�v�<f�=^�\�u}`+�hȃ V����0Q��%
�f�������X^�����܉�ee�|N���z�\d��܂i������V*e��a��|���.w�P4c��ֽ��Uq���l�g�c_m��7���:�=+7[U[\.N+���`����e��V3���͵��AƁf� �@��=��f�p)�2���iܮx���"��Ê�qL=!�X+�3�ft'L�yh*̊�Ϻܝ�G�;	}�cZ�Nk��D� `$@�q��H����q������S���h/}g�W�ݥY$�	�ȿ��Ђic�J3�5 =-�c�Y,W��3L��-������	�f	1+���
XpM���G�o2$�j�|���K%/�k�3(�|�Z�emC{�t46��2���@��׋��_���Y�pQ�ެp���"h�V#`��Ͻ�5bs������(��	�T��F�.�R��@�2<-��<H����=��ʝ y�)&_�ۆ��ݢ�v�ia�YG���o�ڣz!�+wf�e�\�ئ�][ϔ��Ev�4����{�J]P����v���FVO� ~u?$��Rv�ýy��Za��+A��"� bgA�Ҁ�"��royN�ֶE�qYd��#����GAP�JŘ�B�`!2�K���[LZ�a
>����lx�k��ժ��a�~�լ�E=��f����ƥ��L����x�gQT@����n���'� B�!qP�����4�b��� ���S;H�	��him]#.0#�Z&��юu]���ȭQ-�<X����s�>�g�5�� p��fm��0�e:mIr�	�|,���ik��f8h����s	ymqP� V�R�	eM;J��Yk}D�j�a�Ә5�3�86R��3f�=Sk:�섶혠�n"�͓.�D� �����4�B����U�g9]�ok�`/a�f�=6*^i@���Z�b$�"4%H.���NӏM��g��+��P_�9��^(��&J�T�KP%2����s�Կ�����t˛YS}L�Ե;�ۈ2���e����pÐ�t�$uD��NQ���`uŀ�[w=7482���ژ!LfZO@�"�~$Iw�}�Ih����#N�-ޠ�4`���@��bܪ���Uo�f��T-��Y �;���������y�Ǜq1����kh�Y�V
@���,�&[�J�5�Xs�6�y�LȜ�%+{ttjD��>�l�v��G
G�񩠐��|>QUP�܈�(��X�,'q�; ,(]�K	)�̤� �8�.i��pz*|����!�k����œ�j.Y����N�>,����j��1q��x6A�n�r��i�wgb�a�� ��oT�U�����z$���l��8nIﵮω�n�<��}8ϊY���Mg�����q�Mx"2�wD�Ϳ;�i���,^�.pW��NR;�$���Z����I|Cާ���#R%t�@sf��%?H�<�E$������ :u�h��n)Hޯ�н�_w�,��"ť�\��{7��4 �u3����i��d��:�g���ɭ͹Y�/n���� pz���'�o�^�ƚ�BaU�sg?�����n�h���'�6�ӳ�Q���Y�+|�X�`����_Z4Ff�m�*��7�j�#r��q ����w�`k���Q!H�,v�I�aM��f�XZ!k�c~t�Wj��e��j��
��]��ʧ��`��ڄK�O?q$��*�<zw�&V�RE��],͚eh�aA�	=��O�	�#K�k���������z-F�Z�#���|k	O ϠWy��`���k0���7��o��3���y�m�c�f"�r�q斩];�7{��UQډ30RP��������x���Y�Av��2���]Z�oRZ�@�G��rof��ks\>c�K�8=ZǏ��LU�e�µ8W�v�/[.��{��`)�"����t���ުR�����c]���������y� �u�]�:<:�4z>��R`^��p:����b��ʖ�A7��I{kI7Q!D	6^�J6��``�:� ��Wj���y�v͎��>�P*�	mC�j#�<M+_ԿT�!���\sʛ<�S�fĝ�w��%�@!=�<��.T��[Hz��Ͳn{Y;Ig�G��4�M�ϒ�dk�01�R�+� 6!���tuiz��ݏzBր��t���^�'[��1��w��`9�qVeQ�Yc
�����,���,ǿϨ-n��O��2w��dؾ�̹�0u�G��%�$��|�k�
��q�����t�HFk�R"Wz�	�*k�)�bz�����-&]�*!q�m�g5+V7*�J�iׇn�c�L�k}�z�u�F�`aL�k0�.�u�	��x6�^XZ������onT�������T~���E+\��t��b��Z.�ia�Ga�w��o��a{@S�w�]�-Js� �yŗ�����9�������{C�z����.��혩K�Izbh���b}�hq�Vw��P��5c��G��a�����hI�K��K�i��yP;m��LlYT.� @�F��kD�"�P�F�f���nv0���Q¯� !�q`��I�>�a�ȑ�it���������u���&`��_ ���b����|$H#q�o�8� �`U����|����W,]j����q�	�3S:J&:�"��֧!^�!x�y�)\.�Lg��M��߁ ?D %���D51>јM�q��G�F�)����Z����L1O6��0�p�\�+��axI���'��(R	����r����{�wt<�Zh1�	���e���e���h��<�3y�����.���>-��ӻ0b{��0�!�#s{DFg�>0fʖ	��{\��yuL�(,��Θ�2h�S��Z��+�s� ����!ɞ��Ip"�7q��"f\�7P_�iq3���Gm�;K�׳�׻�9rt{o�]v#�����·�Y֒ �-|�/�~���g�^-��[3�O%���F�"�cA '�<�_W�Bꑠ�w8���S#d��vtް»b����� ɿKᙖ�>�];��&���pԤ����E`,��TJu�är�S~��
�6��ถ�ň}au�Ƒ:���hv]|lf<�VR����sN�0��u�Ř���+y�9���L�a����I�R���>"�X�G@f��ū�T7~+A���̠��~��h�04�q6kAIa�֜� ������+ENnù�
���v:gÑ��k��9�l�*.w���H��j;�uS*��^��=����J��	��Q��̆�Q�Y��xp������1u)w*f�es!��Z ���ݵ�)�W�� ���4ֿJms�"����-�k&"�C�R��� ���x�C��z�A`i-}��	�U3�u�y�J8.�u�7��7�(|'q�2u��EF� \�,��Ѫm~Y;�tn����e ��I�ﬡ��j��t��>�ܵ�R1	Z�%@��^�w����J�����f���^�a��nx�E��^��k@�*8�=M�'���}^] �Qg�g+f+�������'wV��TLY����,+�
�P��ӣ.hlV��O��'��"��F��%�yF�D�畡��Q��`\S)D0Fri)�I�=j#�Ј���x�Z���!,�v�;~���	3����Z�&zGzF��:ޖw��i�������R�ŊDHY^�0����
"��1��br?_��!,����Ee��Z�}�x�J�Ɠߒ��.�K�/6{�����A�^JK�+����su;T�����c$��w1����X��� }X�np���� ���~q��D@_}���\lN;� ���I�E��(��{�;Msbߟ�&��-F�9�j!��&��Պ%�>f 9qWᔉ�X�s���M�#bB@G�a1J�]�(����>�� ���8hό8�n��Ҕ��x�6�$;�\��
=�CҴ�b��n����1�gߏ'�ة�w�Ҝ%�� ��2��@Ү�2��i�+ h*��xD�M�NG	��gk޵���PW�q.(��x�.�U;�us�ٳ�k)�E���\4��!����4o���YBd�����2����Z�@��Ҭ�s�֖�m�s��z03
f��в<��6&�Ŵ�6���-j�Z|�u��S(6�1anҶ�I�Ō�C���������t"�됬1/u3��bE�P������ыC��L
�EϚ�k��Na��w�3�� f%!tz��5a��qJiJ�>�&?�Z����`J� ���B��q�K!�u��'�>N�,2��[o�4���L�G�9���m�g���(�16>C��0�?s�0W��ҋ��G�?*KI�uIT&S	e-�,O�7��%
��\w��-�J�`V�G7?�!
��ӄ�C��E�!�=�> �n&r��b4�}"�k����n��V@�}�XP5N���vI�*yOK����������H�ͼۓV�b��^�3x���Ü*x�H���|!O�=�M��s�Ҟ���A��k�^T���,%���d#��W�t���~wRYF���Ýu�d뇔��b>fF?��լ>5���̋E�a}�^�Ҏ���������ʨ��ʄ3>��@�8�\K�����z�|?h�X��N��H?GaJ(l48�:6d^=��s=��	��5h$����e&^sC*�
n�Q"�7K�#W���ERM#���*�g���_����;.����U�pZ�D�X���ղ��,�P�?hZ��|B���@|����	��b�Η�d�	�#���<3w*�+��DM���\Da��m���f��V@��'H�(����3�AtqN��5�~50 �13���c\��Z3h���@q3z�T	�vճD���9,7;�`�V^�1Jܴ���!���hKb����=`N����º:|-"7���[��I'Ɂ֍WA̻�C�;Tfd�M
(ml�h�w�Vl�#����FC{)�o����y�V�o<^K׎b��z,��hu抙��|�6 �[w�h���Pn�e�����Ѿz������b���颦|���O]�*Iv���JѓD�:N����srC>�>_Y�2m�� �8�y�ZA��i�u2�ܕ����$��u��w���&s�Oi��m��6���&�n�_��:�������i�KVә�T�T���~�Q����Y[T֌�ř^C!�0
K�Z��z�R�dVU�X��r'V#$�1���LXXP�X���p.iA�ϲ�;&tu����˖�5h�*IGl��b�{HH���H�ڱ�y����9�:����i;��.U¸j?�j T�Y�b� ƌ��l��7M�C�"'��	Q��ɢh>�dD�9K�f��6	��KB��B�p���+�2s�<p��O�H��!Ee	��^n�KBɈ�ù[�j$d��(R �Z4�j/@�ԗ��V�fl"f>Y�Xh��n�w� !��̓���9�l�g!rZ����tuA�~;]�k��輐k3�ti�5*�ŉ^�]�g�C���tMɓ�SP�M�ݘ����h�L�JD�7AG��t�W!iw�U�%��fL*��H�݆j����a��'F�y��g���r9�k��D]w�YQ�+��gۣ%�1gMٙ��M�rww���z��U8i-�؊a�:e�L����G�kDN� �\�B��  �V�%���t�,�^�"P��O�����:U��r1�s:SU�����[g��')v�4eB��,������k��/�����Q��2�둾�{蹊W��4 �R�"�~X�v�=df�6Բ#��X��j�f8�h��AV�<<Vƅp�����m��A� N�C6u��ꎙ#	����sc�Y�:k�ZjR�gQ���-�h�[�m.���QD�$ؤ�YM�z�d�NXL��WH����_�K�3�̀��ʚ��ֻ�t�f��C�M�mhX�Q�&�s�S�k5�"��\�0�hzE͘RX��gr�*�8J��������C�:���-��!���^'�MՀ_����<��@D�?6/�S�-�6��u�{B����#[m��ќ*�[`�3�Q�^�GlS(�!����,̼r+C�?�_��n3�f����}��8:�AV��<֌��o�9�[+��|�v���Q�+�k��ǯ�d��m&�{�E7�-�;,Iqm�j��M\C�JE�Q08�#��bKp�`(���$�ǵ�ٓ2�������\�Pa��Rm^"����,����#j͢��j�2Ƨ�e��?��6�*,p��q�* 0��~�̼j�k($:�0������:@�-�}	f~���"���P�����g�h���Z�;��"�u�E܌�����ޭ
'Lc�VJ�M��E�L�h��p1���&�`��My�h������-89e���	a�E����_T���T4���1�N)��4����&�����'�m5���+��Ȉ+�8&(C*	�J7[�{���|���K��I(�oG����!���D�v���}SF�+�8BjR����JT̏H�'\L ����[@*6���Q���}M���=��}�N(��T��QNY�`�I^�2a�D�)$��k��]�m- ͥB``�ؙ�s�"�����'?٫H�u��7�{Z6����/q\g�����>�z���n�:�d���U
�2`������l�5�k���g��f
�� �s�5��k���8���/�"%i�<�=2�{����q���p2_�Tw;�/\̭�Ћ���|�#�ό����f��n�`�)�������q��9�a/L�S3c���R���G�S�>,ِ��>?�z�_��[�kz���S��5S;�F$}[$"�%�W�;W	�ě�Q��<��ݢ�	U(}ߛ%H�W���R�J����3&���˝��5yA"z��$^0a��BUԷ<+aBp��ު�#*�vc�
�t�QzFE�,z/�ܣdkhU�|i��S�6}��&��s7��x��c���=��@LH��>�1�FT[It�q�$/	�`��;Lm����Qp~0�<Y���K��B��f�����Ho��7O���tѨ��o���	�1��QJ>t�f�N��:aF��݂3Y�ٱUj&�IX4��L��W�G�:�Uql���R��jz���㾪�D�,i]Y�F��2ФjE)�$�:r��t�u|yǥ�k5Z���\�0���m��\� �w�2"�q_�����9<$n�9�1��И���˵Ҝ2���эg�B�!���
8�&��|U�&{�����̍V�)��R"��4w�=�>��F�K:�^���ٞ�q�uf��-qK�:!e2�q/�u�9�5J���-�ס�"�C{i�
Xo(�����	��
���k����Vz�ݼ!���T����0X��h�J�|���*n�|�\Wdn�=,�U��"��ϳ��U���>�Z)>�%d�i)y�������Z��?b^FܻJ2����ɢK[�&�H�Y^$4�&�K'�W�?ؐ�z�X���\k9=]A!�\c�xZ}]�@�|D4���&o��g�ʈdU)Z
ZkE�h��إ�Xҙ���o��ʠ�Ήq�wS7�i/�R�P�N��0�|��%L.#�����MP�/5�l� 2���&b�Q׈1����@��5"*V3���C���aL�w��7�ڜ�g���]�Hf�����Q����jy��̐�- U��vg�:��P{Ȳ�eI����C%��dyٶ��^D*	� �_D�*��@P�$m��������]C�K"�9�b�u��H\td���+�}4�$б"�(�?�4�:HNO�>WÇ���I�]d���T-�c�,�������L�����T���ր��V��d����/��J��v�@X��?ܪ[w�D�Qud��$�O���"@g�Ʈ4��XL�@|K�)~?�BKf��Ǽ:,��\��C�q��@e�´2_���D&�5�I���Y��Ц������$��|*�|���*kb��/�|��8�N�"~�N�sJ�Hx��>@�l�w�  �h���M�S.��Ϻ0�̠�:�C����K�`�
ģ�c�鉑��t*�K�ț��a��Jeϲ���D�K�j�M_r�t޹��h��l0��{��ӲSŌn]����M�B���bV�I���d�rJ���/֨�ӯ�t���'�m�� M��h͌��7��0��o�ف!D×�8:0�1�٩��#���a�����w3�kXnba����}Y�b�ikSib!E5(��˒���иH�&���H:�Da�,jB�$(m�TP���2�����
h1Z��h��F�����Y1�6��t�ݙz�O���s���F� ����#�`ܢ��B(���W2�l0t����뗙 �oc�N���*�\)i�0�e��tA�ga��Hf
iM���}��X����-�rI�MG��)�-���h�b��dunrҢ){� �>���v�E^O˴)�J<�8LPsz���2����ή���b�K�{�%���t"v��$h����=�D4^��ɜ�W%d.(K��-M�g,����r���Ͼ%i/�N�2��ė�&�;�����J�Ĳ���{�-���>sn����;����vz�����/ݵ�����.���)��&�	A
����a�w�b��^���3��]����L�p�-�)����� #�iy�����*_���	�hc�}O&&dR!P=�&r���x�})�Mэ��D�[�L��Y�Z��YM8*#A
V�R�cWW�#�=ʚ����u��x��U����)�ަ�.T��`��K��	� t��Q��k�����ha����!����L���ʄ�W�QXva�!��jc誙Ë!�6�	Ü��ʺ4�ϖ���n��.� �֙��ސ�V�s�*���r��a����`)`���<���k�$+��������m�1b���N�i��N�9_�-�L��꥜"W�.��ԉ�6k�'��
|6��n0��9,��{���R�z�΢J__�K��#�3S+۬�Ě�*�R�-(��GC=aj��f阭�+c��&X���ʟ�+]wSU�n"�j��&�� �(pc�ĉ�� [��Ť�`��J�.��H!\��7���QX)|�u�Y���h����Uk����(�B��V���Kd�J,�{i3��hw��f8Sc�H��l��r�;қ��#������f������2~z���dy���´������?���|����C�_y韨������������DL�j�Sm�Y䞘�d�^Y�@I��KD6uT*s-�S�S��#���� @k���=d�5#́+�F��muO
�J"F���a1�/Cc~�ya���47��EI=��9�Fq����c�@s��UC��j�z�\> ���3(��S^�C�ZE7N�1b�ܡϢ��&�*8�,)�G�E$��ZĻr�h��T�&ΚGŖ"�BR�K�H��Ղ){;�bk��eܾ�r�L���9�^�1�e�M�6K75[�
E3��Y��*
J����� �r��}�t7.[ʭB5k�/t�]���&���׉}G���w���[����%"��Я�TmJ�y��.V a�d����T�=YM��'��BS�$x��K�kJ�b��Y^U��f�^��̈́VߓE|������}�� �Eq���'o��ƒ�]���AB�v8��Z�_W^)�d��X�i���w��}kɐ��kx��߸)��W��ˎk<����5�9���G����^�����_�ly�����߲,z�/|�SG:�>���o�����/|�7����8>~������~z�l��e��pJ�LC-��ՈnW�P|����)r�K�|F�J��QN3�&Gi7�g͡�(�h�Sr,�6 ����!��|��Y/EMWa- �� �v�ficC��L]o�,�C˯��`�IB�dV��B�o���F�(�Z�M��(6�b5���M���7F���mi3��)�Ѽ^ete��޵��yf�0�>�l|�JᑠЌd�?W��3��Z�ϊ��w���`r�kJ���++"����8����׎5#�����=�z��@d�4�&�w�L��@@�Y/2��g`��,���2��1���Ю��l,G��ަ��\��dX�FBk�pt�+t���c�u5wnZiOc��1�����X����o}~�V��T\�������`�������F��Z�� �.�::
5Ñ�jJ�+��� \�rc���]�]���E�Y�,�b�WǮ���Z����P��f���|w����m-� ,��g�(r�܉}Y�����s�Z�����^��=���u��|������ }����;��a,��ȯГ����ϧ�������ku����������O~O�,�i6K��e<�G=c9��SMkU����I�TS���:yw�D-o�Qt�k�P!#�x}_�O"���,�^&Q�o4� �����'�@�=.
�=$D0v�3L���)-�+p�(#G�v�pDc�9ԯ�F$���1	�I�9��c�c�}����>[(��Օ��&�p��%��!I=kf荎3�	w֮5fuꦝXl�ᰴ\�`�J�|���g�'2�NG���|���Í.���#k}< ��K�^��+]E�mfkG�'f.\5���8Rb')|��pL\��vݹR"��2'L���V����nF�c�}صG`,#��m���k��+���x�� ��8�L�����b�cƠ�������;�����x�ީ�F~<�S{r���XV���Y�9:5b/�����|�`
|��F��5}�v��K���)��w�a�=JzM`���$�o�����4醦k�#_�:��{���\�S�b�m�n�e��7�G/�n���ۻG����O~����������>�iǝ����������K�ŗ��w��{~�/����ѿs��{>>��O��ߋTί� �`'��
z()aM)f�S�lf_  �IDAT��g5�Iw�"����.����~B�����n:Of,NhJD�n�ɣ���y��m ��Q�QW~���VL��]�&� Ƴ���OV����X
����ؤ�ƈ@�hJ�q7X�ð{�`�1�>;�D���[�_|��HCp(	�ڒY����i.��ťЊ�&�-�\<��|���GP�������?��-WU��zT�Kn�5!�f�Yg�0{ ��ī��Xc�4s#'.�J�hoO��u��UgzN+1^ujfAW�iǶ\��U7G�tG8��=�K��3�5C��ٖ�p��|4{�O�Uva�];�����:s�Z�m�:��������ߏ�t~�x�f~������vh�8��ą0�n�h};:Ȩ����
���~��]J��kCBĕ�| m��vzp}ש#��:9Cww�Bj�h���5s6�/R7�f�N�{U+z5Y��y��Go��������������G?���;�&�e�_W��<z����w��^����������O�W~�<����/��G�_)��Tc�d�������v��J�~�Z�������,�O͂!� ���ݸ$.lZ{`H}��k����M�7~��S�p5]E$~�R��q^$>lTj�4t��},&�M/���cg�� ��Γd�y�MC3��:�[E���ta	X\�'�׸n}Ctd�-��	�1o��d��lo��0'%��2�tJB�cq&$���:Y�.��g�w�=�R�\��+!q�.Dmb�y?z��P�����$�(���T�O��}�$�l�1x�~2��rP�����V�-d�1��KORT�4��9R0T��s��-k��#�&)�Y	���kF�2�ofNb��<��Z�V8,V�K|f�H;�ȳ�Z��v�T���۬�<�\�?��~@݉��hF���B�{8	5�1V$���d���z�ƴ����x!̇tm��I-����$�Y,����S�0t���z8#������KQ�Eh�����s�pw�܏������/���Gw��k������6���_��w����g��G�^����Ͽ�ߛizy��Ov�ףE�.��� K*&�����:�y,:�W�ڣ9����k����ڡs �a^s+��n;�"�)ļtiM3��q.&R.��*l���l:k��C4����~�JP�Y�L�lC%AgRdҪ\E��j���;5'��-�ᬱ�m�u�k�(]�H{%sN���W��X�������r��u����z�Q�g���.D5E6���d��VO�W��e���s<�vN������F��v��;��1�� ��,L�̂��*u���ي�4�;L�\ϟ�>�XA+]�~~M3�e�]�JL��#��A��G��I�f~~J�t/=�%���'��{�}��$fQ�M1�OE�7	���!Q�����"-p�Si�Ji��\Z�i��.���6�� ȣ��;�]���#pB1h�U�Bݬ��*H�i�R��@%W&�s���Ȓ�uGf.L@��HV���R�f.M	,��Q�?BQ��|/����	��ۡ��^�YJ��U&""0))5�vW>����m�}��1��d�X3�u������
���*t��7��<S�4M�,%R9P���Vn�L�^�Ӈ��?��w������"��]�NO9��p����_(����z��s��>|x�~���n�����ҝj�&Nt�sa���"���Q7T4�X#- C�'��{����с�\�8�!R۱����5�^F�f��:@��IkMSǇ�RH����?xM��I|�IC3Sd1IQk�G�#��� j�.&eڒ"J�dݐR-%��k���ՋWA܈Q�����2��klנEj����:�b�b.k��Q#�81u]ߢ��o�ϵ���U3?��%Bh�ᒶ0_qk����u� A���5�ɖ��=闿�4[[Q��Fi����S� �	e���
|�<N�1@�C͊�.p�!� ~G�V0#~Քͱe|��q��5�$�q6�\1�㌏�Z�@�F�?�nF�g��@�K)xZbipuh3�֭5%���ZӘ��9��-_yjxl�� !H`��?�րhE�f����ᭉPJ���1�6�С�5&5ܪv�����VN{Rf4X,I�0�i�0	=6��iz��I�)ڡ�����	!�@����x���Zlr�/��a�Ь�_>	]%�+�����&z[D
E��R���l�H�W71<T'LVYꈣ������+�ԥ-���i���Q43F��X���=���OM�y��:�g>�~���O��k�鹷��:d�8��>�������~��5���O�1=m�y~\����ߞ�ﺩߐ	��w��,��� �p��$,5�2@׊^\f֢e����g}�������J�h�*�m�}ۯf��6j\+���`�������@=6�1�QZ�)o@����J���gG餡�1i3QHڄe�� x�!�����e }��^��;��H�Ecl-��w���D,J���FkM*[a4ʝ��{/r�N��H�2H��O�T������k0(onIa� #1�Q��o��a�;������CѾ���y�̤��ᴚ�UH���E�F�iRw��� +
d- B��t-䦾ah�b�# �Ǘb��R�`�Ó�Ǝ�\���X�X�fB�Č{��/�ܩ��*f����q���|Uw�y>/�dc̋y:6m���T(n�ڒ Fi��Y����]�зaC��[×L�#��b����XX���Xp����0�W��Fs�?��x�b������%��'kv�BQBê�@-jYU3��F7���g���^����C�����ߩ���7җ:^C���oz}���ɀ�������ٟ��O�/�щ��H�R���=�������"�nT-i�IT�匉���V̵����+��4f�Nk9�+9��>�i�d�#/4 �h�C�ޑ� ��mL���;(X��77fiOp�}��E�V�
���I��T�Ĥ1��,n�vf�@�B����2UY��'ن�I\Q�z59�7�5���T�l�#��0.3���b<���ML�,�8�U�9��E�@Y��ςQ��^���\0���p����=^C�~6�{q!�}�E�we\�;7�IE!Ŧ�J��s�2؉f3Uc��kK�����cMW4����s|u>�W���]���9hQN���ؕ~����i�Nu�I���`6٣v����,Z$��F`�lX�S|�M��s�ék~t�����V�`����@�]s�X��8.�R:�]	0�Ep�(�Q���횬�ӊ��ȍ�!Q��DN�Oy�N"�Ռ>�^�ʟ$�د�o\lf�;����<�>��˳?�v�oz������:�[g�>��?~��k��2л��}>���i-�f1��TC�z�F��Pr�~SSx��Q'�_�xH0����7,�M��%�/�x���e8Gir�IA��\gу�/�<l��5�Y`���fj	��W1̩��,37I��A�Z���cs�S�V�ӱ'7��6@�Da�S�����
���Ip(��-a��,�:fs7��P�I�'����i>_�n�Z�L硦I�g�+�,&!�#�%����D���,*>rBк�׀Y���d���@(�N�q������dt�
�}�n���P����z�I�'�ps��ijB�z㳭���IM��OZ�L��zeܰ�oY�΁o[���täj���CCW�>�WL�M��<� �{@�a��%��!��0�4�\�FPW`�'�f���Y���݅���?`JҽѮ���)�?�o�U��l�v��-[���
��nM!��@���4"+N�Ч1IM�L��f���;�\�OЭ|/G�=���n���=�=�C���g��7�����_6C�C����I���?�������֟_&����ā2��e�`>LA�c��:pJ�%��޴i@�8Q����&�-d�i����9u�C'����m�C��(�o�.��R��8��c6���U��{�,����TB�NV���"r�t[��O0td����Է��o�2���<L�SM�8J�@*����m��a���!
��1l�f�~:�ܕ�ZE-k˫���7����"<3WL��\K!2֪�q�*�P�>������,2���MƑ�#������`¶���j���4JKYq&�;ES���v�Zz1f%��
@���&"�;?w��`Cv��``��6'�vu��Cp8����o^�^�ԇ1��Y7˷�׮9Z���C8h"�O��B�ե��MJ�	ꬁ�]�i���X��d�v���ԍ��{Pm����?��xu
�`>���'���[Ҟ&M�U7��a��ٝW�ػk�!u�Q����bj�IT{�b2e����VUek2��9�O�~u����������������=�A_��1t��L�����������G�y�"]/W���il�1��räѱ�-_�,
�{���j�U���Q3$\1���Ř�^��h�� 08|>p�6"u&!\2t%�-��͂�ҹn�p���DCԠ�b�E2ӽ0r[t5B1������D�+C`�L�&P��0�*��60A�������10�����h�n��y��LxXKb��Q�g���D��mg��ee��jD��n^76��6Ĉ1@M�]5Jd;���f�ւ j��o�1�J����t�c
�'��/�|��{�#�@��f�p�n�-�F��z'ʹ\��]Ts��ߌ�Iz���&�Ɔ0bxk>�f�o1�/q��;��ۥС�6���P��oԎA�v�����|Q�K�A��Q�z��s��+Vt�3����oi5���m��K1���K�Ef��qF�Gky6���P3����ڄ��j�mX" �r��Y��	�Xm#���;oy-�tH#�Hb���k>�NR����3��^x��V�[���1}��W��_��o��~�7���������ߟ��N���6k�/J���mJ���MӰ �K�D7r��Wgէ�J��ɺ6f��ߊ���p�s>J�w��-��"��<�a�q�2I�H+#/�����̌��hT`�v%2�XȋuSmb&"��l̤�6�k�(I���+��L?�a��&cj���͎��V�
ps��������p4����[)&��)���=������Ka��*��l�V��No��VB%4��"�=�����C�}ݛ��U��a[~?꠩�F6���v�g�B�
Ke0'�ܲIX��Y*��խ�\�F]��^;pM��M���m2ʎ`Ä¼2�����^�������;�ay�!�3q�KL�Y��� Df
�2��|G|�>!�Ä��}S{7��q�a5C(1q��	h,;�oґ˃2܆���"l)�`I*ˑ1�*Q�2�Ɉ`�6�X_��h;�$(/F�{�)��U!��4���YXҒP�ߓ��_��~!4��h����[Bk7���%hV��$���>�^������Sf��,�
#7�����x���o�����=����ߚ���羚���:o\���?�K���_�7���~�����>�C�\�ʽ\��iX�{�\R�J�#m8 ��@tf�B��`� �Vw�bC,�%�m�����6�(��Tb�3V�}��A:/�.k)w�
Y���jK��<Ka'<�jlk���]b��k)Iz��w�7n�`�_�ّ���ݘ:L�	��6���Q(�*��Ã1� ٭!A�y]�y<݈��~_�z��}��r�''��6�G4[`u��fF�0W��veR�l0h�>�����9T��1$s�H���mV<�HB ��f�S#B��`f�IV�5�
x((���� k��V%w*�����Z�ō����JW5#����_,E�TP1��1<k��.�by]z��]�x���g�}dV�i��{�!)��3�'�V׀h�f�h���;�.������{�l��*X��[:O&�j��J!Dv�N��MZ[�|��i�'��M�G�8U+��!*5Ł39����=�6U�90ԒR0��S��Ҧ}&8%��
y<��L�"(�`�Y���U�
�M�?4�u�⸞�	Ӹ�&r�y@��(z�Vt��x��έ����H�;��ŏ:���ED96L�nZ���w����������5o������5�����_C�����z��O�'?�y�腿���]���G���܎sq�KL�yqgʦ�)�}U�wVBքZe"�.`b�ǖ_l������}�#��ĭ����3�0.-ia.����@��'���(��*�B`�Ʋ?/����H�5k����K�t�K�)^��v2f��Q�`�Ed}(�i�6�kƗX����9>��^e�nY<�8��Y��M�x��)SŰ�#j5`�I����h��c\v�m����ʅt������p-(�^3tנ$�:>y'01�ca�����\(�7��/�Z��y��b9SS�\��jvlpE���.�>�	����/�X���t��������!0[�c>>U�K�4�Ӡ,�;���Ǒa��ʐb�S�s	����7�^E��o��c'q�Χ#u�~��[4�t�e�����g��3"��qpl�)�-h ,��t{3�^��w4�بiaӅ���5C�
wF^�/�C�>F�_��%>a']��X�ئ�ۻ)��n~����_�����"����M�����_5CǄ?��.s|��ͣg���6��ϧ�_��!<�)� ��ԏ���R��TȂ�	ȩCW�cD�w�,J��60^��͕���\j3����B����A��#u3V�A\g�cH��ƶ�t&�e�Y�0�cR5� �u���cU)����ѻ܆�������S�J��:��!��]�O07b< D�M�[�Q�fŵ="�R�$w��~��̟��:4+�Z5�Rc	!I��vhx�
M�,�Y�w�.��J �0��)��B�pu����3��iU%(�W&��Uh"+��1Ɋ�_+n�"�ۙ[�.�4�IN5�Ά03�q��H f�k��
<�1	6��s���-=	������ɴ�&U��QH�)�����v� ]�����J� ��kB~�:��O��.����"�h�)M�L�0�A�����݂˧e��'�������H���Ee�is�=�t'R �僀���lЙ1�9;�1?T��C����T/�Ǻ\��99~-$�Sq+���_+<;K��b.��j謼�ɓ�c�l�s������?�����ߥ��7�����:���������2��������M��{��������H�'���f��,_��^"��s�	�(�֦Qded�@��ȍ8ۙF�bѲ��D�m���AW��m�m;'"���#i��@��PQ+���6NaV��b�(��m�֛����΁7��L�	�/$\̳��:%�6��.];hB_���'��}����T�x>��k���C?r�5#�n�%/L���I���Oi3a��A��I��T�;�VZ������f~J�	�ȵV�閒��	m�Y*2�5�f{J��Z����z�����9�Y<�;���i-v���8��R���(Ym�|�ҸV]/eǈ��G�@�3�����k�,�W�>u�̓�lM<�u����
M\�jc��9Z����1���ʭ[#aM�X]9Z�%aZV����<����Z�t�óM_q���"��#N8�����Y����'����4[@"��Ѹǻ�Ňj��� 5k���A�����2�c-d\3ů�E e���{C��of~#���'<M��q\�^��u�dw��ov��S����
�������1t>�������L��l�(��"�}S�@D̈� Dbt9�t׵��g)g>�ɧ��D����?��f��g����>Pd���+���F��pO��5nb;ɾBP� ��Kmq��L�a���b=0^����k���}���ǤxEW�>��H�3�Ey��`͑�tiMd]֓��¶��6�гb�P�<��qٜ�g�{z�����ip� ��a~_��Z���.\'��%|�� !�U����Y�2�Ԅ!�\�"�j�L��@dR���B�+��"��#{j�v�&����R�=N;��D�b��G���GS��0g�a�}�����SR錉�B��]��UK�S�S�紕i��c'½D]��I��nF�+x����I6C����\1��[�E��2�XO�A8u����Si�hV�ЧJ�����V^Եҥ��N�m�O��|�zsG����r�|�s�f!��ZD�!�S��,|f����.��b6K~?���|)��n�Y���|X���[�â��q�kDγ�<��Ks���A���s�ɝ(.ӧÂއ�����{;�r��oz}���)C����>-ƾ����8�;���TΏ4��[k�F0pt 1�����Q�ś-W������8��f�&M�j�(�����ơL��f�	���2	�~͐2qE|��DZ6Q�t�Q��%�EY{00�����inBk�o����0+�� ��1mŉ��W����6�J�q'��䫣d�YC}|���N�'Ҟ�0�v0�Ƒ�������K��2t-�%�a*$g�U�J�-��X�و��{H�pa�L�O�s�u#TEK�� -_�������5a��j����S�9��M+V�����p'V��D��|gBC��T�Uf��:Y�o�&�U0�V#��:N��s*lI�!ÿJ�ݰO3�L@�@`�"�S2�,:}�}���(��([C�a��1���0�mY���Ь@�f;0��c8o��>�f�^��*��.�}���Oď���t���p�Q���+�8&��
du��1
ݛ���	�C��G|�y�=�9մV���3Y�x�k+怏k���A��g13��i����m�BE[�rN:��-L�c���ͧ���=��.�}}|���}����?�n���v�?Q{��K9�!�3�Y4@m�v�ཆ��{�Qw[��Q�U�-��w�`<H��8�(�"R"��R��������e��d6%x�>C�
�o����f�V[�ig.��k}����^}i��x�7R�T��D�:�r� ;2eQ��T�m���4�I���v{���檀I0(���*�����XCkp��nH���i�
Y%�CXh�5Ba��Q�0�G[�3��w�CۣRCohn�RI�<I�O&���H�p��	PY���	�ac�L�`�HeC%:���P	8��M�#zc��N�p�'�q��`�VŃ��3��q�b��pd�EYΘf�{0�UaN4=��������If�]�Me����@`][���f=�S��H����w��%��%ѭ=�JZ�@�%~�n7E��?
0i��u�%lK���gV����)֏�٘��d'��
�0�ݣg��V�==y�%:��[�ᶉ5�YbEK�J���\�
��!�A����%�3��y�����9bs�L��Εv��z����[�9�i��i�)���3���Ci3wQc�p[��R�k��s�Wf��/N��?t��}���\��ks|�:�}�{���W�m�;_�Ŀ�����w,0�6��=�I�ڮRK桐�.q����t#O�r��T�j�#u#��:��I��%��,��&���m =f���0\#@��^C�2�3n��K����kE� ��tO�*V�cWn����R;�?�ӱ�,fR6�I��pMflf�-���+o�Ό��m3��0�4>�{:������r�tKu���l���TV��:��U9Y�C0q.}7�RNU|�'6AΓ�z'��_�8�g��*�˳�
d�S��'*�)�l$��������S�#H�Qr�F|%N�g�
 '֬8#_i�|ޝ�)��	a���5�n���k��
8�΍=8��,=���Ls!d�R);��rLիL�p4ۺϊ��!P��=�2������q��v��CA-DbL��#�{�GE�o�_��.����uy3W�=f��Y�UF^�Q�0��*=\���~6�U�R��|RZ����0ef ��TA0f�x�v�qz9��nXC\��x�1~A���,��%ca������ځfX�-+��|�`�#��d?8#݄�ȯ��͚�?�x�����P.K]��+���iv*�V�OlO���R�2AT�a)g�����5��.�S��p�C��sLVN��v�s�wg��_�}�����6��-��ua�||�'~����t���������~�·g�� _�j`@�fJ��ZE*�4m6 >�3���&��oVŝ��~Bp��^��]@4��/fu��� ����m������m:Q�r6Q�"��?⮠��Y���gL��F���Y�0�Q��I�Ed����H��[�WG 3��0� ��i��/����FR�%D�<V�Of�QF��n������y5�����pAȨ3sumn:����d�n�>����||�Z�M��)�, Z�����E!Pj��)e����j(�,G�PX3:/�5�{�b:H�Ct0t(m=�'�����T-�\��F�Z[b�0_g���Ws|5G��P�	f�Kn�����,�Y=��$�3�G\�~-�u^5O�7y��\��=�A^�I}��0�P��=�Wr�f���๾��4G�x�px ^���+���$Ѡ\�,��X��v��J�����Z=�MȪ�0�\�}��R1g�@3�7����"@����E[��G��?�����{/}=��C����P}�S�8�����X��?N���ʵ�HL�����b�J��˻���$9��Y]�ޡ]���/�	�R�ȓ�Z��k]�Nc͓u�Z ��M\�Gjc�ƈ� ͚�G�	�`�\þ�s����̆ȳG��eW��-����d�r�t\�3�fib?��0���%y.�Z�j钺�5�y���6���*���Q*�b�B�y˒�
b~Nu��eGb�֔���*���<\�}���2�����9
#����}�%��|�<m\��Si�e��oi�hD\3f�p	Z:=pd�G��%����A���T�ӓ�z��&���"�Y��n��#�Q�fe�K�:��[D�2z3�'���Xm)�]�G�Q�"����֝2Xg`����ڱ��f-]_�kꭅ@�`7��>h�aɪF3�b
c��`������Hy[q˙/voע��J?�������o���3�d&��!����W��0��v߸�g[�֣]��D35R�4ձ\��]@��!/}>2S^j������Z���]��ښ ��/��b��[�����eg&�I�y�y\��4�o~�q��~�;�z_7�����E^{�����ӟ|�����g�N�������X�}���v̱v�<�V@�f����"9��];.��f�`�=cK1G`���c����_�z'��[I�d�.��4�ۂ�-�(�gT`�t{�;r6%��h4�B�OR�+n݊)O
�q��YL��y4�F��3CKU��'G�;hu���Cw�;�]���5�D%m4א,������M����س�|^���Y[��.��*~x^㳚yĬ6�J�V�ִg�'8�v8k���U��1�;_�Å@�a��$GF�K�{�w�4\�6�93��L"���)���M�i�s���2�Oiw<��]:$�`c����nX�҆E�>W�f�K�W�X�D�yM �$�$��-.8f�{u�|�̔��	-\!&�Z�jw�x64ʊ)��SZ1��"p�E�Ͼ `����87F�,"|5�:��,{�M�z�h�����(��̻X�͒k��0
O(T�4ǣtZ���JWi��f%�3�kʶ���
r��.J�y`�9�Iig��l���F8p����O��}.���ϫ2re��7'�s����8M����Ox_��}_]񘇎�C������::<��/�O|��,���/0y�DS�E󛔉��=�c�EtJ*�1����̻#4��Gf�L�LIׂy㛮G%�&Q4����iP.�i��3Af.K���׌�ivS1%D�	I�H���,�Nz!릉b#͢��_��!�Z�����"��Ԛ��k/�L��][��v7�4B�Eb�=�w��/w��)��ر�&�[��=�o�ŧ}y�c�&!�g���|߽N���Fʭ(%9@l�bG��F�Y��c.Zꘉ��@�o���5G*C��`d��B�^J䑩)�
`(д
�,�)��՗Xw�f��"k3oO�.r�I;���j!�����%B�n�\<�a����v�ϼ���_�9m}�͵%�'�B�3_=3�:�U&�P�T�G׽�﹒P�q�_�ԃD��^ph�M�5����pĻ2k)�k�iU<��������N,��}��$�a.<s�Jr|kf斁$�M�1�K�}V�h.��n�..]�b{�\];ZB[�52z-��5�"]�!v�D=����ۚ�#xSt|/��$o�q���}е"���w���[��_�}��g���������3�R��>����t��}�//J�?�H��R�6�3i�M+�RA��Q�����s�F��fk�SB��؄>�G)]��`� vg�N��!���\Ւ4�˝��s���o@���cD��,&�&���>Z\��L>�S�N�����izM���%Z��N��E���~9!�
�D9k�V�����bN:��&K%�5���y�:�����8C�p�NF؏`h%�L�5i���qa�e�ιj�^��5�Zj�Ko��_34�/��n���ay���[xҠ$>9Yh'n�"��E3R*�<��!�s�.0�R��dx�H�L�"f�L�ʑ	�:��O�[E5��{*˟��L0�*��L�j�T_g��Qj�]C�u�9�k�m!�^|���-���|�}LAM8�0������&v���I>��*��}��ձ��5@��OӀ˩@���\I�2k�糬A� (-�Z �)�"]�drT�'�vՒp�]q��5 C�V�����
N���"\#:6�)Z�~3����I�j��H��\4t,U��,�gv�pB�dM��#��@�jQ����V���1H�-���N�/.~��ܻ�����}|4t��������ş{qz���D���$��-�XU.� GD�FeMY4SmɝSM�J��ҧ��C���������MߏRY�D��s:5�_CWd��&6Yw%��tj�5T�`��BFLͤ�L�DÔF#]��{��'VN�d�U��$�4���H1I��G"��W�)Ҍ��_K��:�=�o黑�g�/����ߙ/ lMza����r�+�N_�h�Yk�kᜪp,��Hk�kmr��n&z�k���Z�������))?w�㒯���_���:h���'ZI�Mx�hc����7v�:`����nfo��	ڟa�Yk��\[*x*^�d��3��K׸��߰劥B�࡙vW��/[��p�I&B���f��%r��j�����Aq�!�zt嬸`Z ����w��$�Dd"��A+��O��#������-V�C -b=��鄈�"��8'����}�-��S��K�d��R"������22��� H��pݰ���/.�qf��ƥA�a����O��M+�V����1;������gir�z�X.�����H�����u`�nu���d
*ǁд��e#��/�އ���g�������7�����}��׿�)��*��o,���K;�-��0Aʓz�E����),i��Q�U[*�O{������� ��9�y��2�g�G�jM�0�5jRDF!F=�$8�g�5�,��u�!;I��c;�=K�b{�!i�2�RLL���;2��Y��$�$T�V#vB�w��Y>8p�� �SW��ޡ�[�Xl���<X�����a��U�p� x���g!/%*_������ŭ �U�[̘�ҹ�~��+mO/�G���'^N�-4��h��nγfV����wt{7��e� z�	��y��L��L7�I
�D�8��d3�a�B������T��ا��}�@D��N�ST��.m��%H�8��H{�K����r����'Rⶋ�{'- ���t��]?�᧍K�!����@�
��ʙ#�#荿�&8�>�8$m���_�yˉ�մ�N.0�P^,�ք
��kB_��4b#T�fݭX�#��'��1Ip��N��c}�R=��l�d�"���3gr!����e,su!D��X���Ҡ�.A�Uc-��BK��-VDr���p��8W2�Z�L"R^�ޭ%\w�B�e��5�\Cg`t��[
�eAA!P!sf�������<Оb�#1#��ig�G�'�������4E�8}�n�u����������}��7����7����o����/3�N��ۿ���=�����0	2GB�?�(��E" �����������]�V���t���F:�(��V�{W6���U�Q���5k�y��M���r��|����>N�G	�	]h����NBT�@¡^�E'���^�}�������*��q�C�M�B����&�}��@v]�u��'^$S��s�W�@B�+
�d�t'1\N� ����<=��i!
;�/���O�C?�u�_g@I	�Bjs�� [���c�UP�&������ih��Z��* ��@:�z����K��X`B�^���F�k��ɛ�(���V Ø�"���ڔ룖^���S��C�)����������Z���~/׼U��4�5?{��1��'�́������*�t�+�؃��1�$9���.Y�d��X.gv�
�LښS`׺��Z/<b\��ي�0=�ׂP���r �K�,2#�fP9�ߔ�����0�{%���Y�nD1Edx>Y��B��y�
�Z�����iO�u�D!�s�mvߦ���Z�)]p#I5��h�<W�[�w����ǥ���ݳo�������K�:�a��o���/�������O�6�w!i�נ��Y|�-Ȍ=��b�^���AcQ��ms��I���ދRw�����Tb3wՒ:�lML*�eb����M�JLE��lr?qj�4�>��礔_%jKC��jJ\�gl��{��/����)�Q��l׶��[�����ݴJ9jh�q���}��oK�}��z�dF��ˁ�!̳ᓦ��F~����j�F'��!���7R��1ccT|镧�7ӳ��1͂˞jP�k����,n�Yq�~�� �~v�^)��'X�6���s���^"^K�B��E�;׺ꤘÂ�q�̟<a�F�ŒYe�ZDLr��2a�#z�](�&���|����M��YK�1
�B��;k͌�%���ZDB�X;�
:�w��}T��k�ɘ���'�I�U��?[$H-�p���l�?��Q�~�<��$�q�<Dk4�D�Jv�-B��p��� �{+�{М���͸�T=��-{�,{j�Bռ�Lڮjt`�5פGk&�=UXơN��w,)n�Z���bL�:��8U��T_oj�f��A��&�ql��N7���~wf�������u|C:ǧO�4�~��{�������L*��*�`�~�چn�j@���_��i}��FV�k;%dv�L)�M1���-`fi�7H��Y��\I)�j(I`DQTD�I��J�fM�$�eA���⤂�"�l�p�L��$3�j�j1�r)p��km�#��!$�c�5q?i6QTS9�E��1c�n�K�%u�;��[:;�BO8��o��bm����yY�����NZ�hR)R��J م�"���H����/}�C
��>81P��c-ڠ(�N'H��I[I�ڮʖDR2EʒxI�rxn{���c���9�>�v�P�����������6p���{䁅*�%v*-K-�8]/����i��yj}a��8��|o]�S
�H����oJGٺ.�
�̊���@����8Ѿ�F:	�?�?��fQ�$��⮒�EU�7��U.u�$��\���
��[���bN�������>{7�tyy��q&׬�r��2�I[�g�}$ga�I�5��X�ܽ��z���z�e･+�I{#���lU+�L���I��N�dn1�ų�	t�䦊�x
nM��}O�N���@����r����V�͓b�,2��d�9�H���t�7)/���m�ˈn�n�]�D�F�A��)!���Px������h��"��+�~�?�4� �'��y����������n�O�A~,&s[��w��dBD+���4�Wn&�MB�}6�-�{�h��]���C�L5C�u��z���Z�ZNb�Y��X�z��+O�ɜnЄ0����4Z�����U�@��H�ĭ����._Q�	@�y�:��O�����d'($Fb����u�

H�J"X���&&v�21K��>Z��%,i��h�4deG�5��"��X��j����U����8^w!;i�u� ��Sb�Wtʲ�\精JHaz?�'��(��,V�Q8j8��u�\/�e��B���}�FoA�{/)M���uy|i"e[G�vV���1�:�˾�7Eb�<���)E)�����v#��_���ngF�SI�i�{w�%���c�9�3���8ȥ������ᾍYdB�> V����F�S�dI�%i�z��}(�^��ۼt\�Nי5��Uw�<�{�MV�F���Q���LY�<��k6�����)M����\�8^���Q+rg���B��F�$#��JkΣ(��P�B��wx���.V_�����ӊ�?pB'�'��7^�*�ůB��O��?�~�N:�ѠxH��LN���d�0�۠��Sk�֛��	фɁ_�m��[�w\�a
�/�5�sL	��U]�l��?|ә�y�=5�� =tlY}y������U��8Ȫd���7����RӜ'ʲb�m����� ���N[J���3N�q��e{\(�
�����-��.�� ��I��J��A�}�)���Q���[�Î��1QԣA-dxn	)A5��IEI3W�t�)M�+
����-kz�:�ߧ��TASr�͕9�9ۃA��%��S�K�����\Z<nO*�Q���qF�VS�q<K;h����'���0.!�>�s%��� �D������a� 푄�a
yk�"H:@�*d?�"��9Y�B���lѰ��>"���z�N�ٜ��JsOeM4o>���9g��8�@c:�%�n��_S�̔
j(�ݍ�N{�ŵ�?X�w_�L�����}ʫh���?��Q	�9�I��4'ɔ1��ߧv��Gg`Xf�D$�ͳ
lO��{��a����lK��(Qc��$5)_��n ��kxS�e��5���!t�=�~������o)�X��?�J�>Є�*k7*s�)���%i���YJ���þ}:�>J�B�Ek�czH���Ff)���cL泿��!�q+wV!�	���ロq1q��q3f�؅b`��$�`��K�,����Q�T��تC�Iq��T� M�&�ȣ����,�AW��W���e���1g�`ݷT9PT�c�O�)�4
�A�7oѲ��ER�+q��v��o��e��Ls�q��������Ш�ԉ�@ٳ�F=)6x�wܪXr,F�~�0��g6.���I�A	ko]�>��kLi�YQ0���Sᚵ$J�u�@����2��N�D��(��Q�%��8��t�����v��<���1������|�5{<k�C)c��Dnc�#�ȱ4�Ŕ�[�Ρܿ��i�HѫM��`-`����W(���u�"7H\�ŷ�7ރpR�K�\*�g}�S&����	ux[4H�wm`��]���םt/�̙�����X<02.��4�V_�Mv�c6�/����b�n�>���$��ae��b�P��U���^'�%�P�Q���<�`
k1� FS~4�F]Z��MAcE�ǟ��=r��4M
��܀f��������P�a���:'|`�~��	�q!�'�v_�+�[��<Aٳ)QRW�]�@kա���/�u�}����&�A���Xx�A+\&����ݪЊ���$�4`������ؠ*�#���s�=�O)���4!Y�H�If�/���8$�5Ťdnnv!�D��aP���:�>���2@��\S��4� ��,���0�Ʃ��3i���X	u��+���2�J�/�qԬ�՚����6lx�\"�J�4��u��{�D=>u��D�
[}�<��b�(;�^'��$�\�]�Xi�ѩ�P�>�����\l2O'c5iς�z�t���Z�I� O҃Q�X]�U��'�)
Z)#���R�i��|j@҉�d~y!(C:��.�j��Z�J���4�k��g����^"#á$4�^�2$��M}[#��"��Z�����T1���!�+٧�{'N?�Q�$J��ΥRB�����/�_ϼ��M����%���� 7'j�C����.M�Y.����d��d釪!��	���9Ú:�I�Pi=�`���n���z����r��PԖəȼ��M�|jSP����5-.�\�r^��FOTQpJ�zZA�����`�H��h�(fc�Sԁi��/7m�]�7q՛BcW7��P>��	�.b%��y�7�uiHC$O#S��]�z��[��?��6��p>(|`�~��'��?xN�����������/������%��k4��4;�R��u���ZtP�w�ԥ9�V�HW�m��-�؉Uez�޳�
T�2�%����B�Xד�K�Πپ ��]�6��"�k�l�$_T�G,/��`u�r��j��B�+�N��_"�Mq��e��k$�1�:j��
�zu�3]%:B�q?�@E��i��hh��R��,����C9�z�ht��w���,�ɿ��������ٚ�T�#!M�&b�k��GF#�?��y��zL��V�j�\_>+5�(n>�m��b���5��<zk&�s������j��zZ�8Ϙ�o�o�G`e1��wPWi��K��a}MQ*��Qq.��}KeX�m?*@�Xt���\��F�^�7�C�_�ە�\qF/�;9S���g{�ɮ�R�D%>kώ�[�|��Ǟ��'/*�{���L�V�Q��i(H]-�\��p	&y���:$�n'�+)�-Z�4G=������=y�
_�2s��G����ۓ��X���:��B�1��:�q��"<�7f�O=�0��<vz��&���ͮ���π�4��1.}��j/m_�p������k��%�L�>0B'<��S��+�.][�]S�]�����OQ:T}��]cMa����Y�(Y�Z��-y1�����"��ķ�<#��L��L�I���I��_�t���?�U~���X�t��˛�}�1W���u�l�V�е)��I�8&9e0�I�JcYY��4�����[�θNa,	+Bu�Շ�n-C-��� ��Ne�Z| ��B�6IR�n�� �}��5��8��	�C�~�n���>W�]��7�_A?�(Z�`��O�^��FnLS&ƾ�c�q�%Y\�j=��յ4��:����~�[(��V��H|��%��8���N�^�pe$ZM�0�� {
ְC���cix"�iw��̪_�{
�<e�:N��e�d+O��x&��a�TT�P� ���YH=���|-���SZ�Nd�(�V�9QԸ�疆I2��n#��	�.ԥ2�n����h`��9ю�� ���h��dD*]�Z�T:Fqx�����ܰ���u�Öd�'�/�C�S"���d� X��B?�0��U�I��yN�a�ӊ�d�T&��;�%kIn�!������ڻj�9�8�i'7;��?�����o���k�>�C�(G��J�߽ ���l�� ,��nH����D�Ik�w�ĸy�T ��-ɤ��tr-����Wj��q�2��r7��D>jז�P�B��L�畿퐗����f�J6��mD�k����)�
����&=�눦�Q�g:���K,�T�;W��Zƒu�*y"����(j�Y�d���;l��al�i���3+;�X�b��SB���fT렄��+D�[\�MGd�-c��zM�)4DN=�:�µkW����^�訞�]���BCB�
={�����2٫\��J�C���
�btn�Vl�5��k&d2Z���R��t��Iv�F�dL�Y�$o6uA�61W����qtM���K`&}>.��z�4�����$�Irc�׮�#7����o�K	VerkĲ�B�EY,���k�\��O�"�k*k������?v����:��+��8i���p�>�d�B�N��"�i��PO	e�kG6.{�D�+X,� �`�9�A.t�v��kR:j9������6Eɱ���魨���s�s�'�������],͵8�d�q�i�&���5���(��7��=.n�^�Z_��N1u"r�2����_=��~�������'�4|���	�ޏ^����B�^���m�����z�C!e A�8C�Aݕ*�6S�+����%n��'i�g�v�o�)Li���4� 
Q���=����UL�n���O(�>	O��R�M!(.�L�$�I6y�E�f�m`m�e�V��A]��]�J cR{����ikI��$ܭ�`��o$�\˙�� T�ݲe��V`�FژG%�j*�ز>o��EA���%t!Z�⑩$<n�Zq�ry]��%{�����{޹���1���1^�c����Z��b
�2OJ�(D��k�L����I,2�u#-����nl5=�P��"_�z��
��F��M��#���-N��սU��w��n�Jf1��K��[J�/���$��]�:�͖���uI�q�q��Ե%����I	��:�P\���Öm}�^��0	w�]��:%�5H����9M�
��V�e{ۄA�(PRIc2$g�+ٗ6���I�;�f���
�mu���� �$���s\C�O<{c*#\�48y'��;�Pb��佯_\ir��<�������JO������"�����c��(*��W7}��y�ik��ҵP��\/�;�LLCY��5W�<&�@�=��-Z��j���a�[5�p��>4>pB'<�ħ���/|.^x�~���zI�P%�[�LbKNj�ԅ��Z�dnVw|����Wvg����<����w�b�������a�&�=mz����h��cuS�W&tv�Ic��6�r���ꁐזNh|�A�.���V�-]�E
���dN������ř�
��o(Zn�Ĕ�Kָ|�X-ԥg�:%{������h�Z��������RU�f$Ƕ��$��VE!�Z��ΰ��޺��[W��`	yQ�+�ť�9�.�ҬC�#g�q�9UE��r�F��e�7�"5[Hc^ۣi|��w�w�o�dHw�J�.�����b�U��>���zdm�)��Lt�6I���w��MI\�r�)�����EnL�I�~t]��KhI��]���e���=mߕ.7����qE��5�/��A,�M�c#!�����+��1db�Y��}oϙ$�ir%-���ȺF�g�R�d�^�X��4��%��j��[�2��J'��E� �ܔ3= hY��y��~Sh�v�D{496���e6�^�vN8�������d����R��-yF�{o!ç��ͪ��+P��ȍ�̓*�ҵ�*8�r:��.�N��H�i��6�'c�������h���gӪY��>l?��Ϫ�i���\�Ąb��b[/�<
Mj,������<����3w�~�����a�o�2峏6���F尫D���SM9�� ���q���zCɌ�E�#���t��r�*�q�6h�t��l.t��;V���h�L,���Ժ���
eC�3VHS�2�e�A�K7Y�l�z�'�$▭:\�t8C�$��"�r��YZ��O������vKB�*'Ȓok�|���j���a��i�ꦂ&�˔��C�ʁb!�l�,�(<CIpl�I��m�`�ض�H��v�q|��K��d��}�\�J�7:ɫ��B&���}D���S�4�;���ico9K:�V��J�l���<'�*X�ps�ۚ���w�I��&ɘ4;��Awj9�b:=���uP�>s�3���Q�;��d	�Akι�� #Q9+�:��\�g���T@B��F�ޓ*��B�_	+�*W��h�R̝���w,h�"�9,�q�e��gQ�s	C��v�AP~�m�?/疔���e��NVr��2[�{2B >�l�wFA� �7��e/Fk ��|�z9[�q����������:���Q�]p[�]�?�{����U\�_�}/j�U�6r���q��R�f�Rc�,�#��S��'�`ԺWM ���qSw��Q#ڸ�ޔ���12G�0nA�,���1�F��t#�c,�O�Af`%���d�Z�a��*h��J���?N����(2�%���C`"��ǂ��A�(d�1-�k�o��*Q��@<RJ�5����2c�E��aD~h. U)��U��N�
��.���O����f1�%]��C��=Z�в[��v�I��$Yk�4��n����bm�w:�U�B��f1�������a�8��xC�ߏ�	V��ٖ��9�bR��7��ra�1��0�kѪY�屧,[�+7���J�ܼ9�v�ބJb�9�װr�a�Z�,q݁�A�YQ�4' J�'ae�K!�J˱����K��(��#4�Xs�A`K��^U[�vtTN'�9�i��`����,��M�=@�[2[��)%�(M�,�n�*T���AW��ؔ� qd���hb]R�@�pJR۱�T/��хp��H���Cc�����a&e��"��5OĿ�mВ_�K�*]$�x�h.: ���:c�)6�K��PuU��?W;O���n�M\Vc�xI4�ڋ"bJ��f�Tʂ��U�^�0Q�V�|F|N*9?�9Y�0&}N���^7-W�C���R�Zr�/�/��������gg�����n'�V�N���O�+_�2����E��e\��qH���&+I��<��~�Lw*��Q���x).ҏ*��FLP�#�6^�i��1w���ܻ�@��1��ݫ�d����S����-�iK��4�^�OU���*l�w�=���/{��Cę
Ӓ���j���3��� j[�<Y��a��Y#u��뜅r@YHTz� Y{��G,�K^���J֨�-��ф�]	CHc�n?�۞(y�zt,�m�h�JYS�������.��H�5I��+}��_�x���f�cܲ\��W�/��W��QQ��V�3�7�2߯�,�uȏ�˙�"�}�ʥ�\�0�"?W�N%��*8�R���{��@�R'�����V1�<��mɸ@�.��h�K|��ǵF=kV�i}�y/�v�:s�N�b�oUMΩab��Ɇ�\�.Ӑ�=g�'#d�ܕ'��S�똊G)�(:�ne�]=���ȑc�n�{j�+�,��%�R���v.�o��C �qD-YJ@��u��I�Mq�y;;"UR�kQش�,X� ���^3X��}(l_���i
�����PY\�����N5�ԐJ����E��CX�u���r��zE��F���b4q�y�\��$�X�պ�śh���P}�'?����9���x�O�k���������/�*��&}]$Mo�DX�轕j�4ԥب���:l�K��]Ǐ�#~��|����	#�}��V+dn� �{%i�aZgb6W�4+���|��.1zq�rIP]+!NZ�ir-٫�h���l��R����Cd8}d�DՒ��?2�E�!��?k԰X���͠*B�.�����{� ���$$��������u&���z�ԉ�a�Ꮊ�i�A"mZ�^����J�-m"���Xيl�|R���C(��+3w�`8���J��-�
�uގ8��T �+�_�n�.1�~�h��3�T���+��}>]�qK�YJ�wb}$�2��Eʍ�%{���:tM��9u�WAz�GU�J�@I�,T��^A^�P]��-�J�L�+�QsRc�2fA��ɳ��9�|�f��s�dM�������HF)i�:mV�� S#�r���G�^.�dܩt$�FB� ���i$�Ž6�3B���Tz�_�Z�S�j��щ)򽤿���Q��T��<LZ< ���-%���0����Z�(be�q��i/�s9�(��Xʨ�u�S3 ���&cG%֪��}n��` �EP	2���%���Y�W<�3�g�Z=Wt[C9 �+P/1����m��w�=x�����ے�	=����<��|�կ��O!�ZF����u)�I|7K�G�SѲ!�x���N�y��jY�`��;R�7�]1M*�Uʁ5IPE(�N��2����^�o��H].��$F-/r�U�.B(e@��TTg�6f)z�@b+��`]�Q"���*.�����u�ЊF\�M���x�D�CF���R��PVm�l��*4G�{Ɏ�����<=�M�ǣ�@n��uL�f;��;J*X�nzq-���C�1�'j�E��w�v�����x��䚫�L��o�H�b����� w�+XU��ϟ�2{M�-F�FTմ=�����|+�^�q�&�g(Jb�t�Dʺ7�
�J.�rԎx��3�lu��5V�2���U�)�D�٢\,�}�'�,'h��C�3�!��3�f��B"���Rڎjx�n�l/�qWX�%Tu��ƽ6�[���ɂ\����i����F,��5�?d�
��~M��fz�,��(�;��K�,"2�����J���-���RA�����o �A��	��9潑-X�5�H�Ѧ������_&�Q�&���(�%"�=9v�NUVQ�ίT�؃�=���.(�AcI����N�µ�=S�ሢ�{I;r�4���+(6N�-syZ��j��cH�7��_�����6�W�=�p;�%�z���ϯ@����C�?�/���?��gC�|��ǆ�� 
����$@�����֮d�W6�>N4e���ׁQ��Xڧ��m�wy����$��..A;�j�f�`����ԗ�,�`��3D�����*����|
��$ӂ�_�7��SR����͚`WpP��Z��%V�3�CT�!m�-��@�XIR�t��И5k��HV�l�CqMN�IcW� ���hIqRQ]��%#�ѦCa��~p0��t(ܨ��%�d����IHl��Jb��t��Ԍs��E�2�{��PB�^�����\��Z�J�eܧ��L��]g�k
�7���0�F�������ⵃZ6����H#y-�$�8��Ϣ�d��K=4� Ւ�փ�e�t'7gn��� �0�9��K��5%&�Ui֒�~�	���19|ڗ������)ד�,�O��19�^u$����T����j�������^嘵v�:�6���E��	�=,���ZR�j�O�f�	�LT�C���Ʌ��a
o���> "��I�8�4KnJ�� ,��D@���|ǩ�3UO��q�G��fYy�dY����?��-���\���@5�6h��<�|%��cbŻ�F1m�7��vI|[��ڠ���ј��a���7ˇd �m�ۖ�Y|�y8^�w�}.����I�^jQ��HO���C�Ƣ>��?&�$ǉrE��=�荹���d��n7���D����`�.��h��t4�¶�*JҊ�b)�RwwaWq�	���I	'$��͏�Y��5g��T�����,�54H�Q{�S�N�U^_�c^�Ѭ�&�����3Z%<a��W2�tDx�;�噄N��TŁ��� C񺌖7e���V���	.�3��I�Ww�( D���d0Tx�U��� �*B��Ư��O-�0;|��]�d��m5%0�2w���q�P��!�g{���d�۾�mkC�w�ޞԘs�Lً�uk��F��6I;��Z���{b͉�����L9-e�"�n��HP�ӾZ���Ui��@�A�#���A88#V9�zck-�Ӊb�`��i�&͸&�ǀV�M���U�v6o�H줎X��������D�Ǜ��!-0/Tֽ��}���G	��-�m���j�35�$\RI�'
/� �6�l��x 7��v�B�9�aG���r�q�*J�8U�?a��3 xhL��@��A	m���P}`J�����X�)7�ph��qw�����XVc�>�J��_�\��e��be^�M޳h�ǦfoFl�ȑ�c���j��c��w(�^�f�����O}nWܶ�N�z����P���֟�ׯ���M�#A����EU7 Iz��%���Y�>ђ/�]i2�%�A� L0䱄l�v��k�6uф-b��64 ST�byۈ�8r��q&�;+Y�pbA�d.1�ʬi����c�f���$�O I���$�
����3H�-�zm������ɪR�z���3�*Q]��#��e�o��hw4�ɯDC.J"t"\��G��A��*����RAM%y�mwx.����h-�C��H�ڎ���p�~ 3_$�ɵ�h���j��!�۝�}��ys48�u�y�<>�|��3�D,,��NvKj9������
E�!�CY3]Iι�V=�<�i	�*REԵ�h�!Y�e-J���F��B�Z,`���A۱��B\f�myźi����Tޟ�J�z��2�%�H����� ���b�ɉ�3iX��QL�a3��\�O��'e��7({/G\^OϬY�Q=2Y�P����
!�\ͻ3�sȹ�p��DJ-�zɌ�G���˝�}j"e��j��=��{�ۭ��P2�%a���R=�$����/�+X"m�Ŵ[�I�9��b	�lR���;}w�+0z�FQV�h��M������cA����>�0>є$�Už����TR02W��p�H�5��|�z4W��r�B�.�D��oլ�/:$�\U˟�Cz�r��nw�քn���O3�߸�\���g��������!4?��Ie�S��#$Gc�<���9�b� �U�U�2m�-��!Z�n�ʈz���Y7����J2vp�;&Vݧ�c��ц"p��������~G�+'j�]1���A\���k�߭UI	�5Qc�Ԓ�s4��F-
���!n�v��V�����غbwk�b��+{���'P��.^��=�q],ީ�0��ȵ�+ֳ�ܐ�̍I�\7H�[��\Ԇ�h��.�0Z-Y�H.�Z=��s���`��jA�׀\�76'���X-8Y�d�w��U���%T��ג��sE@b����"-��Y�GgP9�a�e?�d�h@I���n�0�=6Z5�	�L<�5���ֹ���s�xr� ��:ƽ�
�j��O-�$|?���Ru2��C��FؤDp�ZK��
�J��l������ZA<<i}��׮f���^k8E�kU�wH��a�~�C�!/�hF�Bk�#�2ds��W�ְ�Gr����V��\�����Ӽ%S��D�y���I�,I���
g�:Vd���Ǧ��G�RP�]σAHq��O�q��'�-�V�m@{8�~$��C�A��-�r"p��̳0���kv�x�H~�"4��EA�KaHN��*S����*�n�TH>����LHk\=�&+��
���aYD�?�"?�'�j�0�2��]Q<���V��Gqm��\w(�i�������	<��!�	�#�@���g�����z���C�Z]���B��'��-����J&�����"n�G$��PmZ�.��`�m�\�<��S����jYVy.����r7�:���TTy;ZU\sJ�6j�H�s�� �vF�>)�UK�k �:r������l���H���G2'�Fk�}���9���X��Ζ��Zk�Ce�N�����oL�Wm���X;�B�AR�
��E��p������.��Ξ�g�(�q]47�b�~␥��NvN�oT���5s�k�ъ	h=-�^���.q$�6���E�B䤣�	$vj��F�v|�Z>xz]���^Q$��T�E��zy?z8��q�,��Q���e[�1����p�)F�R��Qq��~��ِ�k_�U>��t_�}�d������<��T�f���M���O
MF�A�"�E�t�%O��uK��-��r-�w^�>[�k�Q�q�k�G \��Xq���Zs��4����j��p�����S�9��%��W�R�{1w�ZH�hl'��&q7�hw�bFY�I��d��6n��^,4�Uh�u�%�tpB���Ǘý����!i�y;�%�����Xն/���|Ơ�"Q�[i����r>J��
�j[��Y�:��CDJ����l�C�|4����=U�%ᶳ|v��	W:i�f�QbŀY�0�H�玨S�Ԭ�gMA�Q�{Z%��C�a=b{!��G/ʤ�B��0sJ�kv:{���5؜��j���nu�9Y!RWr���]��l˟�o\���{o�'��?w
�B'<��O�+��[p��5��ۻ���_T!��!�3�.rS��I�[�Q�vu۳�*k��ˤ��n\M"�Q���z��c�C��E""-�,�m�V��e�ns���� h�%)U�M�� G��I��c��JL�W	�H��Įa�~Fb���fyJ�9r�#*�X2�7p� ��~�]���#�5J�.����]6�Y��D���c5�HDQ;�|wH�<�hN�(Ԯ�G���jl7��k��*�u�8���u8IC7p"`�y�(uӲʋ%~�~�3�U��9��<Z�QP���w&��A&�H�Y����Q��E4�A�Ȃ�e��(�"�����mW�t��G����l�Ӿ�4��%�dE�p^���t�0����7���AY}=�(�.D]�&�Fk0AVV��aZU0L	[���1�(�$��p�uv�C�l��5D�Vl״��PO��!-I��Z-�;�pDb�j�"*��rW���B�ˣ���2�Y��� ������#!$`�d&P�~5H.^'Zbʽ����Q�V����U]m�.Ħ���#�-���)��7��v��+۴��Ks_]�����JH��Lu�vx�jT�������TNH��j���zsX�sV���Ð�R�V��W�\.q?��=4�q1�:=�\�Kwy#����Q41q������ቅ�����9���k�.�-d��iv$��<��*fu�P�zr4���H٠�<��5^a�B%��h��F\*��(x�{�ʆ����Xvb��.�ZF)�g"���J�ь.{��g�Wb�V���Q��Q�X�bY�I|�+�BI|!^�f���,����1}�������ٳx�"t�C��,o�7��ē�_��O��V�O�e�yLÉė��Q��q��D+Oba|��Lgس�'km��PJ
��Z�Z-��>Z�&2o]�&��nQ�p�8$��e��]� vF+}�b��#�wx���-#J<�i��sſsc��<b�H� q/���%�Y����Z� '�v��AK����+�~R�e�[�����n�����W�p�����5\���/���2.�U$�׸G���]�X��B}[/:�h@7�Ӵn� R�p�\��U�w�C��v((��t�׳�;��.���>���������^v��� �n\l�M�����nׅaP7"+����!^c��~��u��w��Y��M����e�J��A'�U�S�H�BR[��s���a���FJ$h�C���z?Fϥ��xS��ɾ<���$Dݖ��&�
��޴=�yy�=�+.q��?A�B;$t��}�V�uw��D#��<`�/Ń�b�-l�lmqQ��X]8�;T���0��AJ���G]\v��h[�K$�x�kz��^�k��P�����2��w�ڽ�_߾�� �u�&$X�qs�r��'
���?h=�m���u^>�_H�[|�v���&S|��^��>8�͡AM�;�Dhq��M�Vx-*�^ց�N�~�q��H�UN;���5\�}� �����ݏ��}H�w�НG�=���p��Н41w�#��q)���%en�zt�ā�Ns��Z�T���z����:����{��w�No�c�Q�5I�,T�F	u}�D4�@�X�6�z���0� ��!�� �s������h�{R��n
�O妍O����js'��Z�|ܰ��(H���Ԩ��2��k�ѧ�iE��2G����-����x�?���7��y�ﵗ`��rG�9�#t-�~�wP��p�Ƶ�;8�s(L��������5�!"Yǎ����L�x&$Q_�@B9J�hr�es�I���d�����Zp��y�S3�\H���r\��[��	ʞl��O�to�X܊�FΐM%Q�c�<@�e�)���>�Qk���J�
��@?j�pnyG�#~7���Us�(��j9���oT�����[H�#���/���U<@["�����W]up�{�׿ԟ�A�Qfi�K�_3��?uir��iK�5�U�<X�Yۜl�dr+c��%���������ݠ �"4i�^���~l�K��\���~�#$�����n��l6��n 5���z�����1?�-���q�h":_��Q������M@	����|�1�
:����n��Dj���Mlɶ�f���py� .��.Ƹ���N��,[p���~�|�;�] �P����:U�m���&��v7(�#�B��琻���b�"j4����6������q�9Uזg�_Y\�pyu�~'��o�@}3ԋ�B�ڰ�ߣx�f�}Ŗy�4^�!���R1b;��_L�K�Hx�,]r'�����Ac�T�-c�Xi�m8����w�F�;��&�L�{AO.���UؑK`��:���Dq�ł׏�B��h�{Y����vp������\�w��߷�ۑQ�ˇ�Ck���=y��:�wᛞ�ϵ"�?���,��!Y���q�d̮ǟ��S�n��c����F���e`�@��<}���ND��a�{�q����[.��n��Jz���u��$<�Zb�[��l^'%s+k�����v������}WNy��W��/+�r;��V��Wi����Y�F��پ�󲺊���������=���O��w��HB'|�G���߅���~m;�����PX�d����Ń�ڡX޲�=R�&��(]��еW���K6�KLJL�=nM�y��ꂆPb�c��>b"l��*��)��ޟ:`��6�a���
�#�A@�l�d���[�*J)	�&�Y�4U�������A��H�0J�_��K�a�d~����g�:����VF��hӄ�JU-�@�~ַQqx5ٯ���Z���^����������HG���hli�~��m/]z��o�	��ٿ�����ݖ��+W�c?�ɗ�{�꿼z�$�a�D�ۊ\���=���:,ֹ:��!�� ���dǡ�Y�f��F	�A¡(o=�+5K�0>�+[��*�'��"IV��K0���4b�>����R��R�BIh�i�D�I��`$T�2��p�Bi�X��}�2O��b�\���d��B�H���ˉ�(u�'i$V4Gc�3�EB�#����;���v�:i�o��^Ajg�8�:���7^�]?��uj����Q
�uj���9o���~t,m9!Z�v/g넚�7p�#gҺ����vB�r��W�n���.�;6*���oO���z���owpR�~�a������Ο��G�k}/��9o���_Ev�P�n!+�t���aN�woK��q�\�DbC'������͐�7fb/�8
U2���w�d�G4j�G�J֕�E���Yy���%�4��/�p~���I�h��_F%j�ʰ�%)׭J'�`�K��?N>b2�ѧ�6��L�d��߬���@��+�t�R�g`s�;��	w,�z�3��W�
���`5|#�.~%\\���
��>4�^�?��8�Q����<�O$��Y�͙���'���2�lOg[Z��ru��%U����"�ٲҿ�	���F�����gPK�̽Ρ'���.o9�k�VC�5�T�E�	:��)�V�~�R# �Q(!d�u�H�+����� �����M�x}h���������U��.�on��-
��,W��/����?��
\{�X<|�¦�s�>?h�s�={_E�z����ۗ�f�u<g|�RF��e{��1��������֕����Cv�$��H!��Ą#I��=>A��k�xf�'j%�T�eXw`�&�Hڿ2T�I��Gz����m��%>ߴq�*�K��5͠�1��F-5�*�!*�\8�2��@zcw�M�7�|J�+�DCjC�6�ɐ6'h~o�t�z�h7�]}m�߻֋���$}���,shW�w#�k{p.��:}�����/����+��e��[�%��
�~x	"��;���������;o���Ґ�7��sz�܍js�2Z��'�6��u����G��?��~�nG�P����r��2��8ԱC��lJRd]��N|��4�r�* �I�t�����6��dH\���k��l*��ȵ�垄F�)_V��:���b����J+dU.UG�=��O���!X�t����K$��ߝ�KnO���m_&$�o���l뿎g�J�!Oȣ?�����;��	?��q�~#���W��r�8�%H7�L��O��~.��n�f-���dِ�HIEÄ�7�5�3��57�F$�U6�&Lc?'*�;&⹲֖�
%�!@Bo�^�c�t���I?�	l8Q�`����T�R���)n[hK�,R?�0�S��-�s�sp��\::8��^���ֿ�@|�^���f����=���܃�!/�5,P8����gΜ�����>��0�k�������j�.s~)��K���%�N�ڲW���TJ�n\`h�M*��U�'�Q�"HV6?��9.��a��!<�÷m��?��Ko|�k)�T���1�_�����.n��a�1<���~�$�\��uX,Z)���$���8�N|����u�Է�ݓ"JCZ:ɭ��J�c��IR@���Gi����q��km����3H�<�+E('�-e�e�����H>�(P^�^GfPJ���_+�#��i$Q�t�fGTy�8�8���"��b�:�T.7������t��>Ń~���쳴U�ͻ�����ڍ���t��:}	�"n�� id\�H��Y��u�41���btO">Y|����ӕ���!
��՗��jާZodͷ��fj�X7�ȷ${9�PʤB�2��ي:�5�*����w�"m{�!�Ԗ�X���$-O���s�5�Ggw���}$�g�����h��[��~��k/�CIM���
.�}8>Xܩ.@ǿ:�}���{~��Ǐ^����w��/��������'и�h���3�$�����Z-������D1$�b�b�Z?*\TRB@y,�X�r�k���ٚ���+�d��/�v)�L^+�8���<bd��h�`��`Wy��r��1h5J�<k�]F���,L|Z8�]z��?�FJ��f��|9�����Z��̣�l��yl\�;�"t�O=���<�?��|��+9�r����ٕ����>R��'q��萺�����4,�Щ�$��H	]\�b���&�b�2�hY�v�K�����3ژړ�T��5ר���j�r��~♭�ƭ�7{��ó8�x�")d������$C�tc�8��ษ��98���s~���K��w��/��ڷ��wp�O���1�;w��ӟ���������1ʧgК|��}����z���Ç�j�4��g}�m/V�_"�י�Y�Չf$SZ����X���)oП�2�M4`'�(\6f8LYf2����ÛF�s),E͠�w����DI��F9Zd����
���r���Bo�3וe���;d�kh��j����WQ���ܝ\�t�)��k�|
�Y:ᡇ�m,m��~�����{��p?�,����a{W�ǐ�?�W��H��"��C�z�O\DH�B�9Qt�i����Y�Kq2}|��5sR3�?��Y�U�mm=ZWK<;8�jNT�4�Hڌ�,t�~�עl�m7�*�s�,Z���耖,�1�%F��`}p��ѽ/�q���_;sp�6�o�&��;����p8���������y�m��}���s��j��'oý��O�����w�ǡ���L�|h�Ȣ��{�d-o�zhTlHy!֜u������B�y�|#�2�����[ו���9��N�0-����9j��t�Ci1�ڕc�A��$�)ɓ�Q�	ߏ2\���'U����_����0��LP����;ys�{N�zl~�l	�0uURS���z��2R�ej,������_�{C�°[��{���Cx���^܄тG�χ1!o���?�c������\*rB�9k���E)��[[�ɐ�=�h;�4��l����i_iz��[TR��N�� ����j��q��qLK�:����"�`��{��їV���}᥯\=\���K?��t�; ��'�����|�$��}�8��<t/T����rN'G9ԗ���c�2<����!�=(��#C@�-�|[�����]�=2��c	&��A�zγu��ReI��)�|�&"�[Ge��X�6�Mr�Ř 
06�	eh��:�UT��>�K&����->�?�5�
�ĺz�m|��R׿c�^W�Js��;��g�Mf�>�0�����Ԕ���K�C��}}��.�[H�oqV�嫰~���C�o��S���U��R�8��de�zu��zf��7�7�7��q�-mkf[���1�1p���)Y���#nY�֋o�bt}r'�m��]�!"�䦪B��h���n����i�r������4�����/_���g�y�_<��'O?���}�U���08�;��G��dI_y�۰���&��d�7��_|��?�{��Vi�[P#�&��������Q�܅�~�:,�a8LCZ#!���u��9СT�ID�Ȃ�
r�'9^8�$,iD�!C��F5�q%{��Y�Xq����ax�o��ȚjJ)��O��N��ŚH�*�N}
�B��F�����Fc�*�G�]l���K''�|��q_ ��ݯ�Ï���o��?�y�3��"�)��'���{��p8�=��V�M�"8f�m	��p8�9�	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8���o��<"�*}    IEND�B`�PK
     t$v[d��   �   /   images/d3b73945-fe79-451b-b309-b64aab767520.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     t$v[��9PN  PN  /   images/779eddd4-9cc6-4216-b155-89a4f50be07b.png�PNG

   IHDR  �  �   ����   	pHYs  �X  �X{�M   tEXtSoftware www.inkscape.org��<  M�IDATx���	�dw}��_��Φ��h$��.�B6a�x6/Jl�l�<�^�B�q|��>I�N��<'��/f�el���ZG�A#�H��=�=�{��FHH����u���Wսu������o�[�Z��j    s�%   �9'�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   ���Bqqy1~�7��b,*Fg1:��Z.P��`ԟ���6G1�F}ZU��h��q*�ϲ8�^
��Z��b�����b<^�����bl���U4���?-��qQ1�@�U�W\taԙ��ǣo��(�,]л敫��ؽ-���F�p���v-�z3���8u�^��ʝ:���h�m�tq��b�A���$$�I�x�,��|��.�ҀԳ���5?�����
��e�b����h���aC���=�.�z����4��{^����6�@q��b��"�w$!�I�x������b\�r�t.]=k.���E���ѱxE4�wFKGW�t�D45�WG��?��_�F���7�+��KQo�w=������&s�?�X���$�Ͷ?�X��o�Q\��_�ś�����c�T�����S1xt��{wL�6�:����Ew1�U�b;����E��0�:s�xA|Cq�_��]et/����n�%�o(}U@�*7 I����e��q�с��h:/��uY>FI�¥u��2Џ<~o~��8��!?����,�׋��'������sD�3'�������/��K�zm�~�ۊ8}4��  �Dy$������|%v��q��oF�:~f��p��۩����Q�z_�,�̺�E�W��ߊ�g^?=��9V��ָ�m?=�7  �Bs[G�z�['F������-����Q;�Hy���b���E�<`	tfM�"�V\������_q�b�{?���  ̖��FW�⿍K��x�ӿ��wgn*w$}��~�����E����ά(^���-/O���̼����ҟ�����  ̕r���_��8��]��+N�}�ro��b[�5E�o�1�N�/h7_-�s(_�ڷ���ˉ�� @ˮ�5n��x���]��3���b���E��PC��*^��/s�_�h.�� ����ƚ���y�����hk�DKS%�|����x�U� 4��$�W�ܯ��W\[��oN�T.N���b��]E�>�F:5S���Xq��j9�ֻ8���'b�E�O��-�h��;b�X��K�Z���w�S[cE�������G�����@�(��޳�x�?~0�O+g�;�>[n���5 Щ�����s��8/�������^�aJ?ga�W��)F�D��lk.���v��ŝ��폝� h7^7}����<���Un�~��ֽ���o�g��x�*�C�����W����OEǒ��3V��ŭ���+�Á�dP~�❗/��}sW��;� E�����~2��_��G����=���H�p	tΫⅪ<��k�(�R-Z{����s������K��U+�9�,ho��˺��� 4�r�Sy4�=����H�����ɏ�)�}W�>p�tη/cey���=����=�7��?�fUO��K������keO�@�Գfc\���{��1>:\�Z^����@缩T*?[\�ؙ�K���Xt�g�w��o۴t�s搝���q-������Ŗ?��3��^l��Z��π�@�s^/L��~�������������C������-`>x��I� ��]������<{������Ŷ�g�H�u/̘@�|��bL�o_�l�#�fA{K�����μ���p<y�T  ���?G�/�����6�/��̐@g��3X��.���GKgϤ����)~�q��q��h��#�� @kWolzϯ�ÿ�/����b��_U���3 �9�[|��Ηl�>V��Ó.�\��O]�"�u��8���ظ���&N���C'�v��Q'i N[��Ʈ��0�'=No���?0��T*늋Ww"6��#��y�+Ǻ��Ӻ���'1�~�T<�7�N��Ș0 `�ۼ��������3sn-���T����$Й����/��X�~�oZ�7�]0�;�؃y�10<  0�^ty,���q��o��g���9`�:�V�T����Lo|��O�|�uj?�邘|���=�o ���#� �t6����z释m��j�jÕi���/����`å�����t�[7,��������ϔ����}�  ��`Zp�8���r���?L�@g&~�̕5���I,����u�~h��X5������  �կyۙ@/}0:�$Й�J��Y\\<q��9V���I�/㼵��n/�����9  �êW�5�~�w�:6qd��b[��Z�L�@g�~:�|�ڦ�m���]��Z��������9O�  �틖��W�*�<q9Yn#���#`�:���3W�\z�nZ��-M��C��{v  �O�m��z��!Й��t]w����0�W��9�8^��Ҷ�  ����O~�w�LN�^�@g���knk���xم��{.Z�qN?��q��H@����O�eԛ����H*����z,��[#iz���okԛ�8�m���*'�L�@g�*��%���1�]+�G���F+{������v;�&�F��ãIODC���Xk���E��G�u�8��ZZ�k���߽}b��f^_�VwL�@g:^�J����.�fA�9������l�P  �|Un7�Ko(�'�@�3ן��u�@_��zN?�#�� ��ֽj��'�5	t�D�3K�\i_�t��bI����� 0�}߶�)�Lǂ3WZ:�&]����>~���  ��;��?� `�:�����5�%�ۚ�-�G���;  4���y�0E���<s��m�Pkm���)�  �����ON�'^�@gf*���  ���/3$�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�$s���طo_ԛ���h$���u�K�� � �������V���  �J�  @   �   ��@H���������z��֭���[�(�������@ԣ?���ŷ�7 ��K�$���]=�Qo::;��4����z,�� p�y�  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @ �{��F<�ukԛ���h$�=�P��G~5��������ܹ3����� �t�dN��M淓�����`�l�?.0w:   $ �Xz���C���hM�mQ�z/��P������ҟ�c�{>����+ �{ �JsK�v/�JS��X'��:& �&�   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@�����  @���T��X\p��Y���r   �L�SSO>��O�̮��  �F&Щ�{w�������旼}����G  ��	tjjpt<���}�VĒ�>܆Ǫ��O��  ��	tj���H|��q���X��#Z�*q``8��'�|�  �$Й��Չ /   /&�   �   	t   H@�  @   �   ��@gF=��<�/`�V���h��	N+�G��S��^�!�l�>����c���/G#Yq���wQԛ#O��vD�Xv�-ѱdep����{�_LU��'fB�3#;��t�t\p��yNo�}�7�Q���'�2��i��XZ�Ჺ�=w����b4��>�	��<�Ǐ4�s�A�  @��x������W�aV�ҷ;*��;v,������T*�~_�Gw��b��=��.޼)�����.� ��o�F�v�����[��s��c�Ν�(�-[���Qo��������K�.�j��.\3��y࡯�����S$Й�g��;c�5o��;m�uT4E�yQ����?�ѶǶ�s�a��y��'�m���֮���Xz橧*З,Y���Qo����9(�8�r������Kc|�������,�ـ)�   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   ��t,�cO=8�wZ9�3*ǏF�|�t�Z����͘��m��7���x2{w�Fr���\���wk$'N����Ѩ7CCC�ٍ���Q�_�ZulgT�g7{�m�²�)�Lǥ#�N��_�d0��@�/��?���o?81�߶?�ub0��ٳ'h\'O���۷�Y��;�4`�:   $ Й��7�)����������ϣ�?�s�(\tYԣ��Kj=��߹-��h�]��{���Q��\��8ypW��o�K�3#k^�㱬؈f�{Նx�~)��:/����n�4���E��L����.Й�   	t   H@�  @   �   ��@  �:��R�K.���:������c���14:   tf��xϕ�cuo���������ç  2�VǣR�f�Tf�@��Z�+�׬��]�/����)�{Պ����Ğ�  s�:6cÃ�^jjj�����ӛjM�SSׯ�}�8?�����%�o�  �K���"�Oq^}n���XT�NEKGw@�	tjj�Ү�.s��h+J}x�  0W�GG^�g��^�Y�47Ԓ@��z���"V~����%��	  �3՗?�q�ZztjK�SSM�xR��   �@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �NM�����  �f*��n�5�NM�>>�z�&]�oh,��  �R�����ȋ��^in�5�NMݳ�x�juo4O��o<��  �������}a�7����Pk��:00w<q(~l��hz�Hx�@����  ���:����щ�J���"Щ�o���[7,���:��R���q���Pq���  dR��v�@gV��E���  ��&�   �   	t   H@�  @   �   ��@gFN<�5��=���E��&��:��F����OD�h_�<z�l�z3zj ��z$�WFKgwԛ��O�б��z��7GkϢറ��8�����6��PV�ȶ�|<`:n�wwD׊�ӎ=�h<���F��֟�+~�ףޜܿ3��w���5���X�Შ7;��S��/F���C��eW��6t�@�=��:   $ Й�}�mW/���ٽׁ�Q9u,M�:u��J����b>z�[ߎ#��[�n]\r馨7}G��C�=�b��q�UWF=z��G����(-Z���Qo��������.�j碈�e�z�G����ľ�)�LǶ���^��w��6�?*�F��Ͼ(������>��S���K��"����fۖ�*�7\|�}�������4T��X�"z{{��<��3�tvv���������_{�������@�0E   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ Й����h�<���iS�᨜<�fdd�E�vn*棓����x_߼]ǓٿgO4�����\���wk$CCC����ftt48���1�_�\�؆����r[��0E��vx�Xl��f���x��G~5�_��������塇'�ߎ;�����[�l	�r���\��S$�   �Ό,�tm�/\0U��]���/Z+o|S4�]���{AC��R�;ף�1�r�qk._����=�ў˜C}����oL�@gF6���c�U�03.��|���[ײ��c����4��EK=����=�̀@  �:   $ �   �   	t   H@�  @�Y��T�=m�\�����qjd<   8M�Ss�b�nâx����ib^����/m;'G�  ��	tj��-��Wv�`^�W��U����=���t  r�Vcld8���6k�_Kk4f�@��6-�zQ�?�]-�ƍ�㎭�  �T�C'�8?��<�3�Ǌ�hn��5�NM]����\��'�rۑ�V  �����sq���#�������Z���Ү���\�����  �+/�߻mL�Ss��*��~>� ���hOjO�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@���ƫ�u9  ���Z����S#���u�e�Ǫqbh,  `.U��"�^��Z���C{�c�ҮI�y��@�U�A `n5�����hT���7��t�C�	tj��''����/y��������  s�R��������Ĭ2��p�� Щ�r���;GN�ƫ�-�֦�s�:wl=�o  �"қ�ڋ+��M�Ss��j������buo{4�~``���  �G�3kʓ��86   ��@  �:   $ �   �   	t   H@�  @�y��Oǁ�.`�^���K���w=;��S�X��kb�k4���ά��� ��?���`Uԛ�w�Ƕ=�b�m���?���'�j�Ⱦ��������0��v��<��7�g���h��Ѻ��Gj=�ֽ�'�2Џ>q���(�_�z��<����� �   ��t<�ڵ������Y����mQ9�L4���ѣG���T*�˿�/c>��������`r���x�[��f��g�}�S�(6]qy��;���K��|l}��h�֭���Ψ7�cǎ����5k��WuхQ]��Y�ϝ�'1r�)�L�Ѧ���]�iVﴩz"*㍷!������2�/��ʘ��\� 8�%,���x2--����`�º\�������H������7�8?7�k��_�Zu�����b[�p4`�kk	   ��   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ Й��F�bϽw��VN�8�������j5>�G�Ѿ�{��{r��y��'s�Pc=�ݱ�.�c���������/�������c׮]�<v�TT��ջ,��L�@g:֍���~9�}e����,�_;�?51�����]<Ww�ߑ#G��544����r�=6w�.`�:   $ Й�W���;^ty�T�/^|Ϣ�W����G�h_T��k���Z���w�G�|{���-�(��|O��h�eΏ���m��x�t	tf���Mq��703�=�<��@Kg��X'z�l�4���e�e|l4`&:   $ �   �   	t   H@�  @   �̊�=m���câ�h�Tb��pܿ�D<v`    �̂+Wt��/[V����ml눍�;�[{;��?�  ��ccQ��T���R\4��NM]����8�kW�Ğ�Cq��  smlx(�G����T����c"ԡ�<ʨ���-x�8?��:  s�:6��8��W��>-�{ԡ�:5�vA�Y�Y���m�10<  0WƋ@)e���5��Ԓ@��:Z���:�r �9U���HΚD�	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   ���x�zN˝�b   uK�SS�㱴k�e�6�  �S����i���|��Զ�'c���I�y��P��  ̥���~��JSST����QFMݻ�x\��7�t��Cm�q��#  s�����j������hj����.
����jy,�n}�m�����ų}C  �{�[:[�:^zš��.�N�95�w�ؼ�k�p��J%������ԈC� ȧܛ�M�3+ʳ�o9001   x1�   	t   H@�  @   �   ��@  �:3��kG�x `�6���h�]�6�w���Q,��Xy�mQo��g��t4�o{ot,^�f�}w��D�X���U�ӆO�����:ypW�Ltfd߽0k���y�7����ߣQ���'�2Ї�5�z,����C=v���h�7_'Пg���{.9t   H@�3��v�^�����;���㻣�:t(������T*��g1}�s_�g��L�W]������ݵ;�����ho����Q�������Ol�F�z�����z���/�����X�jU0U�����}���1r���S$Й��M��h�5�z�Mm�Qi>�����E�~�k^���_��@?+�����'�mKcm�,����\���yOl�����;1�͉'��kmm�ŋ�Wu��_;�ۭ{�#�ԉ�S$�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:�3�j5~�#��с�������oē[�F�<5�d�C������  ��O��<S���O��D_��`~��  �J�  @���w'@���a��{fv��.�[�� ���2.���bD�`S6��8N��q�H�v%���)lCGb�@��K"�#�����$J��ؕ����j�����h�
��ٳ���|���׽Ө������   ��ņ�LMME��
Nl```�u�5�v;&'��8�f��֭�^� �!�!�3�<sn��۷�A�V�k۶mq���G�9t�P<؃'�;�-[��K_���E?�p��� ��:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@g)�kMMĞ����OZ|<�����kjj*����x�޽;zM���=�:����~222ccc�k�e�]��Y��C���;���Y�+�,�@g)^2;5O|� V�����`m�#v׮]�ڷw�ޠMNN�,�y��w��x�,�@  �:�r����}Y�b��-x���9z�/���Ϻ0z������X���{�9W_[.�����-?F�7��>ˬ��];�/�y�R	t��W�6N/X��mg�y?����6�y�ױGl��ʹAX��g�%�{��:�"�   �   	t   H@�  @   �   ��@gU4�*.9}C\�u�������g�hL̴   ��*ض~0��3⌍����K��'���  Ȥ�nGT�U#`�t�j�Y�;/;�D���Ն�w~�����'c���  ���Ӛ���Tt:����h4��nX��*:]����q~D��x�E���J� ��To5���8f^�݊N�70�1��:]�7N�0�c�ߺ.����n9 ���=;���p���WM�Dwy��U����*c�P3F&:  'Q����.�U@w	t��>c�BT�v  @��   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ ������>  ���Ntg@�	t�j�3Sq��>���l�M�  N�Fs ڳ3�7�*�^���]FWݺ����<��_{�`  ��V�o�H�~n^�����<[�aet�j��L|��3�8�#��'G���  d�Z7���Ӟ���:ګ��:]��=c�wl&��`K\�u��z{Ʀ���ާ�  2��͹�M��*v�NǍ��   ^�@  �:   $ �   �   	t   H@�  @�e�w��brdw�b���������g՟�����/6�ual����5ӇĞ;����+~"�6o�^3���1�������1���Y����m�X��v,�@gY��,ũ���@?ʡ���~/�Ź?��{2�'�?�W�cm˅���@��7Ů��T�+~�z�~��gF��� �   ��R<2�n��x��W�I���G5�T�v�۷/&''�۴iSl��{[$���b�޽�/֯_��zj��������D��O?=֭[����1::����p�v�i����xFt��xU��o�٩�GI��;���Ǚ��Ī>ic��Q=�֮C�	�ذaC�uV��jZ�����:�����*зm��7o�^3==-���r�W?���sƥ�>wu����_Ձ�3`�:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @���|z�@<��?^�g�/c"X������������h��v������q�}�E/���c�=�F#z���t0�zyܫ�徱�������S������$�Y�M��l����ʛ����m�V+��ǃ�orr2�_>˽�~����'��H   �,�e��Q���	X���T>�i�s���������E�Ͽ��^������,_��ߊ���oF��<g����g�����[����T�ei�?�O	`y���R��c�h��SU�,�4M_v�L   �   ��@  �:   $ �   �   	t   H@�  ��Dkf::�ٹ�e��  P+q>;9^n�ߛ՚�*�ގ��p@�	t  ��=;}L�?7fn+z�ht�@  (�-�ǿ�%��:�  0�N@�	tV��u�hVU<3Պv�B  ��Ϊ���7ŏ^�5���-79ێ;��[y:fZB  @��u?�����o9f��@#�:���`�p��'E:  ��:]ua	�����^|�P��K��v<   �L��UW�x󼏹����Ň���  �L��Ugn��1��yh ���  �~%���F���5�8  �^%�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@��Z�΂7���  �*�NW����7��1ӭN�N�  ��	t��ݣq��N��o��V�t  ��	t�ꁽ�qϞ�xՙ_�������CO  @��t�'��#�3q��[b�Y�ͫ���_������L;   ��@���׿�ȁ��c���CѬ��[�}l�q�   GtVM}����  ��'�   �   	t   H@�  @   �   ��@  �:   $ �Y��#��  ������j�ޞ�<�ǉ�E�,�葉�ɱ  �^Љ�zU��Ǭ
X$��R<sd�59  ���}��u��$�Y�}G&�  X�:�v��lAo4��3�Ǭ�X$��R�ydb|�c  k]�={���vo_�.�c��Y7�#`�:K��#cO>  ��ufO��~�����E�,Z��y���z��jl������o  �N��v��W������z��3?�H����yQ}��C����^  ��w��96���~���X��R�ǡ�����v� ��T��=;s���fT��'���7�����,�@g�n���7�7�#  `�iOO���j`pA�g�����
X��R}���˨��{k��&��n}  �Zў�:��U#�z���綠��j��K �Y�N�3ZUU}�[���[✫~:  `-�f�5ϱ�����=��h=�%����<����Oe�~=���o�  �	sq>Ϯ��������7n>��,�@g9�W�{�h������p��  Y�g�K�O�������~�ؓ�Ν4��z��D�%�t:SUU}�L��>��ß����_��  �l�u^¼ݚ���͡uQ5�?s{������>�/�:�����,��+c{��_�).z�?����  �B�3�ռ��Z��y�hDc`aǞO�2���s�{�2~5`:�RrUUU_����X���@�௼'  �)!�i�涖��	�Z}�ys���׾s�8�귕������+e|+涢&�}�[�E_  }��R[�`����a�>z��������U��Ǐ<xG<����s{�²t�����]UU}��k���������Ϩ��^ @�(�@�S��|��wk��r��8�Zq���;���ɲN|_�2)(V�ϕ�����];bǧ?���  ���)q�F5��1�nQ�f�'��C�}�ȏ���~!`tVD�����7����̇c�˯�S_�# ��:838��gioG�l.�����7���p��_+��+@��bʂ�%��L��>����v\�/�G��  ���j4��<S��&Gv�=e��c�?_ց?�B:+�2�(�����?���߹!7n	 �^U�{���ټI��%���\��G���;��k1}��#�F�xK�
謨N�3SUՏ�ɻ�}���������i4�wl �ZQo��/��8�\��ث���I��+��Zӓq����C;�sdV�m�k˺�t�
謸����Dz�%��e4��~W������_�w1�~c  ��z����G]fma��f�<�E|n�xy-�ף��l)�z�����������̪_�k�:��+L��e�����*����j������ջ��w �m==  zN}l��`�;��;�w]<��Gf�߼�rY���] �隲��X��e�eT�vm��~�����q��  du�{���{?2��r��e�#]"�骲 ���;��g�jg���w����?�~��  �������}o�g�w�y����u�Ot�@��ʂ�s%ү.�����^�����0��w[\���O;;  �d������{���ѳ����N{{@�	tVEY�}�D�9e�+e�P=�o����mq�[�~\x�/.�Z�  �\황x��|$���њ�:��:��8?�
:��,؞)7��P��r���hԗ�����$�{������wŹ�{�˱ �*�uѝ_�x<������OsWP�_�E�*謺�����(��*��z�����cn�p���o�s�~sl8�  ��6�����o����gF�w���g�:뮀U&�9)��>q�%��Vn����ѧ���`���b��^g��Mq�+^�^|Q  ��t:1��C���[c�7�v��B�z����z�N��IU�7��K���ܾ�����57jC[N�m/�"6�wql<���p�1��3c`x}4� ��ǒ�NN��9���/����ȃw�m:�G��aN�����%��]���k�X��z�Z�Y�竚�� ��5;9�Vk��,�Ke�nY�# 	�N*eyg�y[	�F���2~���mg�Q��)♱g  ��S��2��}���(��d:)^`�txD	�M��2�f��qq[ʨ�o:<Xa�ׯh6�U�����v���aÆ�F��&�;���3A�6m�5�^��˝ �zyS/wbh�Z���	��><��(cGߊg������h@rkbA��_8<X%7�t�窪��X^��7�y{���7�\�/�5��o|��Hyﬕ/�*����~-�k@Y�����^{M � �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @8���������5������l6�j4�ưh������n�g�4&&&>�S��{gvvv2 ���p\ozӛF���k���e��d�"���oo��`��   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	���y����     IEND�B`�PK
     t$v[w�'<�  �  /   images/44e1934a-57d6-434e-9b76-9cc9cf9f98cc.png�PNG

   IHDR   d   �   �=��   	pHYs  �X  �X{�M   tEXtSoftware www.inkscape.org��<  qIDATx��]Y��y�o-]��>�F�iFh$�c��b6��I생�NL�<$���������)ǎ��Ā}&66X�� ��@B�f$�m$�>�ޫ���oUWwuW�t��D��4����֭��˿�V D�2$`0�	B�!C��!CȐ�!dH�2$`04�IQ���6xt���[XO���(Ļ@V"���M�ƎCtI������ĺ��sӾ,Afjߊ�o��T�N�B˲��q�*�C�Cz�4D�{\e�����̉C�<uġM3h�!��N��NÇ�y��W�n�cۥHTk����
��J�H��0d��Ma�����V,��?"�i5
�^�=3����,�Ű�Rw�T�Z.��b+�(@>9)�_V^�/�?��gsȌ�=���/�ա�_4�z��P_��������ۍ��F"����L҆���i�h��-�FZ�o ��x'P�$Cvz&���~��\OOvÒ�; ��S�.+p���@�[��-��g�о~,����G�d27 =v.?��?}��m��x��z��;>_�t�go��W����>�<N��	�􁪤NL���	J��� S��dc �����w׋��,�@R5,��eM\�YF�"-X�id���"#����qǵ��3c����0�z�h��H�����޲���}��>�� j�B8��w`�g����o�'�.�O�M��Dv�#G"��dAF3�+�wt��&0q��3g�s%�ш��K�82�)�q���͜FF��%�!�� �;e����A�w g�m����W�����u_<����z:c*8;c5$57E�ZƵ0��o@*
Y07�Bÿ�8Ά���@$�=�M ��gY��Az�%�AQ粉����R���ڣ!�p	�sn��� �W+`��.����N]��"���4Lku�Ym��n~ߛMK�C��u��a�2$`0�!$��N�Yi�5�{-��zD�t��d��t�l�A`B$WTZ{�[��R ���U�C[W���؛�� !�G`b�V݁~�KZ��R�h�x�ճ����څ���Gv��^�g�%�+���u�8��\���"0��m���0K��S�T޺f��c���O�BE��0����gN��H,a��� �-���\�f��_�S1�b�,K0>6�����-����������4Xt�!`�v<�^�4,]Z��1��v��Ld���u�p�&���AKVC��e��yX���Ca���2-`�Z�R|t���0�i�����"0M��&��x7eTl��6��]���4MLc��EDp�5�h�8܇i���3��CB,�!,�rʻ�3�IP�LԪ%\�Y-���k�	�ū�e�*�$V�|^tݺ�.��+˚5-��5��'I�f�C���/M�^�=�Qt��(Ɯ�7W�N!�j�ǝ����L�$��[Amiw�!Bf&/Z-s����,b������W���
���La��w4r��ҝdi3Q�O�fH�c9d�����Q}��灡8*�~ �t�,iҒ�½����Z%o~^N���ȕ�HR�p� |�uԘ� "C���0~ݶ�U
r�L����`U�x�h�p��(���x��R�����~��_���Z�+���[&w$����;�䇯�������͌1Ϧ�/��f�M�.ĺVp�c���*0z�2�P|��J�~�jg9S����!��G7Gh&E	֭-тĴC� �g�A�s�@���׻6nX�2���x�cId�ϸʐ��\�٢Z+�>1|��"��j*�]}�!����M+_�͐�D�O,L ��`>�a\��ộ5C��h�';K�ax/�d�B�Q��]R�V뭊}*����:����k�*g�̙��_�%+��EQ'��[���dD�I�D���f!I�2AKV���E�UŞQ�hz�O�-cc*Ix�8V��t�s/�>��-�'�#a	��fջU�m��У�ڄZ��!���a�3R7\	;#1���Vp-Y^G��wo���kK`��l�V-R�s�����	P���p��G!�2.���(0|j�r��L�ŠcS �U��t�b��V��vO��
-b��f
��AZ����#�w*����d�.�2�V���!���X���[T���5GÑB�ygIoD̔* ��n��L�ꖺR��\jGۻ`���`�b��Q�ǫ��=�|̝T�M��f�ø����_�$�an���mt�� 1�V��T��Z�l�_O��d�f�\Y\� �}^�0�Xk��w��*��Z�.���m�AY��5!�>�-]i�	�s�X�#�`F!�я2姼߶��ㄯ. �aab�f�=ˆ�d�,�,�3Ė8h$������-��ͧPU��IE�`B����]5m�f��k�l[*n�'�x7��PS!i2��(�_M�Y�k�(yҗ��c�̟L_����S�
�
�	Z�m[�"�%_�*��*�(u�5�ɜE���^��/@'�6�&���,�͹�i����l�;�&�y��i�m�Zkg)�
�4��Cv�U�Si1p3o�~,�zKu~2��O���Iѷ���M�>w
�N��iz0�i叾�юe�!񮕆�X*�$��-�����sҸeM�;��e:y��!�{j�1��M��]�@K��i�x��s^2��!2�����u��N3��ax�im]�IB�U�g ::Tfˢ���[����̈�5`�½#�f�va��]B4�6���6�EH��tJCs��u�,�g���xy+p]�e�]�/2a��C�U� ��W2�@�9-?DX����^�T��g�u<�nZ4`�g��4��{CޚC��]dZ�0�	S#��d�C�����A�\���VQ�fI*�o�!���e����~�X&C���J3�ܾ��d�旟�f�Đ}Hʤ�e��:Z�E"�Ȭ��QA$��2ʄ�Tʓ�tMG���G�);P�z^��Dd�o���a��E�C�5��`t�-��4pϐK� v�>��;�*��F��: �� [g)0I3ǥ�hSN+?�͐����X\Q�6l��;���q���+m�$������b}���k�������Է�`��Ѧ���f8r�2y�wp'�Q��r�"a�w���\����X�*�^�X��zj�ۭ\t��HȐ�#�]%�V�д����w�rz
�&���Q�#H�+|G������t��i�C�5q�u�Ϥ�+ܽ��AH�����̆���ll��*V;ٙ1��~��b_�E��A$ϳ'}<����$����"��*���b:v3*�À���nF�Q'�y]L�&�)�_�)�T�6X�%K��6��V�d���R<*4R��=�t
S��5L줃4�d�(̵x�/��߉h������?�xZ�ӳ�z�
C��-	�Ae9���Z ���j��f�?�Ԉ����i]�-K F����泐=�����vH��\�y�i����G!7~���{��{<~��($'k��ޕ�D�g������u�Cj�m���>{Ί:�9�̴��$?��^A��w�0$Wl@��d`�Cp�*��b��t��=f�Z�tB�6�����lX;�:96|
�H�Ab銒/g�����,F��si�w�$���W2D��_?ꅣ���&h�:�\�0�0]��L�V����c����Cb8x��!Qں���lYZl��1T0��(���Qʠ@�rP������vh��vٲ�Ӟ����-�Vi��K9�(We~�"1$&��c�9g��E󛺓����+�m/�S�g�a�%�u�ruD��t�)Sb5�/&V9��װ�~h�E%�`��rP���^ʟ��D�3��F�a@ F�Aǲ	_��Sn9�����4���(LN�����sC�)mզw�҅yƴu�3+��c�
i��+3��]�]C������#�f4�-�-���o�d�/�ge��e�,U��!���2d	��ֹL�뤞 M���ߌ�?}�4H�T��dR�x�����	���'�.�=�3�6@]_<���7@6����dJ��Ժl�F ���f�����d��"�6d.�Q'6�|�7C:c
־n�t���9��Ql����a���94��z�FW��-��[�Fd\b�YB3Imis�}�4+�g*��H�_z�] ���oPLi�e!{o�����]�H|����%x�M+_�8k��&`z.s�����8�za1"�W�%�[������l!�s�)[#�����9�!ʠ"w���H���];�y���d-G��v�dg�����Q1�%�Ƞ+Z�	`�M�߭��.��{���&�#t=a����i��FY����l�|jֵQ�*tUYN���̤h�L�f�hk�ۯNm�z�WfCQ���dJ!=+,�˲8H�$�8�	��$���E�9w�x�ψZ�,�N�2���=���-�Љ4���[$��_���v��N�!<� ߶۝A55
�o?��KDȑh�s��\X}'ĺʎ��0�}�����SK� %v~��|�#�J������ʠ�Z����?;=&�NlZ���o���V��Xw��u�i�udI*�B�T�(r�n�ru�t��/���d�\D˒���oCU��OA�"��fƚ�^ؼi�˖���Rp`���8��#`��*Q�D�n���`G=�nv����A%�lZ�, ��>]��Tvn�)�t�]�Q���� ��JG`��f���"�%�����d�"�*r�8贬�{�9��n�Gϙ��x��������C��x�Π�����5�ѝ
���{����ǛD�U�a�͊��Ǒ��������t�5�Ɂ��.�Ó��P�/?��s2;�|�y�����-X`��'V�H�b���J#��4��5�I��e����f���=
J�#�L+-�8$���2Xs ����xv���bf�|#�9{�
��T�tR<+=yN�q9���t���Ͳ�\��`U&��z�D@�S��*�b#���eȑ�Bl�e3��3�E�Jۖ��A���D�&_	S�a̳�30Hsz�x.���i��3�.��.$V�����N!��ͻ4(i��XHYLK�M7A��+S�uY=IOL��oVx*-�]$��� Rݞ[?ƍ���9����53���|ٺ��H��;z`��Ae���6�(�vxh�F�w|�Oe?j��bȅ�HӪg��b���H��j�J1�N�(?˱n�6�X@��-��jis�x�L'�T�i ��__|�b|���0�XZ����*ӿtUĂ�,��T���M'��R0�5@&MVb��^?������F��ϊ���u�{,�z�W�,����M�#�����!���I),���C(�T���KCo�O}gN,[rr�rP��y"��l��3T�k!S����`m�6Ȝ]�����[���O]��?�6H�X�ŔUX~�#�=�<�j�g!{�u�v�m�ݲ�v��|S�O������SfP���n�u�:Bh�6����u.�YdH��߈h�B�G_�(���9�ҙl
��^A��3��:��o�P�C�d�,o�6D��A���%}!mҽO�t��%����!r��;(��|�:ln��V��p�-��Y�>�@��w��}�`ц�ڴ?h>�JDZ�0�Q��|�:u^N��qv��A�c;�\��-,+�-a�0��L����m�F]���\���H�-�����w�t2_8�{��[��ʒ����av4��d���'V�tU��e�]^�}��4:�DkE�s�g��!:��Xi1i_ ��|Kn�F-s71%��c�Yc��缃�>e@$�e�����hl�̤Q�}$"�*�a�$ ��@��Ȓ%E�$z����}Z�����s�G2!�Dz�����[R�|�2�ڗz��D���C*�(�����A�\����[w}^0�\�jE��=w��[n���\m��vb��T�?x?�d��/gP�a5n9�fG�*�V��S�M��ٺ�vA:���6<I���#��P�S����\��m�Z���z>B�ʠ2���оvKu۵���]�� �AE�s����'��.MgP�Ƚw]�tbNNe��������H���*N������?��*|VD��o<Z<,L�c��?�὆�!CȐ�aA�����F���|,��l�y��h�!8;�3�&Q	�k��k��ڔǐs�����!i�g��"��Iτ�&�$IM�Ԅ?Ą���7`z����^���Z����:��h�z`� RI�:��G����+�9��_�?ߊ-]�}ō��v�U�G�Agh���+1r:>Yr��zdѕY1��~=��+Fa|�z��2˜CGG����r�g'����>y�W?�~�4Ő�����?�����po���7Kj$RKs���eu�G��%��N�c0�ɝ���KVr������Zұv݊%�Ov0�9pb�{�\!M��^�������5},�,&/>?������$�zon��|����[cڠ��`"�~����We����]-?s��o&������x|i̞;~�C�A���V�ز����ܰW�$�צ�Dܹ<�VF�Q7�s�
ovn�ʑi�t�ev������G�y�޲�s����_y�ɩԙY�dU���`W�C����o�H�?y"��+��K,�K\ө�WEט����~q6�7����^�i��CG�W��35��,h�I+��܋O�O-<���0�;�W�..�=��GW��g�Ϻ��30�5+�o�O�H�>�.�ڽ{w�zT*f�uk_���=��ݻWD���r�L��ܫBn}�Q�E�4�ˮ�Խ/-�����|}��]��$`0�	B�!C��!CȐ�!dH�2$`0�	B�!C��!CȐ�!dH�2$`0�	B�!C��!CȐ��J2��Y���2X�N�i$ܟ�e�U�}�bt����ʃ��_�h��֛���P��lo$ܞʼ��n ���]�P�(���v߯.;C
�D�Q
��1�X�=�'�kZ]��D���<Ӯ7�����y��8ܟ����+ey��D�_Q�ʗ0��^(��=��:���j8_�\�=~Ԏ�7M�����egH����Y��{�[L�RV�2$`0�	B�!C��!CȐ�!dH�2$`0��48�_4O    IEND�B`�PK
     t$v[wJ���  ��  /   images/f9728bc6-2422-4ead-9082-90351081a874.png�PNG

   IHDR  �  �   )��   	pHYs     ��  �8IDATx���	��e}�����sN�{���  �NpILbL&���'&HLn�F�u��%��Y43sI�b���q>���I"��+��4�4��Yj뽧P�j �s����?�.h�p��_=���   8�:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @: <�6��䪹��|X�&�L.,�t~'M���L���t2�ٙ4�	�l6M�����l(uBZ�>���f��?�[NL�~2���o'� �d��L�L;�]I�<�o��;����W5 �: <��û�;>-d�K;�lX�f:K�>f'�t8��p;mW&2�b�s(>�F���7|⍍�dj���̤���X����ه�$ݒ��9�z�}���[ ��@``�n�f8��8��ɞ��U�L�|�W�E�К?j#�2O�7x��I�B.������?|V(=�p2�9����O\2��d���Ω�8�J��d�w>o�����F  9��@����[.��j�ON�:�d�x��Ei��B��4�	��!�6�������k�ۍ������U�|'w&��]��Z|u�We�� `�t ���^qB�&���3[��QI6YR�4���1�b��<�ւv.,h�p��z�D�ُg�o�إ�Z��s��ұ��^��� `�t zڍ7�X�w��gwBxq���ʵ�ݛ;$���I'�)7C�P
ݏ�������o�̵��϶r_�w�m�λm���I  
�@O��o(ݿ{�w�'���;�w�|b:ӫ�I�ۅ�Px|��5�ڹ��'��\��F�������� Ϟ@ z�7zd:+���֋�Ӹ��d�S
r�l����Cn�^5��?ټ��$��N���w���� �� Dg�������$���������ڒ4�D03������6NitW���u��Kv����3�]5��nZ< <=�@6|r�±�ɋ���/?�}��N�Ƕ����~|�\�!�^����_\�y�w
��?e�e�n����  ���!s����/,��]H~��c�v*Β��N�S�����\��͗|���ڕ��ض�n��� A�0�F7]3��=����B��zh����N>�7�W��>f��K6��F����P�|���� (���ۼys��/�v��^=��rb'c���N�^��
�l�����+���r�k6�S �#��6����c�C�?���g^���&�i=��X??��o�؟�e�U�����߾��Wo 0 : Uw����W^��4.j���f6�3�ʶ�J�ՙ��W���5�*��[FVW>zU�N �>%�8(ֿ���uJ�?�T�3��ζg8���5
�S���'�oY����'7��o_���  }F��ߴ�7ZC�׍g��2�]�L�v�=��]U_�}�%���Ul�޵񢍟	 �': �Xw��/^�(7���luE��]U���¦7}������{g����m��	t ؆��0���n��U�B{~�C��k�l�64>��㵷���\k�/�ܽ� �$���4�w�G&�ӵ�w��;i;@dZ��⩏���^�=�Z�_���� �C: O�M����K6^�]��V rIhM�گ��/[��u�+����Ƌ7> �t ��+n�bE����z���f������d:�j���L!�+k>��S�f�τ: ���y�Mo=�Z�_1V�xY7p��4����K����~h��.7����{��  � �7�����{J�^��N)@��d;��R��R㗧B�$�����k�=  "`��n�f�]�q���دw�9��J�T]�[���������y׬^�:	 �0��}`��kC[״Bkn��d���r�����k�?��~o�� b`��}��_h����Dn� ��m-m�n]{�G.}�Hk�������z �CD��� �ɡ�_W���i�	������5��O�ټ����ٗ]��v �a�����7�����?�3�o���� <�4tr�B�ōv붵������v>��$����M���=����j��I2��r�u�%�������k��� ���n]�*&�O�'�Oӎ���,�r�Ò��Mk>������o����  �H����t��Jc��
h;;<7��f���Ks�>���ѿ��5? `�t�>q�M��i_?��<9 U�K�Vgծ��Cks�МK�`:t��!ݐ�����R�u�L��i�=.R+�/h�[�^w�e�_w�;�> �A$�zؕ�\y�O���z�~x fD;�OO��K?��?d�7\���� pt����+�x_q|m'�)xf��䖍,���M���$I��^p j�ک��ֿ��e�o��h�� �#��c6|r�½��7���� h&��I�O,OUyw�:٘���KvW��w�v'����b��O&	��H�/�l^����|�-��b�; Ϛ@�!k�7�k;�=�*��8H�Z:٬v��C�����FrݏsV�?��4;;'w�wN�l?2�h�ښ�~�{6�Z��x�Q�n[��+׹7�gK���7�wƯ���/O�Խ�t����U�U�'��B��]>kY��q����ڵ��M>�~trg��nX^��ʶ%Cc7]�������Y��\� ���� �]�=��Yh��˘鲧���j�����|%7��v?��ҽ��ɶ��[�Ƕ�j��@Gi'���P�5�G����׵�����o	 p�:@�W[?���`��n?˿43�2/��8y�I����㱾ml[s�16��^�7��-�r��+.�x�;�g � �"t�7�=瞿�(���-�̄��x��4:�\)�\�>ݳ��/:��Q��%�Ƿ7ܷu W֓L{dbx�������^���^ �g� ����+V|����7�ͣmig&��m/��􀶹���ٹ��ʉ�N(��j?��ֶ��[�=0_ٝ�f'K�՗|d�1Ci���^}��  OA�Dd���_2>T���m�0�v�v'S�~������-,t?N^zr���#���jv����m�|�$���o��[��o~�o� �It�H��������7v�L8vM>�s�,��g�׷u?&ɖ}[�y���Iߗz+�Z����[���u]��  ?ŋ@�Clt�5�����&�p��M�N�油�{0Rɝ�䔡���nݿ���]�5����N�S������?c��YW���'��������G�����KӴ���V���ys�|��yG���wD�{V�{��4����������b�U����Kn��w߽��c �@8d.��������i��ݓ{���'��Y����任�o{�oC�Ql�\8,�?/���W���Wo <�p�}��M���I%@DvW�����S��;{���'4&��v��xp��fw��ߴr�����y�6�f� M�̰�}C�R��08b4�Ix|1;��9���{N���=o��J��y_�}6;i�I;�̝�ݼ~��7_{�� X^̠K?��/'˓�H�~Z������ɜ�^#T�ܩ�N:nѱ�{����T�������Y���nY�꺋�{W ` E��/@�ڰyCqof콵|�� ��]�]�?��/?m�ǔ����C���B�HC'79�X��C돾���] 8Q���O��|�=�������s�G�;�"6\ɝu�Y�G�;���G�]�S����Ӵ��,U_�f�9sk���`�t�i��}k�Ndkk�G��"w ��_|����w<����j����#�G6l���V_� �0MF7�.�7?�ʶV�!�V-�6��Pq(z@�z�峖��ZZ����7���z����R�P?3�3��oX��W�4 }O�L����^jn���%zЮ�dUqUO�2!�9f�1���,/|�o�v����J��k��W��'G7]�/�|2 ��:�A����=�6���8_�G��i����zP%?�;oŹ#�M>ֺ��ժ�ɞ����5�O+�ӛ���W���޾; з:�A4z�[N���}0�&s�����=���xxq��������߷���^�?��o1>>1�i�U/��X �/	t��d��ѳ'��ޗd�� =n�1�i&�N1Wʆ���2'.>��b���W������g+��k�J+῿�����m�}�� @�� ��^q�D���~���7Y:kiO�f�f�^|�G�C���w꽺���7����e�/{�;W�� @_� ���������ć�L{v�>����=��'�"��������}=Y�\kI5>���7���?�jO �ot�����\U�5y�T��	��/e�F�{������.�ν���ܳ�������H���r�^߸k�ޏ�n��妻���,u�9�W7�2�a �2ݳ�'���T鎭_�|t�Ѿ�7�{j{�����sܡ�d2��	�N�,^R���/Wk�Z�Mzo�Gg+���k.��[.�E����,l�䆅;�{���m-`٬�Ӗ�\)�+��G>{��C����� �@��,��m/Z�7����������#_�~Wm���V�1�|��y������~��W5 =M�<CWn�r���ޏ����U
����N�,Y��V���8w�S��6��{o0l�䞤����-f�_y�Ж�4���7j�6@�^h>o{��7o��իW��'�O� ��E�\4<��}��o���9+
�N�y7Ɵ�ǇK#�s���s[??ًgx90�M�l���������3G�;�4�27�Ň�\��&{jwH-_;�s�;�a��k =K���잏�=_?:��r��9}٩CKG~���EË
'/~~��~��K��;����=~��U�UsV��ù�������-�w�v�?�S[ޫ�ڋ�~h�;���k� �$�p��x�o��Y������S��2���x���G����=��k��P�g罍�ǂ���Q�(6{y�;h-���W�3���{w�SOC����뿵��o��w��! �s:�X���WL�����T�dNYzJy*�K��?m�����d����k�k�ڻ��j��r��y����O�[�OXt|yNyv��۾Zk��1k!M;����KG7�n�x��� �)�g�tӺWV+�ׇ>�`hA��gU�C�z�r&d2�<k�S[>3�kgwyv�z�]Q���5V�YQ<n����\��g��ZV9�E�;�~a�W��Ӑ�&�k�\z����z�Ư z�@xk޿�����������p���OXt|)�`�\){��s�?}��'�4��F������=�|p��fw��q�+�)����K�r?ԋF���ze�H'�)��4�a�=����� ���`��ˎ��j��	�g��;f�|)s�ag-^|P�ϚS��;g��C_x苓�tn����{�������[˧B��E'�G�hE��+f/<���Z�W�-�Bknfn���M׼l�ŗO �'��D����l��V�5;������sV�=T�W�%���ZZxޢ畿��;&��n�o�
���B}圕���P������=�q���*�B%{O�|}7s�U��[7o��ݑ?��S~p����r���=����KO*wCc:�����x�m���������[�omn��<j�Q�_�=��b����H�s�]�4��H��8��7N=\ ��@�){?8vu}����G��(������9+gd�~7b�\~�P�Y��S�c�n�uϨo�}�m�j=�I�UsV҃0��P[5wU��+f���+�I'�c���W��z�W7���� �� ?f�ͣ����W����R��9w������s~6�͜����O����z��G�Fy6��z�+ۿZ}`��ӗ�V�����/<��o�c��n��5�	��H���n����w �$�~�[�8a�<yU��=�����y�sW�3\Η�=�����[q���~n�V�~�������S��/<�|��cK�L����[����/�}��&b#��픪���]���_�z��� �� SF7]3<Q���TB�8l�a����!�y�y�3��6���_�?���"�}���Y+Ϊ���l�� /<��<p�dw�@�X+�Z\��M=�� @tz�D���Uy��i(�1�-���r���9+�������ƚ�ɧ�m���Ǖ����{x�t.�^|�F��E&�QGz5W=cݭ����W_���t`����N�'�} 3�7�.=�r�#������O*�7&:;�w��Ώt��߳����ɝ��54T�ٳ�B%��#~n�3�v�ښ�;���׮ߴ���^|�? �!Ё�����~y�R�����\8{�YC�g-+�u'w�}ؙC�=p��X}�������=ɿm���ӗ�Q9l��(��D���y���|~b�9m�wB���4�j�=�wm�Í � Ё���}k�6g�ߞ�NϮ�=!��g�[u�Т�E���=��:o�S[n��~�53��i�_������j�����^ ����#.��qowO2���{6�^zU�h?O�A"Ё�5����i�=��/e.Xy�pw[���sV�=��?7���?����4�+��8w��m<��D��߶��Q���ǎ}h�O�:���x1p���e�Mj�׽>텇_8<�cwJ/ZX螕�{�ݵ Ob_m_w����+�^0��'_�tߌz�����y���w�L�뿷�W�۵�{�g �TO���\����t\��=������_0ܫC����ƛcIw�4���F�g�����N����*����{�������N��v����4W/W��t͋7^|�d ����@ټys������N�Y=l�0�}�?7\��������\�Ot�|��It�L���w��7�;�,9��Fru�31�<7���n�I'�/�V���Pz���� 8d:0P>���_7+ͣC�A�_8��>z\���sV�5tۣۖ�x͡����5�I�s��Ӈz���6�sV�5������ja�G?|����� ��@������j��[��=�G\82�=98������+�����&�S�<��������y+���z�ґ��ӗ�V���✽�	��B���z�[?��׾m{ `�	t` \t�EÍ��5�|�Z)_�\�����j�t��t�Yy����1i�;O�{�{.����z��s/M4':��u_#D�{��Xe���z���'Ё�0墫k�ڂУJ�R慇_8�k�ڟ��Ë�_|R��~��i��I>������p��+�\�w��'�������F�qr����.��� 3J�}o���p�4��У
�B��V���H���]pLic,�ne�4ƚ��g��ąG��H�Ezw�ݙ���lU'���&!B�����6_�?޹��� f�@�Zwj�m���ޫ[۳�\8oչCsʳ{�����rƲӆ&�������1��t#�S�^�H�es�V�7|ۖ�LT[��Hlg��Fho�z���#Ё�����*�V����v����-,���d3�!`��嶉Z�]���#��;&_p�=w&��������?3��b���.��k/��#�!Ё�5z�[N���[z�)�N�,���P��p9*\>=��It�B\���%���~�H�Mw�]��;�3*_���j�L�v2���[F7]��/�|2 0�:з����������_:jޑ�0�����<��ʗ�}���������C_��n���=��ˋ�,8&����E7ٽ�i�/�v�c�� �N�}i�-�]6��86���+��脲$�A��/:>���{��ӽ��·爵uؙC�y��<�I�}��ɮ��v�L�X{���������� L+���+n�b�����4�2/w��3z..��	��W�����m&��3m��P�R��O\|b%��L�d�^q�Ч���x�U����NH����_m޼��W�6�`	t���˭�w��r�1�|��Q��΁�Yq��Ӈ�ݳ�~�{w}�1Rɮ������t��9�����D�F�衕k-�����S�	 L���5�_s~=_� ��\�{��������E�͋��b�]��\��];�V�������=�Z�{kA��J���b��Vn�����o�x�c�i�3�h�d8�ew;f�1�/?�2(w�?[�B���?�����1]"�I���m_���#_<����N4&:������X�={���/i�Q�����P�X�˩�� L���X����1�������9+�:�gj^e^��e�}e�W�����4����/:�#�C4�=iZmLv�N�������2�w�W���������q�\sg ��@_X�y]��o��5@*���́�}3c�T��x%��Wۗ|�o�NYr��t�\�N;o�'�~�c?|�]��i��:��1��? :��N��v�=/��r��9w��C��́g��%�/OL��#��������[�����+�8h;U����7�'�kcI����}I�5�	���=���_}�k��5 pP	t�獾g���r�7B���p�ag�r�������Y+����OOL��@D��]�]�_��*=�Yi�]�O}��v���K����}Xa��ݰy�ǮZ}U3 p�t��5g%oOB���S:~�����Z!�Ϟ���������a�[��N�闷���#_0�T�V���tj�ǚWL=�� �A#Ё�v�M�g6��sC�
��	���7b5R�-Y��՝���'�g�wS�����t�W꯾r��z��� �@z�p��{�Z�b��9{ř�aUΝ?Gͤѹg׽�G'��{w�SߺoksP΋O�vH���[��9 pPt�g��u���)������J9_�7b�I;�=[�켧��m=�I�4��^n�����5o���� <g�Y�|��ǧ���UsV��^��gi�?t���m�o<��z�]X�$ө����*�e��L�=i��ֿd�P?�Wf�U
��)�Nq�������}��w�ƚ�Cd�����n}�Ƌ7> xN:Г�#ɕi�����"�Y��Y�N<#�N���G�U��M��!N��)%��?O=\ xN:�s��t�/W�c{�׎Zpdq��BW�=C�M>ֺ��j�V�vv�\�T���7�u���yێ ��&Ё��n���yw ܉�N�X#it���7j��ok�'$�S
�ڟM=|c �Y�@OY�����G�q���*�l�'�L��T�7��qw�tv�=�R�������x�;� ����V��3�3��,,Yjk��^���ǾS�����I��Z��;�}m �Y�@��y���������K�ok���%_���ɱƘ���㪅�/_r�%�߽��c�gL�=#�t��ʽ�'-9�\̕Lm��[ڻ���4���@'����d��� Ϙ@z��{F��U�	=`nen��yGO)�$�;���Yn�j���W�^�:	 <#�	�Y��NH���.�����yR�)�_����=�=^�Cje��P��k�� xF���=��,6)���*.Z��)��o~��z��9��F��� ��1/"�����C5��k�L.s���O��GZ_�����������lZ�+���� 8`�چtCv�'��F��/<�T�W�{��}��_��A�à�T�?��N�<���&/n��ȕ���1�.~B&���~�����o`�4�׿o����k�	 �D�Ul�v�'->������I�]�]���P'�ٴ�y��õ�"Ёh]v�eG�&���]��[5wU!��������0����Kn�����_�zW* �D�]��Iw&D�E't�Y=��4��W���@hg�Y��|o��� ~&�Di��͹�
��B�����ܲYK�F��@7ο��+��c��9�V��=�$��@�tG���*���u�UK��?!��C_���!΁i�'u�,����~ �i	t J�r�������Ë�=?��~��w��9�ӺG�Z��uS� <-�Dg��F���UO
�{���\��C�������O�Yh�tC��-We�� ��@�Ӟ�yC����V��/v�|ʃ�lܳ��F x
�\2w��c�q��� OI��i[�"w��畜=����]��g)��:���@Tֿo�KƳ��!b�K���f--������������A�7�F�q�%7\2��k�= xR�JRIW��������^o�;_����N���	i!������} �I	t *�|���R��Y9g�@On��F�n�xFڥ��)	t ����_ޟ�77D��yG�2��@��}�7j�����j�'�yߚ�7��� ��@��ʶ~+D,�͇#�^l��m�-{��NxV���gr�ߝz�_ ��@��!ݐ}�㻣�޾r��b1W�����4VK�|�.ہ�$��J� OJ�Q�����s۳CĎ�����'�v��m_�L�Ĺs�9i�'n�䆅W���]�� Ё(�C�+C��V�����s�7�Vm�9�	 �Q����D�N�w ~����������'v�"vԼ�v�|Wug���8w4�b���.�~�@���>����H�3�̊��2�۝v���w��`g;p�r��F7]3����' ?"ЁC.
/[5wU!����j_{���Z�fk;pPu����/�zxk �G:pȵs�����r W���u��V ��B��A���R��FO�+B�F����+�r��������wW�4iۧ ~�@���e'���-�j���T�����켧�h��}	`�2�W�r��W_t�7 ���!��/[9gE!���D�e��� 0͚��+��� ?$ЁC�׫�>)DjAea~�8���G�^�I �n�Br~ �G:p��zϾ&��^��b�a�z�����c����h��]t�E÷\~��� �@�¬ܯ6C�2Sߖ�Z:P��I;�7�f= ̐NH�.�^��� �@�V�}f������r����p���7��Iw�3���� �'ЁCb���G�
�:l����{����|�`8`�%�4�Y$ 3M���xc��B��峗�������h��Uf\#�\�:��P I.����9�J�20�����!��Nnɲ�/�z�?����!�)$��H-Y:Pύ߳zbI��� �:ph�r��C���,�v���f��A'�� �����-'�e�Fy�y![�t'�����9�f�q�tC���Un� �@f^���!RKf-�gB&@��{{�X=�$ө�_����w�&Ё�Φg�H-^<0ϋ��h�[5��@���{�@�����.���Z4�p`��칿 "�ʶ� n`^�q��u�ζ�����Pqh ΟO6&���]� �$� �@f��ϝ�l��ґ%�e���4��ģ�K���7�����1��50/F�H�g�H-Z0ωݫ���`+ D$�ܖ�[��F� �@����C�-�����n��"= D&��wϡt``	t`F%���!B�|)3\�B�n����s Ji�sb `�Q�\�<Dh~e~~*�����f����ɠ8`�	t`�\z㕫ja�P�Ђ����޾}lG+Ma� Ћ��N�o���̘����Z�Ӽ�y���o���V����4�x�� H�3��&��e���)���@���]�v2i&=o��'� ����d�cB�*��l!���n����v�t��f�@�@fL'�Y"4�<��Wϻ{��v z�LzD P�1��Z"4o ��w�N�����v ~��$ (�̈u��U&Bm8DhNyv�����v���@��l{a P��f��P���٥�}�|��nu�$�� J�3��vN�fra�8������N��$tJ�Z�@fD'�)u��G���$�v���/	 =�����������ȥ+B�f��{{w8\'��@��:�N}w[ 0�I6]"4R��@�5���v��t�� 0�:0#�\�(DhV��}om��s����a` 	t`F��N�Sy+�J���Ƙ@zJ'$K� ���ۼys�_��
i��P��'��۵N�݈��<�SK��� 0�:0�>߸{qZH������V.��:���VρޓC` 	t`��ZQ�+ʙ�Է�����t��tBR	 H��/Ӊ2Ї���|��s�%�SZ�y]����� ����2QNp/��}���VЁޔ�z�z�-`�t`�����r����ۧ���N �A�y��$w��L�N��*�}��v=�Ёޔ43�Z�@�_.�"T��z�{�ݰz��l.�  �L�N'�@/�J}��^k����4Ӊr~	�t���K�aV�P1��g�k�t�g����(��$Ё闦��B��߁ު	t�we��Ё�#Ёi�	i!D(���{�����L1 �L�L�*�|�ࠩ�������O� OB��.M3Q>���
z�Ӷ���N6�����E3�g�i��5�l����@�f�8Q�h�M�[�s�l��%椓��?��2^���0����=3�-�~�ǒT����A�@�]'Ms��p&��.I��g �̀N�+衯Wϻ��c�Yi&�u*0p<�Ӯ��l���|*��zWR�S����vS-��m)7���=������ui?Q<	�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �  O��h��2��s�dB'_�7 }O� <�N'�U�M.:��C����Z8�� @��  O�X)T�vy_c�>7 �4�  O�2����$�V�5+ �4�  ?�М���B�J� ��@ �2�����9�k|I'� L� p 2�Lgd�T��_��i. �A&� P6�m�~lb���p��_��t�>��!Ӫ�*�\��ods�d�~�����]���5 ��@�S�f�8�ora��� },_*Lv�C�ɟ��k L�Ї�Fyb�Ĝ`.}._��F��:?��� 8�:@I�N�^�5�-��{�B�><d��\���$��D�jjSq` L�y�{�Y���C�y�~��I���� �F�Vi�g��\�5<o*γ�N���� 8X:@K��|��������L&��̟��LMl?P�_�`� =�QkTZ��-��n�/y4��F�O认O}��� <[�{w%�]������^�{k�eyw�Ƅ�!�d�K�$d杼�eN�!!���cb�:���[��p��c��wf�aBl�}1�ٖ�Œ,����.�����[����ߪ�]tI��������F�@]�ͨy� �BIdF���닅t���\uq X ��jg��Ec���xq�K{m���s�I�5�@  ��@�0���Z#F�s6�0^8�e��X�l�hF��� �t �ǧa��F�l�!2q^��N�~�  V � ���4��H�D&����j�թ�� �B���8>�.[��g
��X�6_�Z3[  +�@ �p|�]��l)[K5ʍq�� �F��%8>I�R���܂X�Qi��� �t � ǧ�EIƫ�
sb�f�Yj�Z� @�� �G����fa�8+�j7څ�bsB  �" ������l���y�8Y�QJ�X��������  �e: �ǧ?�zn�8Q�6��V��/Ԉs @O� �C���r�_0q�H,��Lm��J��
 � z��ӀQJ���Ҍ�P,��tu�8 �� ]��i�s(�
��c��b�0��\m�h��, ��t �"�O�#���D�r}�PDn�Du�֚�  =G�@�4�<�?FƋǽ���H;չ���g��  }� t��� K�8/Oe��X��f�<Լ� �  t]n$7�ʦb!s�au�:!�8 ��@  ]�-f�3�LU,d�f���+ �w:  �L1��-e+b��|u*h9 �:  �T.��+e�b��B}2hy �:  Xq�l�Z+̉���x��.
  !� ���2^�0^8!�j,6G[�ֈ  `  �7�6��Y�T��,���1 �B:  Xq������D��ڍv��؜  ,E� �eS��Ek��o���B}J  ��  �E9*(M��?Gb!�dk�i �r:  �`J��8Y<�*� S���8W ��t  pa�D��빁X(��Tu��J�8 @�  �B��xq�K{m�P�^�Du5q H  �/]/�2^K,�ڭ�q��v �!� �yɏfS�TC,�#�,����?s� H^�  �9ˍ�N�s��X�糋�u�S @�  ��d���L!Si-�:W���(-  $�  �*�r�����L���8�0+  $�  ^P:�^̍��R���d�r @��  ���L���ω�j���� �@� ����^�0^8!�jTc~�/	  �@  ���Va�x\)�b��bs�Uk�
  �@  ?�q�vq�8ck�7��R��  �  ��\�'K3�Q�X�Uk���	 ` �  �C)��s�U�X�o��F�1)  (  �u.Qa�x���@,䷂lm�6-�g
 ��"� vq�'�Ǽ�닅�v���W�s ��#� n�8^���^[,�W���-�  0�t  ��.��{�%
�ȭ�V�h�] `�  ��H�D*�j���P�չ���9 `��  �l);�)djb!i�6W]�C�  �� �����bvQ,���j�a� �!C� 0D2�L%Wʖ�B&�ks���3 �"� �l���͋�j�թ�� �!E� 0��W/�N��j�ɠ� �!F� 0�ܔ�,�g�R�rc�o�E `��  �8�[��ҌR��B�Jc�Uo�   � T�봋Ek�Ym�Z�֨  � ��tF����0/4�  �E� 0`�Raq�x�qU(j7�|�Ҙ  �ct  ���ǹ빁X�o��B�8 �4t  �N�'� �Q�J)qG�R��}�׵�A+��檫ļ�   ��@ `0hIɂ��_�M�+�v׉\��&�ͷ�c�w'�v����  � ��R�,�j���E��9<Ɂ8�{�8��}^����x�Ы��V�~��  ?B� �t�T�8o��C������n'��h�繑	y7�|�ǋB�VOTWk�]  /�@  ����S�^}�8ޝ�ֹ�;K�nb=����#�,����?s� �9� �����y],�l����H����Z�xge<  8':  I�J=���Hk��q ��!� HG�*�,����G�8O  8/:  I�HK���XJ��Q�$#  ��  $��v�b�8�G�8�
  � :  I��Wieo��Q)��  �F� `;%��q�u�r� ��  ,� ��B��\QN)
  X6  Kiё�qM�Gb�Pg�8  �"t  ,�cf�\��b�Pg�v4��  �2t  ,�l�;*�0J�&� Xa:  vѝ��勍"���|LQ�  �8  �������b�H{Q;"� �  [xb�)6���q>�D9  ��@ ��S�⩆XH�8Q�8 ��t  �͕Z�u�Q�����b~�  ��t  �ɑ�J9U���J�zL4�  �/�  �#M�v*b)�[{�)  =A� �J�q���R��8O  � �Ӣ}'�,���8�H2  z�@ ���q�ϋRZl��8γ  z�@ �wB'��k3�n!�GE	%'  �/t  z@��ܬ;�y$6
t!��  ��!� �2�N��8�A��@�  ��@ ��t�Lk%��(��8�G  �� @��8Wi� �
�F��D�hT)%  ��t  ��1眻�-�a�_�s  ,B� �*�L���F�N�S�9  V!� Xi�,�q�Eڋ�q ��t  V��TU<Uiq�8W�  �!� X)���8�������s  lF� ����R�b#�U���b�B   �"��K�`h8Ҋ�"6��\�8׼� `;^���0T:�؄k(i��� �2���q�$VFN��빑  � +Ik	�� X�;��*�,����yZ�h:~^�.���L:�峁  � +Č�~�D�9J�8��E)+W3�q>*�d��j{a��|�g4 � + ���g�|��Nƙ׶n5��8γ����2��l&��2����!�`9��v�w#�z�a�EGN�5qn��������V��u�B�wŞ� 0 t �@Li>:fF�E�	l�8��Ϭ 
A8��j�Ly�R��o �� �)����8w��ӊu��8/
�JiU�֙� �@��`vS���>�tg�vG�b�Pg%���2S�͌�|1ϔw H0 �Sڇ�J����-6
uF�zT0��0�Ly���� 	E��9�@�A�
��'�8�[b�H��v4���$3�����g�t&m�^	 �3#��,̨y�z���ʢ��(�^Ԋ�u��hԛ)s$[�K�!��L8Bm�)OU�Su��7j�xa�V�s�� 9t 8֛7e��S5�P��錜�bV���u��B�u" ,G��s�8o�>�͇�#�8��B�8oFb&��s[�Dz����r: �"���'·�#-�v�b#�U��cB��h��y�I�<�ڬ�x�m���Ͻ�o : <������v�b�8ε�s-)��lgFԳ�����E:rˡ��{nx�3rϧ � � 2q��
���1U���b��-�_;�"Z9��С�ƿ�Q|k
�IV��lyZkI��:%����[���}�>�G�n�S��:mqTg}�2�ۥ+79��{�7;�{r�%.��û���+�|�\�����'��ͷ߲��v~� � #�/�1j �W��/ҪPʷ�r�l;�T��ݷ��靯�i��? \(�P�Q��s �.�Z���#�#����>�G��^* 0�t Cǌ���q '�JOJ��fg/��w�������� �`�t�ZOy�&zC8 XI��t��w�W~�����O���g �`h,Ź��\���S-E�Y�������Փ�}�z�������� � !���q^K�!���LL���֏���}�q�k���I6�0Ht Ϝ�{r�8��Y�t�ww���G���o�w� :��W�6��S  ����ި5R���~<3��n���y�=$ 0 t �\`�M �s�(�s���SȵҲO?uۍ��ow�s�n��#�,�L �i�ڞ�0.��X�a:t���#�;* �p:���l�<� ���ly��t:��R�\�������>��s� @�� N��v��  VD��L9�������e���o�o|z��F  ���0P� t̅�  V�9�0Rl����BZ�z�?t��_��?s���"���Y�:q ]W�j���k��Y�n�V��y�K�3���"�3�c"]  ]��2GW�|F�L��տw���O���_ $�` ��9� ��]i6�ugw��k����]����ol	 $� �ر z������v��Ǿ���� 	B�H��vl��3r��ٺi܌7{�o{�/|�}��� @BpQ ��z�F���p �'fyQq�`�zt�z�q��6. �:��2�l
 �c��0�ŹB��r���z��?�W�_ H @"��-�lT$ ��2{�x)/J�SV�GZ���p��o���?- `9@�Ahvfj; X��hzf=��8N,�Cw�q����� �#�$��Z�:q 1ˍ�պ���Od�.���7������E �� �Yo�� ,d֣�z>�vD�陿��N	 X�@�fj;���̱�f-��G�-f�o��[?�{>$ `)@b0� �g��kJ��������Z:�D0�&�� �3S�ۭ��Τ��ս�mg^��������s�% `!����v3mR  �Ь7=/��rW���c�v��o�����i�Zy �����  #�re��Jy릺�Y?����U|��	 X��^ V3�$�tI $JN����"�̌���ۿ|�o1��6: k�5�Lm��j���h�%�ig|o�?�O��_ �� �ǹ��p �\�9���ʱ+ `���02u<G@�ٺa�E��?|�g��>� Kp��J�g�� 0ƙQ�|ֺ��ǂ��W��@`�u̦Bfs! 3#�Lsw]ǪQ�F��{�mox�g��� X�@`�f��� `дM/_��b������O: +p�*f��c� `��~��A��kձk����������/
 ���*����2;�缜U����)<��] �ϸ`F�`��۾��f�֢�y�o����w�Q �#�5=���n��\!g�Z�������_�w] ���`F�`8�Q�L.�v.��,�� @�� ��j�y>�!avt�m��k�x������ ��b }����s 6��k%2���� ��@�wfW_ ����t&�E�vr�W:���/�t 2�f˳-ЃL���m�s�g��ُ
 ������y��� �ab����^ʳ�\�rP}K��@�:��j�=�a�}׶@��� }B��09Z �������}�{��������� @�� ����  ~��d��֢�Go�?� z�@�7� �ہk[�W��Z�> ������  f�SF�uk�������7��?��� �!@_���  9����2��B����;�{:��"���� K̬*�e�&e�x� @�� z��� �S�i��u����^���?}�����y�!����3z �q���=Q����}� @�� z.�Y �q6��^���	 �����N�Lo <��段��y��Im� @� z*ds8 ��A�x)/K4�Vn׮]�o��% �:��
X 8���@מV�?�÷�w� �@O�)� �i�x�Z#���� z�@�3f�"�� gb�qkuin �@��^�9 �E�k��x�zS%�!���� gc�:� �n����w�Q �2@ϰ� p6f9�XD�?�J����& �e:��0g۲� p6Qd�r�z��%!�� ��'�0�jD `'�f�mo��u�2� ��� �Ud�kF��q� ��DFV]l �eۛ�-��
 � ��'l�� `/�,J�=�z!�� z�' =�5#� �scf]y�+��<���'o��c���# ]D�艈� ��䛺��Qo�_"�t��뢈�s ��뼩kW�K$�K ��@�u�� �W��z�hF�u ]F��:�: �<���ю�	�.#�t#� ���D ��@�u�e�� �gۛ��9�.#�t�� Ηm#�
� ]F�  �:ZGb�8�S ]F��>-�� Ώe�Zi^� t���"˦) p��� ��@  �ul[��:�^ �t�f�8 @�� z�@   �®�| ��@�.q'�t���*���s�����$�!d�wa@� za(/j���������J;AWān��P���5@��(�Ȳ�2 `;M>:��ӌ;  �� ����:#�*  Αm'�(e�O��"�t���6 ���w C�@�}\d ���7w`�� �����U �|Xw� � ���P;�  p�th�1k�A�:�����uy� ��0�
t ���t]E� �KV:#� z�@�u�� �܅aH::���) �Or:��C��:� ·#�Q%�� t]0M p�t��ۻ�t �@��	D)�9�  p���2:�^ ��DFi�@ ����F0�x��A���O9 ��k��V�`0z�W�z�0��8г�  �&���@�+:���}��� g����5 Ê@����#툣" �B?L�et �B���Q��M �� �sw- �u:��	�~�M� �3k7�\�Z<���+�)d �3i5[V]�2�@/Y�`��]nIk_�0Q �<�f���%�@�K:��1]Q����  ���jg�2��!$ z�@�S~��dt �i�-��� �Gt =�j�ҬC ��Y
%!�����ڭ�#�C <����m��L:��28�fݴ�  ��n���^u��sF������f��.� �g5ꍴX�(�k:��k���h�i� ��(ӁXU��9�~ ���� �j7�9���t }�4w ���s�9�~ ��Eg��XQ  �-�릷���@_t������`��M?��9f@/� ��Yk�� í^�'bz;#� z�@�7�E�W+��$ ��	Z~.B�ʗ�� ��@�W�z��)d+ :�j#/�a�@?� ���X�ā. ����k6��X��s �D��+3���� `��ꭂX�@�O:��3S�% �H�Z�ns8���7@�5��8VL��| <���0���]��3�9f@/� �P�Ԋ���  ^�R���s�t �F��B�ZO�KyO�N  ��4�����[�}���JC� ��@`�V�U̎� 0����uG�/4��`t@/� �Q]�����+JB ����l=?���:��#�X�l�Ӭ6�q�� 0pj���G��m�܈�)� ��@`�j��ɕrN|	 ``�~�m��֍��2��D�K ��@`3�ި4FX� ����X�ms�%��:��#�Xg������� {n����Lo7q�@�� �T]����9 $��jq�b����:zn�$ś� ��@`�F���J���r� H�f�Y
���-��u��pD� ��@`���Jql�8� 	��ȭ��Y�����)IU ��@`-sV�Y��ʦj H�z�>b6������w~�x,��u: �U�����S�]�d��0S��Sb��=7�*uT ��t V��HU�����  �2_)��.$�S��G ��t �3#0�B��  !��ƈY�$2q����Y��2� t� *s���ꉖ�s1# �CQ�֍��]{n�����X�G�.#�$B��Qi�fGr �Ve�2j��p2��H�T�s�κ @�� c�����3�9�E j�Z�v�m��v�BFύT�j � � Q�s呱�YQ��� Rfj{e��K]h���5 =A�H���b��� `����M�.tz��v2 z�@�8f�{*�ʻ��� `�f�16�SۗdU�� =@�H���ɵS-Q
 �o���3o��������v����� �$RER�]5�� }���-ϕ�b�厞{��z�G�. �:��2�)[��h��- ���ձ(��7<�E&Η;z^Ѕ� @�� ��Pɼz���Gf�ں9 "�i��\��t-wc�%y7wX �Gt ��zt�l�RH������! ��[A޼A*[���%Y�g�8 =C�H�+6\.f�|C~}�:U��>� @ט���g�^wnFΗ;��0�P*�?* �#:��ɍ�����a�K'.���-ΰ�; tC���c6/)2a�b��A����}� =B�H���_*���a�\���}e~�]� ��*s������X�87J�xD ��t ���2rњ���~�wݖW�ܷ��r�o�;� 	�(��Z���w]뢕�ھ$�
�
 �� �.^w�xn�Wan�d~j�u�/?q_5�" ��]k���մXl%��w/~�-��/ �C:��q�#������y:L�_��:�/{�G:K��B�M�P�/��r+�F6ʶ>��� �!@�l[�U���a4���|�����8���|�~�]��/��L����vcT� �1@�\���s�qZk5��,�d���w>� �9��03?37"�3���m����?	 �� Q֎�����9�DQ��f׌đ��{�{- ��9�|nfn���Ԍ�^w���JOMn}� @�� ����c�Hߐ_?��?<�`[  g�ŝ���=΍nĹ1���|�-� =F�H�����_wA����Җ�pmP~��n" NC���0�0��g��Xw�d��{�> �$��.��\����\4�}Tk)?y�I_  ?��5q���qޭu����Q�V�> �$B6���-�q�H�E��G�� �0#����1rޭu�KF���;�{�a�> �$�9��u��p�H�6�m4~���+,���4����^�����( �': 빎+��xE�Dzm��ϗ
u�!evk7��'������� ��@`��I.�[�� ���B1��L0\"��8�֦pKF���Go��A�>!�XM�����k�Ƒ^]���BS	 ����3s#I8J����Wc�U ��t V+dRʍt�kDQ���8�[�uB������|1)q���O��R��׽�͟�O
 ���j�fU��}�\��:�@���I|���q��Hw<7 @�Z�T�/�$!��c��&dr�o��o7 ��@�uf�#��=���A���r��?���b�Ƿj��)
�M���`��j͑�|%+	a�ۛ�=������6�>#�t���"-˙Ny`��8ҿ"?}�Ou5ҍZ����r�ˤ� I����kc�j=%	��87F����� �3@O�� ������q�K^��H�7�t8�|���U� pZ��ly��jw�
�e�S�� � ��gV"ҟ<�Wځߙ��:nW#����0�R�c� $������HR�Q[��8�D�`�+��@ �:��2��M�/���އ�W_~�v]������Rͱ�;�$�~�|b����ڗ���皒�w�f'��������.7���|��g����^͙��1l�\�g]: ۵����B%#	ӏ8w��G��o X�@�s+�G��?<G����T��Wuf]z&
�l.˺t ���S��L���D�77��ƴL?�띻v X�@�+�3�����������.d]��k��n`֥�Mqԅ� +(��l��B)i�͍~Ź+��p�~S �":��Y�H_�����E�٫~FO'�~���Z�,�
�B��t }����Oկ87���}w��� X�@�W+��v]������5z�誮_�)��Z-�Τ�S���r�<��)�F?��%���
 X�@�w�-�J-��VВ/����\o_��'W}�V�� �/���@τ� 7|���]ڗ�3΍�h�Ю��W �2: k��9�a�W���ke}�֫�W��(��b5����T&�N��2�D�Z5����Ŵ$T��܌��έ�} � �����>$�ͪ��%���Y�'���]�SA����f|�I�XQ�f�s������������#w���/ X��ϒ �+������ުɫ/�^�2��\����e?�h:�cFͫ͑��b��6_bK�;��jw���X��ϔ p�B.C���d6S9.�み�W_q����I�?;���n.�kq���(�pb!���-qn��5�����Y �Rv<[�i������H7;���ү�r��rӕ=�����	*�9F���57�y����R��M��y �� �f.���M_3]�������~Ŏ�K/֥w��0���� ʖ��%��'v��0��&�m�A�}��oz� �� �g.�L�/��t��c{e�� �_~�.�J=M�+��L6f�i�M�<:��z�>R��S�p��y.̶�\��� �� ��0����nw�:'����C^y�+��U[z:B�j6]�����y�M�� @̯�K��r.�皟��Ǩ��w��;_�s���@�� c)�Wb�w?����ˑ�#�'/�Iq�gW��֪V��S����e��1stZe�b���3�|�l��T����'��w $�}Ϣ p���)ơ�w�:_�Ǐ�錨�����#����t�d��\6�ҙt+��f Ι�^���k���nشܩ�H�Պc� $� ��
�r�ů���90�Բ���Δ�k�]�/[iO#�Dy���Z͖k��{)�'�q����NV��R�C���0���]oe:�a�z�S��u_���w�� @B� +���\��ç��=��i�Aȷ����;����:ɥs=��i�㤲���q��'��0t��f������r>B�h/���͗�Bc�u�V  At �_�m�J�J���G�����sOwFӯ��z����_u�Q�����X6%�O.����|�8�̗�(_:�FN��1���l it a��:�K��������x�����n�?>�O�ez�~Ŏ�I:����Y���\:���L�L` ���(]]�����}�������Z�W�`�;v}V  at ��-��^����C�ٳ���|�̔g��;^�7Nm��0Q��v�[>�N��\�͈:� �N�ʵR�V��,���/�E���э� H��{� 0�<�U���:�0�^�K+h-�������_�k.��n����]�������#��p��>�}��k���p�η�\� �'� ��U[��ȴ���rt�زo��'���ayɶk�����v���L:�0������y�Qo�uU��/Y-���;>�A��� 0�قz�^?rh�|���H��7�l֦�ѯ�����.����}�V��Ʒ|'�3��8�u��T����:�>����=8q�� J�%Ũ�xю�� H0�@3��_��rY5����{�QY�c:qH���+7^���t�]�w��ҩT��f��uB�5��ʺº�ֱ-�B��ٕ��/�9��}ߗ>$��D���p������Ϳz�`�S`h$� �azdJ����N����#�w/��̹��?�90���l�O�գ��:���}'�e]���l�W�j��q�j����҆l�����w�uͶkd�0������>��Lg7�ړd���_��_ H8���\O���ɚ�5�����r������%ٲj��v۵�����av�Qw�J�r��Ӈj���f�:p!�sc���5�5)�q_�������DqB��{Wd�N�%m�|�T8u�����. 0 ��, ˴ez�Z7�V�o˞#O���ū����엃��:�ޯ�t���B��"��Xz,=���b��H�H}ω'��V�R���ܦҦ�xn��v���
c�����ǿ�9�1)�8jnd���J&R `@� ��9.�.�N.Z�]�ѯ��h�Ҵ�'g��5[��[�6K�wW2#�*T޺ܺ��֗��f�`�Pt�r\/���)]�T�QXi$;�n,�/�-�M����j�K��/{��,M���g�$u��p��[��o��w �|F��flMgm����C�ȅ�bcQ̆t�����/����%Q��dnR��n{u[�^<"�O�v����*r�n6�l�VZ�[_Xޣ�/(.�+7^a����?�/+��f�%u�|�fgӗv�s�= �@0�����^t�l�ޤ���We�^^�ǝ]��O7�����H)W�$ԣ��ߓM���et��ԏˑ�Q�Y�֪cX�.N{K�
�Ң�k�jޠ��k���w��2S�$�\�3��|꽟|� ��!���GW�׽�u����<ԙ��\f��������t�m~Q�7�;Ui��N�tnZd����q9\~ZNTOH?���T���+��o(��潼��ރ?���������3u>ܷ�[f:�	�k~&ŰX[�Yu� � "���㪫��X.^��s$ۓ�����F:�Ǐ쑽���%�.�Wm�R2��5Wɝ��������X��Z8,��E��s<���&���67���L����u"/�6Q��_}�k=?�mF͍t�
6��^w���	   N��)��/�i���7�ƊM{7��z8������ŷ�͆ub��)���e��&�9Z=*��I���n�_�I�u#k3k
�s��c�Ė�-j<?����}R^��2(an���[���|�-w�P `@� �֍�U���_֏~T��=�CE�<��PvǏ{�K:��Ie�6AJZ�eSi�l�"�vE��sr�rL*����UH�Ԛ��tn:;��H�Jm����1���~���׵��e:���b�����c! 0�t 8�q�/�-�6�o�����mlvP��S�#�w��kv�s��zU�QER�R)�ֱ-��~'֏׎˱�L��CzE�S�)g*7���MeF�#^���5E��w|�<��C]����~:���o�ݟ�]�G��92����W�L��Γߑ��V��zT�f���kw�e.�b�(�2���f����j�j���b�Y?Z>*��%�JK�)Y5�J�S2���ԙ^:y ��?�Y��ȡ�];rm����j2�<������ � � �i�ȴ��*����z��2_�_��6k�M��~�Q�:�E��p��TJlfb]���c2�.��Tʭ��Ʊ>W����\g�<�B��%YU���8��sc�<���J�I-��w��=�X�޸2ann�2��T�z�|펫�^�F `� �nT��/Hy\���u�߼�u���O�w�>���bfTp�̾�m��*�j㕲ab����2����ݼl�$[ƶ�ٟ��We�Y�c�ǜc�	��3Ȧ�2Y����L�$�������+����̊Y�#Og�֙?W1,�/��v�Ϳz3�S:��[�[�#���^� &�0V;�^$[Wm��-�u��|%͔g���,�q�t�%�}ն��<O��3��Y��5��l(��+O��Ͳ�9�:V9��ͅ!#�C��)�D~\�� ��OH��J�(�m���c�և�wf��?ڵ��=̍�ε7�ֿd�n� "ɸ��hw�|�ܭ�n����'���� ��ԋ6_%�ۡx�Ay��c+>jf����o�{�'�M�K�^,�\I���
/�xyU��Bnsa�V�D�Vşo-�q��N�f�Z���*ù2���f'
2��yJ�N.�xƩq�A�wfҘS���a�|i:� �D�p}{���ڹ�1�!C�����C���;�{���7[nk`�{r��z�E/�m�	m6�z���+v4������q>�l�� ���D֍��~���DQ�$�h>�����Ƣ��Ӂ�r��[��\m.�k̇u�=q
�����d$;"#��7�O�?%y��\uN�)�{��]���07<�Ee/��;�sǽ Ch`/��烷|�{�?xݞ`�o���m5|�l*����b�|�e�P$�镞�n֩?5{�s+e��c��h�E�K�$��1Ym�7�48%��*�J�M�M�s]�k?4#��v�5W_ˍ��֪�$l6��ȸ9u`$7"�TA��b'�Sf��)��:J��-��@gm����~�a
s�ю��l��Λ��� C�@�Sw�z����7���O�m��:ҍgC}����Ïv%ԍ�fU��=���tF��Qm���%rT���({ی����#�H*�����f���_�G�v=�������F%Zl��Jk1b#��ȧ�R�$�	���)J)S�D��1n<��IfF��yB�������S[�n�;����[�[ `�� z����}ۇn��=����?�nd��N�_��2m���>�hW�\2Ǚ�}�s�g�}����MF�2HL�G�D{Z�^����
��;��N�
�aկ��v-��5��X��vM�A��(H�@nW�ݴ�ɥr��rq���x!��8��q�ɑ���%m�z��~y�ؓ&л���1�3r�=����o��� C�@�w����f"��8��C�F�3�~���������>��Z�����zgWys���m��vn�TFճ���)�+�bg�W2f�=΀��C	�fЊ�a��A+lFM�L���o�,�<�#��J�MI�Ku>g܌d���AnvO7A��o�r;���Kn�~\���0
����c{�����R�n�]�����E���|���?   @��H��7�֞`�_N0TCF��v�g�(��=��������}=�V�ܾ������[Wm�L���H�x7w°3�'�Y#�.�O����`��V��a��~d>���{a|O���#hK�ݔV�6?.���n��rt>�s$/����S�
�vMx���_^����H��7��'N�:o3~���	߸�Bhis��ޙ}b֗w{
�����as��n�#��]o��i� �@_�z�G?�oj�	��ۖ����%�|����������&�5jF���As3�!�t��'�wFW��٠.��7G~=[Kf:w�|�����9��DU|���7:#��~?���8�M�ǱG{�=~�����i/�Q���2��3��)���ک�~���?м�b��I9)e~�\'�>�R�g���I�W���LD�p��Y��}q�?5����޳�m�܌�3����-�� �Y:��3k�o��������o����}��Ҥ\�O�K�]#�-Oy�+�ԗ�s���߹��3#ꛦ6ű�n�F�/�	b�K�O��?�3�'�.vX�磟Q>���OǍ�h���mw��n� ��@`�]��u�w����{�o�ʹ1s\�9K݄�����ӏuu��a�p6#��fFi׎���q���� �Y��3Ǣ�?��̑C���=��ü��tҒ
���ް��]� ��� ��?��?p����߭���9���L?77���9����꨺aF֗����X=�J�Ol��e�0&����>8w��G�87�{�i�ϗ�2���E�t׭��  N�@`�]�ܵ��߾�棏��
5������t�K��/�٨�a�q]8ֹ}w�w;��f�����ck� �e�g�������Oˡ��2�8חc�-?���7�8�^q���  Έ++ ֹ��;gv�ڵ�[���9�f7�u������އ���1PK�ͪ<��c�����ℬ[ۙ�zt5�k�3�Ƣ<�p�3}݄y�v^?F�_�x46�Z�/���w �"�X��o4�7��}o�����/����+��y�@7GfE=�0�|]��=x�α^k��tF��ı>�tx��F�.G�f6�����f��?�a?"�\M�_���mozӛ| ���j���3/}����~.�Ô�$X�Vkn��uì�?p�@�fdSY���U�6�J�JS��㜙 ?V����L帔k�L[?;��;��k����}�e���[  �@`�O�㓯}��r׾h�[C1\���a�t
���n�K��i/݉�8���ȔL������F��W����	��c܌���@�Q~��_-�,�ۧ���+ ��B�H�?{���v�o����M���s`��L�7�F���Y#l6�2���/�ɏtb}�4�9���:.�>��?��zYfM�wn�2�y��9����Yz��ǋ�h���?��]�Q  �@��޾�����_����ߍ�Y��SG m�u�LW6�fnO}��}�rd4?�'K2Q���ℌ�%奈�2#���N����;���|_7t;��(g]���G�֖Ԧ_��ֻ8F .� Qv�e�7��u�ʣ����JS\I�'c}�E]
9���nF�ق6��渹��O�w]�����m�Q�J�r2�kq��!^��m˟��a��ʙԓG��̕w��9 \0@����;j�o��������^��r"��'��`�vs���:q���7�^��}$?"�숌ƟGr��6b�>�/�?+����#�^�J��	r3��X�j��a����J�zw�7?s�=� ��� �����/��#7��[�o����v=FS���-��#�&��Q['��z�����q�u�R������/şs�Ph�g���7Bj�ڳo�,>����0y'e1u�{<�F��mw~�ֻ�. �A�H��n�����p��,��W��_����gA���?��$���&i��/�B{"xԗ�Tn�}D@�(�&;�� vY����L�m�JD�B�E�J����V�T9�s<؋�К�K�dwv��3K�B/I��>3�����y��ln�$M����g�-[��W���Ȩi:2��<���5�}>|}��i~n1��%=K�b��z��8�v��Eq���{���4�\�陃�`�
�������c�����?w��>���ǸS�O�%y�z�s_��\�� ���@�۱y��v��9�w_����]p΅g�<���*EG���p��v:��j�ڛ��:�Gy�Bތ�޹h�	=���M�Bw{c��7c�����sc\���ͱ�}�V,v�bv�^ ��S?���L��ç�7��n�7z6��;�=�~6�O�������g�����xs>��F{D��9����'X��������� �Wh�֭k��S�Y�|r��=/:��B�W�'��#����Ճ��4#��G���pd������
�����?�k� 8!:�V�)]=r������߻�sO{ʏ�,����I�H��*�ē.א��������g�����? �0h;׾g�ߏ�c˿^���5���'�z���O����m�k�Y8�<-�K6�V�'.~�\��u�}M O�@��x6�<��9�O^�_���+�q�3��-~��Vv�5�#]�w�#OSw�zz�]�s���~��5���G '�@���#��ݕw_��[��\��5k��� p8Ď���7�Ñ���xkX�/�}Z�n��% p�t����;�v���;�;���]t�E�ȥ瑎�
���x�+����3n�ݑ�/ �t�;6�X�aˆ_���}�S.^��P=��G���w��'���!�~��e�Wg+_s�ȵ� ,�t�m�����ߘ\����}������b��.Z�Ý&��P?2ڏyx�G�O�q� �H�3����|��}�_�����ڵ���X���"����������F:ϲ��=�V��Qs�4t�c]=r��������V������c��b�R���G��c����_���١�ͱ(6
�3�3����� $C���k޶iǦ-���-�?��矶f��Ï8:|�0���\���ҵ��G+ H�@������p�;�����Y���~ړ���׻D�m�w�w������� @�:��{�u��;wn��_�˥k~梳/
��M��U�|m�����,y�5C��	 $K�eݺu3qx�Hu�y_��Kv��O<m�Z�����~ja�k�F��& �<��&K�7�a�;޿�=w��|qoo�P�כ����:�w��|�P �et��pݻw�o�Ν_���O�8c��/8��N�ԕkkoY�d�˜��z:�18t���F�Fθ�޿�i���\xޚ�B�����kU>x����%�]y����$�������qx����K��o_��9瞽����E:� ���+�;m�ڷ�6��2 ��:��P�8��qX=49�kw��S}�yO�_!ԁ����d��]k߻�];*�� ���������'._������]�ۿ�_�'̢�w���?���׾5 �V:�<�1z�{��+o���GN���g>�kq�"�̛�0/���.y�뇆� ڎ@�'��x#���^�ƶo�~���7\p��Kz�u�q[�譟Z\�ً�\�Za��:�<;�o������}�=˺�(ԁ��;�[_�ü_�t
�p�\z饳q���;w��ڭ_��╋.��l�<�E�E3k��~�����C�x�Ct����??w�{���]�j��9����>����Ƣ鵅S?�㫞�K��3	t���Щ�oknלּ���z��8�����йB�C�v��Ī��_;�� J�,�k�׼�R���=�o�{�]a���郧�B�:t�B��`c�۫z�su��?�{� �p`�����/L�����%k��9���
� �����X��������}��/ 8�@H@O���ׄ�;g�7���г�7�yڙaq�� ���3��dk�0�s�/n-�� �at���bX=�*�{C���w�����3N	�,_���%˳�tv`����_�i�e�/�t�D-͖��`��<n_�г�7��������t�6z�+��^ճ�׫�~y��M �@H\����W�����/��K�/�������cꐊ�Mߖ��XU�_x�7^z饳 ��@hY���a0�=!ܳ?��z ,�����X=�������O�^u�di���{�� <�u�ך�)aM�)aw�'�U�+|7�/�3��D+���`X~�`����ӵ� ����eKò�C#�aW|�5}w��lW��0_�n���߳�{�sK���Q]_�w��]�<� m�y쪰2��Yf��po�;យ{��=���8>ͻ<��}�W�a��wԮ�}# �	$��P1/�Ӌ��m�랙o������C�:<�,�7XQXq{_X�yǻv�U ��D���E�u^���pn�)�ý3��m��{�N��Nw�H��l�7�������? `t����
gϘ�f��۳�����v������Ŭ�/m�Y�-����� X`�C5�V�̹-��p���s׭��v����n�w__v�(���I_����= "���C�)��ᔞ�!��'�ߙ�N��Ʈ�`�A7��%5O]_�Xr`Y���,�^���zΩ �(��ɲ,,Kò��s�����w�c��]�@�7��'t��7�w-͖޼���7�._��� �����ʻ��2��^9��/<?�����	������y�l�ށ�ү��\35��� Z�@���_��Ϟ;���CaW���+ <7ׯs"u�]ai˲e���&�9����/� �t ����}y_��~f8c.��
4v�E{�Z���s���j��Z�XԌ�0X���aq|rw�T�2 @� ̛fP�a/�`�9s�����} F�����f�e����g��|�@��faE�������� �St N�ft�R<en��|K�\���+^r�1����>��ƃ�=�u�o6���'�K�kYai�aYqiX�X��� �K�p�m���8|���Ν;�o�}��y��]�v��e��f�����VVȲЛ��_�׎��_�����  O���֭[׼�܇m?����{�s�[6�T��f������.ٞ�bV��E�/�x_�/,-���-�Ǐ ��: �z�[��oqxߡ��<�����<8�����=��.L��d3E�~b4C�'���E��Z\XC|`���
]��N�X�c&�h9�����C��~�/����gg^ppf����gN����P_<�8�;�5[��w8]1���ߏ�lQXRX�dK�?/.	]��G�F܊�&�h+�_�=�?=�=���=��C^P�ן9ݘ}R=L�����0�Wo�,���=�a��^�Y^h���5���sa�sī�phk����Sh�zB!/<��q 8�: g�7&�5������nذ8�;?����������3�~�L��j6�/o䍾P�{g�=y1m�1g������Bb���sc�1W�͏�� 4�K��'p=�Y��(��,���y�P���5�f�V�*t�;�U���݅�}py6𪮬;ď��!=~<ŹHL��� �v: <�m�n���mIںu��F�񪹝<����s h)    �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �    h9y�� �f: �r�,�T*}�r��  mB� -�P(\�[ �	� ��F��� �h# hIY��*� �&: Ъ�^�V�_*�� �t �e�y>�@[� @�ʲ���5 @�� ����z^(B���za*���X� �0� -.�LOOO�T1̟_���� ��: ���K�<p�@�dy�oߺu��6n���  -J�@��������Y:T��W����^��s�; �J�@��W�������b��<��eq�# @� ��<�/jG�![c�ճ�hE �@��;�pA�pq��<����۟y�W|' @� ��)n/
4#��z��'ccc/( @�� �b��S��7��;00pC��W7�� �: ����vI��ŵy�;��
: �����ۻ��?�M�j�_�xe ��	t h�7o~�R�ܕeٙ���7c��T*�N ��	t h�=no	��<ϯ��j�2 @�: ��,�>�ÊkSl4T�V{J��G $H�@��)n��?��y��R���� H�@�6Q*��V����<�C���Z-�> @B: �����*�š��?#=�t R"���|,n�<��G�+�J�\.�A �t h#16�)F�Wb�>'�X����~�Z]Y*�� �@�6��������š#}����減 X  �̒%K�h���[cl���h�V;ull�m����  @�@�Y�~��J����3яכ����7 p�	t hC�b��h4~9x&���������HU��= N"� mh�ƍ�W��O���맦��??11�s���� 8I: ������*
�<t#4�C\�/�799y����W � ����譕J��8}Y��8�P(�M�Z��R�tc �L�@˲췃@"��g1�%F�G �@ �X�ʛc\�I��&�x��y���J���r�� N� m�^�_�����8]x\]�?V�V�X� �g �ܦM��aY��+O�[���s�����<���&��dY���\�8�xB��xff�[�l�dӦMw �' :�����J�R��O��Ӻ�������r�� �� "��W����?�ggY�Ÿ��,�J_ �	t �,��<���k�aE\Ͽ�T*����  O�@�R*��V�o��O�E�e�1�?^��.� �q� �ab��Y��?��7�E��b���u=7��  ��@�T,/���}a���O��J�߾}����7 � hÆ߫�j��h4��y�v`����l```���؛b�� #� jxx��J�R��k��c�b��Q�p�: t�r���Z�>;��D���;w�|úu�f <� .���Ȳ�qzQ`��n�޽����^;44t0 ��� ������j��1ԿC}y`�]233��� �x4 h>z훕J�5qzc�z�����7�����5� <� �)�˟����,�~/0�⺾�����1��#� x8 ���#����.����<��8� A� ?d߾}�����'�[k���8n p� ����וJ�Y��w�8��V���J�� �� ����k����y��q�?N��W*�]q�?  t ��xi�X�b�=7p"옜�����ȧ O� �htt���/.
�H?50��,+��c�J�g���� :�@ ���ȿT�՗�y�����mI\�?ݶm�s7l����%���T*��qbb��.�wW�۩�z�/��ꪟؼy���$��c2::z����%�B�Ƹ;�WY�=����O���^244t0 �q: p�FFF�\�V_��	"�Dx����������#���R*�n�����,�>�����k�˕J�o���u��"���622�������"���>11q���� C� �K�\�|��`1қG��&�gw�P�d�Z}V�T�+ �: ��H���/�������&�皸��{����C��'��'���Z��3�F�fT�M\�h^��� @�� �6<<|����='���|zs�R�B�\�� @[� ����1$��eY�9��M\����722�� @�� ��)��w�j��5���ݟ�/��z~lll�ٮGh_ �W��û*��K���q������~�����8}{ �-	t `ޕ�����^�������̗_�V�]*�> h; 8!��ǧc��R����H
̋<ϯ�������ȿ ڊ@ N��8\Q�V��r[�,���%\�?��~��K/� �� �p�Ri�V�=#���0_<qϽ�;��c- �6� 8)�����T*��'�,[x�޿u���lܸ�� @[� �IS.�?]��~&���wW�,�z���;w�|κu�f -O� '����W�n����w�<�ػwo9��9 ��: p�5O˞��x^�XlF���[��W�j�O� hi X�����ر�'8��{I�qi��޼�����s�5�%���~��}7�pë���q���׳���~5� �,� ,�C����j��M�J��m�T*�*��� �$� $�g�7���K���vq�� @K� @2=+��8�/18��כk���q�G ��t  )�r�s[�n}~�����{V��5/��|�Ν;���� �G� �i>��V�=����؜?8�޽��8n �� $ixx�ߦ��^033�ɸ���1+
�ٶmۇ7l�� @�� @��������]��߿#˲u�c��^�o��h �et  i����8�z�R�V���c���fו��; -A� -!��D�{��a���x,������) �: �2b�drr��1��8�U\�7LLLl�5 �<� �������j��y�|����)�ū��� @�: �r���oٶm�O�����,;=�h^R�V�W*�n $M� -iÆ�#���"�I�G��y�� $M� -+F��NNN�d����+���U��g�J� $K� -mdd�ޫ��ꧺ���"��s��Q�� �%����y��&&&^R(���������[�^�q��� I� @[�#��1�?c�y��fgg��7 �$���ь������������?*��/lٲedӦMw �#���244�'F�˺���7���G�*�o����t ��lڴiw�����l�e��ק���?44t0 �� ��C���������s�,[=33Ӽ��G I� @�jFz�V{Y���=�>=p�eA�$G� mmxxx����K�����e����nݺ�?mܸ�� �� @���V�]������)�0;;��8t��t �#�����
�����B�˲�ұ�����ǧ I� @��z�V{M������������i? H�@ :������T*o	߿IZ!t�7��� t�r����Y�]:X��_�e˖eͻ� �@ :R�����yq::עb���8~$ ��: б���;200�8�$t����� t������������q�?��e�O�ر����� J� mttto�Rye��cuU�<=������fq N� �\.�Z��R��E��;��l� N� D�R��J���Y���?� �@ 8d߾}�������/��܉��GGG�g `�t �C�7����z����W��i��dY�<�]�, � p��������[�<�1Fk:D�P��8l ,� p�R�tS�R�.N/"��g �@ x���xQ�^:@�ek�l�rƦM�� ,� �0���������_�S��³� ��@ x###_�V���_�P��I `At �G�e�H��xeW�6�:t��%� ����j���8�`hsY�=# �`: �c8묳���;���������j��� �t �1\z饳�J�q�����<?7`t �cP*�>Y��6���C˲�8�C ��  � �k^�T������A`t �c���s���t����.��@ 8FCCC+��G�ڔ#� G� �,�>�8���7 X �8�V������� X �84oW�V?�o�I�,� p��<���m��s ,��@fgg����j�/�I�P�F��pOh_��,��@6mڴ;���eY�z��zw��ٽnݺ� �I%� �S�T�9���yw��ѿw�������o��@ �\ �E�_�~���y6o� 8�:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $����$%Gy>*    IEND�B`�PK
     t$v[	^�G�  �  /   images/9ba3df0f-d630-43f7-8169-617793654d93.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  sIDATx��	��yǿ�sfvv�ОZd����XĎ�;N�g[(���p:�w 
`'X�B�1�������#��:@ ����c��9��|_Ϭ4ZV�EB=5��������]������Z�JU ��
D0U��*�T"��@S�`�LU ��
D0U��*�T"��@S�`�LU ��
D0U��O]�f���� 8��S*V���F���!�=�J��@?��)�������w��ςfܤ��%�c"�4�w�������|~R�o�p9����ƽP	Ȣ'���y�q/����;	+��j�����ܬ	K?��`Bq�� ���}�|a��Ȗ/�p��W��i�>YB���E�h4�nmlj�'��<7���M�ŏSV<��G�Y^�O	
�YNg|.~xE���#�5X����0�~n!�����AD	�o����9t'{@���S�v^��G�1Y���eC���#<����g�����)��>���=n�lX��"!���@=��A����R�󼻗�E,Ə�Xl,�X�� Z��JG�C�����F�o{�#3�e�u �������ֲ݀cG]wh�|],(er�Ӌ��M�}��/�}7ƅ��#�
�Vl?�E���ɍ�:�������lu,�reI�p���,i˵�OK��DKy@ K)�eO^9%[���:_��
#e��>^��?��� B��N>��ke,RW[Wbb�D��=�~D�b"�����;��N��*����Y��
+���a(������ ���j����gƷ�ho��l+�2���%y���l0On�k�7���xRKJgM8���f��n�z3�$�*�riC��u[v`����=ʭ� Y�fq�-����ƹ��2|>�i�>��+��
�j�.����dw��
ZɎ��;��v6LҦ�N�k��(��4�X\�K��|=���ZR�^l_�0�-e�6Ct�Ȳ'�AF͇֡z�El��-(��S[N�u�vQ��Fˀ�s�n{5Gq[O���n�{����g'�U�P�kB����;^�c�� ���|�����;�*�P�W^�9ʶ�$ M��� Ŝ�*lR�$}z��8Y�P�]�5jB�������0@s���D�\ܾ�>o���;���:cg|MVY]�N�V�����h��I�.�-^KE���v��P����r"�*�!ޠ�l��m��S�܏�|�-/��g��������9��Zb�<eh3�t��+��֒[�f	�7�|Ic�@=�z����JZ�|(������=t-�C�~��ֆ=M
ڇsY�E��������`]��LE!�����PNE
���0v���X�!�NI�H06��dmؽѤ����(��a���O���1��~+R ���i쭉��
}Ra��q�:+�G�"3�m��޸�mK��n�cyh��`Z.n�@w�梧��}���m��^�º7v�ɟ�oy��!���S0��܊�������1�A��N �ϣ�z�K�	��s`�O�
=�V�ͩ����RwEV�u`�CA�p	�(t[0Ǖ]H8q(�"��*X��j?�7���q�F��QEր-�`gf�C` :��'%�DƲ�Hd@�?����(�
L�FKJX�����i?BQ>��3����l��,H�5��*L�TIe�����0�9� 3iN��DBwʺ�L��F���>��Y@�J��Ѝ�%��d�NʨȀP@W=� �R͜C���S�"�C�Y˕���R�`���x�$(�0o?l��X��N��;%�u5Vܷ�)4pB8�VwG���B�B�T<��A�kyI�h$
��vʵܸ$K~�9Ս�*��ɶ협1t3c�y��Z��sT��$I�U�	,1�ൌMb�6�V^H�]�c��"��D_q_��Y),���<��u\��<Y����?�ӌR�a'���AH ����%�����D/�$kpL'a����A
�ш``�ɮi���`���/���O��� ���lL��8ʵ]=��7cs�U���>�Xڲ,	�SL�X�V3��TI0H��A�4)�A�ف���P�(�8U:���R����4O�.������@���stS�讜p�R���~N�C a���}� �1TS	�� C
a����s�3˴�X"��Uv=׃���5���^��UV �uϕ8r�-&3�5�|K�1,��C�ـ�M���ޡ���S�zl�Q0�@MM�-�i!'����H��^���2���D���
�V�⺮$�Cs7P$E6A��᬴Q�P�@��_G;�ԁ���x1����ZMm���Y8�8������6&��iy�VY�Pm���]8T?	��2�d	����oC��y3r�JP�@Ё��j���/l��\x�E�۟��)��g����Wbeo��R۲�XL��r<��mnز ���bю����x�TtU�p��Vn�k9����凶�0��M��c�1M:��)�u�m��sgI�e��?�D������d�df_|`.>�:��a�w���8"B�i�f�3�K�\��?���R��Xp.�W�|	a|'�Èn\��C2U�l@PA@�K�(�i�6\���y�I$�Ӱ`����c��ޒ�(h,��M{�vWmd��qa����ވ�K�2Y��,g�i�1�塐��C~G	�RG�pe�Rd@�����EX�/�H�<��b,\������,�rP�`�A�.����0s�#������!*E�ʛ@)�k;���A��n�Ƒ�W]}}�0���.�L�2,�G�����G�i:D�%)���[ x�*��UEWt
��ذ��.Y��O���(�G
d�;A�(ad�5)�.+
�3o�=���[G�#!�����X"B��ѐN�ǰ�X�! �������u`����oow[ Ƣ�y�v.�<�j�^���!(�Ԝ�Q�����!��B
���*�`Bt3ܢ�\t�p���x-t�t2��:��K�E�1���C}�u̇`H��y���&A�Gv\�Q҃�pBm+��<���->�sC�GGa���AD���\O��gR�?�\pUd?�қۂVx����"�\D���R���m_3�Ϟ:���p\o,�;LV���'ue����$��5*�D>�K� �`��
��K�8i�{�b>�3y6�������)�;��l¸	��[2�Z�ף~%Z�/�v.������O�
��y���t�b;{v&<���4f�!�Ӻ� s�	����q�6�0�P֨��ul��Y���7���~���[a执��T�ڤ5՞9��DO��A03���
g(@�s��nA4Pb��Mz������ښl�u�vēj���_o�|���)�n�Ӽ�u<uc��aYx���nߒ��!\��^}/��ϦT�;g�ɭ��ֶu��ͩf8�����]�L�0]��`r�P2v�3<�w|'\���T$�������0�Hh5P�Po`)���*?m�a]�:���{��
(���hgY�$��5�Utk��b�����6�UAׅn)�!O�9�}���Aظ�mxi��ɂ����7��q�qjKc�J�HhQ�a�<�(��h�Sr<i{�Î��|_f_��?Qu������w�݁��&�������}��S�)�ųϹ�˻[Ͻ[���
D� L��4زwd�,�w�oc��'c�6�YBK0]�hŸ����`9&�<62�5�`8F�n#Y���~��TXs�������ƣ7<�Pd@�\~'\�����`#<��0��y��_O%S��;�*��Н���h&U1����r����h��X��s_�-�"@Vd<�O�~�t\+�������l�����Q(�"�߿����۞����Bx��o|�G+?����<���i�6ih���J
��я�acyL��(磓�7��7?�TY��z��Bz` &�8	�r�7}t?���l}����lk�Y������Q��=�vc#�Y���9�o$���� 	������%����*ҷ>����!�u����>��,gH�`�>�y�ǫ�?,��Z�F�� l>�-�	lA�<�^tf����0#��|ӏ@�}��m�����x�� ��a��O��@ ��&�v��0ض��.��	Xݴ�S���Dcz��$l)A��!ɒP˒���d߱�?��ҙ�,x�} u2���Tv #)(�kL�L������̻������0_�D�m�6��L���@���.����1����BK	09����A�T߽�@d		�T�~�9��$O�t0I� LʒMফ�`�|������a����o1�~*A�)Փ7>�����ܨ�)l�UQ@�?�
D0�@ȕ�-7rm˗/�u� �0��)꼺�����/@�X�B�N�
,�a	'x���PW#c�����F؄\�cXh��7����t�RM��n�;�K��a3:χ��a���p�hU��uPG$j7�+��=�����r+��}U<�e˖�[�`�+,��'�`����!��A�x $��(4���x�C����G�z�q�4������y��S�_��L,Y���B���yXh��H3nN�Bͬ;DZ���B�~���X^�2Ҙ�+��B��+W��k��ʭ�i�MX.��+����&�W�<.����P��xn�0(o`�ˏGؔ,�qD��B>Q��͖���J��[z��*|:��
]����@�A��.��1��;p�3�����i��װԖ�_:�}	�����)a%�c�,_.V��hHUT"��@S�`�LU ��
D0U��*�T"��@S�`�LU ��
D0U���W�cfrJ�    IEND�B`�PK
     t$v["1^FHo Ho /   images/e2a053a3-24a6-43e1-ac97-395cbc045e87.png�PNG

   IHDR  �  �   �r��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���1mA  ���+w!`0�t ^z )�-(R^$E�}i��_]���s� ����\k�       ����|��5 ����cp{��朏��s p'         �%�          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     ���<F��~��k�fq�\��PVeqU������T��T��aIl���6�4���%��5�j)mm<j�j����J�"" �s>�V��@X�3�x$��?;3���_�y}     � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	���7�o�=���������r�l��ʲ����1(5���z��7       �Z�vm�1�@����}����c�3?�7�۲7�S���?p��͹.x�%K�
���q�GF]]]6={��#�8"�u����o����///�~>�y�>/         ��k��o��F�ڵ+���Ν;���cǎؾ}{6���Jl۶-{=I�~s
^E UEEE444dӫW�l���ߺ���UUU         t���ټ�bڏbϞ=Y�e˖x�嗳s�l޼9���g�>�;�\.�썍�q��G�QG}����޽{g�         ţ�����z�󝝝�u��,tߴi�[�q���}���������������c�9歨�v         `��r�^�ze3x��w<�w��x���^Ȃ��lذ!����ަ��>�?��8�㲨=���#          TEEE{�ټݫ���ׯ�b��������6x(UwJVuuu������          ]�{����ܜ�~�v��>�~��l�}��رcG@��S2�8�,b�O���������          HEMMM455e3al���/�O>�d<��Sٹm۶�b%p�h����'?��2dH�766F.�         �B�o�d~�<���M�6e��ڵkc͚5��+��;E#�����YО�UG>j///         �bҧO�lƌ���y��,t_�jUv�ٳ'�P	�)huuu1t��lN<���          ����!��ڲ��������}��ձe˖�B"p�����/ZZZ���'>��z         ����ʷ��mذ!���X�n]tvv�L�NAhll��O?=N;��         �ֿ�l&M��ms��b�ʕ��3ψ�I���d����)���E�MMM         ���իW�;6��_~9�ꞏݟ~��T�IJ�޽���5���\.          8�����7o�U�V�_��X�~}��$p��ѣG�1"�          �NCC�[����?+V��Gy$��]M��a���>dȐhkk�SN9%���         �ë_�~�L�:5֮]˖-��<�����t�#�<2F�g�qF�m          ғ_f��ܜ���۳����}�ƍ����C����[[[���,          (=z�c�f�nݺ,t�Gb������C�gϞ1r��8��3���>          (l�|6ӧO��+WƟ���x���;�	'��ƍ�aÆe��         (.�����֖�ڵk��{�������q�9(�!�СC��sύ���          �42$�M�6e�z�سgO����TWWǈ#���}��          JS�>}b�̙1q��x���O�S������RWW���q�YgE���          ���)S����_��{^z)�����Y�����ڢ��2          �TWWg��?��X�zu�}�������;Jccc�{�1r����r          F�=mii��g����+�zꩀ�"p�}����ĉc̘1QVV          p�����_�B�Y�&�׭[�vw�S�޽cҤI�v          ����2dH�^�:~���Ɔ��C�^�b���q�gDE��          �F.�����:th��o�%K��K/��63����7n\�;6*++          �B>t?����SO�B����7�iӦ�4	�K\MMML�81۫��          �����a�b���t��رcGPZ�%*�`�ȑ1cƌ�ѣG          @
***���=F������{��A�^�\pA80           E���1}��3fL��W��U�V�O�^Bz��ӦM�6��7�         @����W_}u�Y�&n���ظqcP��%���2Ǝ�'O����          �B����_}<����t��عsgP|�E���%f͚���          ����<[�<r�����<�@�۷/(�"�����͋N8!          ��t��=fΜ�G������nݺ�8܋L�[)�sNL�:5**��          �����c���q�w�믿6t���^x��	          � ��E[[[477��ŋ�'�
���TUUŔ)SbܸqQVV          Pj��k���+W�/~�رcGPx�N��s�F}}}          @�;��bРA��_�:~�ᠰ�TmmmL�>=��          �_=z�/�8N?��X�xqlٲ%(�4|�������.          ��6t����W�w�yg,[�,:;;��	�HMMM̞=;F�          ��֭[̝;7Z[[cѢE�m۶ ]�1p��X�`Au�Q          |4'�xb|�+_�[o�5V�Z�I�������<yrL�4)�          L]]]\u�U�|�����c���AZ�	�������hjj
          ����r���'�pB��'?�6��'jԨQ1{�쨩�	          ��jll�뮻.�.]��sOtvv���=1ݺu�9s�Ĉ#          8t*++c�������-��[����=!������իW           ]#�_���ӟ�4�x����'���-f͚�          �juuuq�5��=��w�uWtvv]OM}��ok0gΜ�ԧ>          ����b	�����rK�ܹ3�Z�èw��q�W���          @ZZZb�q��7�ƍ��#p?LN>��������           �ҧO�����zk�X�"��.��m����cڴi�5          �������KcȐ!��_�2�x����w�����袋���5          �����G}t���?��۷��������/����V          @a4hP,\�0~��ĺu�CC��������/�nݺ          P�z��_��cѢE�bŊ���bcƌ��s�Fyyy           ����2.��hll��K������r1eʔl          �Ɀ����;�#����C���".���1bD           �i�رQ__?��c�����'p?Ⱥw�W^ye4(          ��6lذ���?7�tSl߾=�x�QCCC\s�5ѷo�           JÀ�뮋�}�{��/N�~�80��ꪨ��          ���e�K_��o�9�|���������������           JSmmm\{�hѢx��G��N��1><,Xeee          �����lyvuuu,_�<�h�C[[[̝;7r�\           ����y��EMMM�w�}��'p?@���1k�,q;          �.�������"����w��#p? &L��ӧ          ��9�󢪪*�����	�?��lʔ)          �a�lWWW�m�������&p����"���          �����=���c���"��!p����b޼y1f̘           8mmmQSS��rK�����	�?@>n����O?=           >��ÇGEEE��G?�������r��vq;          p�����%�\�E�����K��?���ٳgǘ1c          �`:��Sc�����,:;;��#p��M�g�yf           
�G��]�v�m�����{�:ujL�0!           ���:+^{�X�dI p���>;&O�           ]aҤI�{����	�ߦ��=fΜ           ]鳟�l�ݻ7���(e��o���1k֬           8f̘�v�e˖E������5�ϟ�\.           �|�<w��,r��G��|�����^zi���          �ᔏ�/���رcG�Y�&JMI�q�e�Eyyy           � �7_q��o|#�{�(%%�y���}.jkk           %555Y����=�l���$�����ꪫ���>           RԳgϬ{��7����z��������K.�          @ʎ;��⦛n�}��E�+��}�̙1lذ           ('�|r̞=;/^Ů������Yg�           ��3Έ_|1���(f%����Ĵi�          �������'{�(V%�80.��(++          �B���b���o}+���E1*���G�q��Geee           ���������o��[�F�)�����<��޳g�           (�%��N����v�ݻ7�IQ�3gΌA�          @1ijj�iӦ�w�Ťh��#GF{{{           �s�9'6l�?�p��܏=�ؘ7o^           �9s�����c�ƍQ�.p����+��2���          ��UWWg��׾��عsg��
�s�\tttDCCC           ��>}���_�������3
YQ���g��O          �R���'N�?��QȊ&p6lX�{�          P��N��ׯ�����Q��"p����V��r�           (E��z��q�7�֭[�|��.���֭[           ���ݻg}�w�����BS����ɓc���          @Dsss�}��q�}�E�)��}��1iҤ           ࿦M����?cÆQH
6p�������(//           ����"�o���سgO���gϞ}��	           ޭ��1f̘��v[���O=��=zt           𿵷��O<�V��BPp�{�^�b޼y          ����r1����b��푺�
��܋.�(�w�           |��������w�������
�'L�C�	           >��N:)������L�޷oߘ2eJ           ��M�>=V�^�7o�TD����b���QYY     ��ػ�(��;��)00�.��4�R#�A��c�&z�9ɉ���$'�����I�;!ш�b7�=XŀH�D�I�����DQʔ;3��9Ϲ�/1̝�e���     _ݺu��+��o�1�����Z�i~׮]          �#WRR���_=rQ��M�6���??           8z�]vY̙3'6o��&��+��"�ׯ           ��%�\����"��t��F����7           (?C����z+f͚�$g��+��K/           ���_|�A���F����=��5
           �_������Ϗ|0rEN�%%%��{           *�i��3f̈�F.ȹ����(������           *N궿�������سgOU�qr/p?묳�E�          @�;��c��SO��S�V�%��f͚�g�           T�s�=7�x�زeK��9r*p��⋣nݺ          @�)..�"��￿J�9�w��%           T�#F�K/�+W���?CN�yyyq�e�e�           T�������K㷿�m��r"p6lXt��1           �:%%%ѷo�x��w����<p�W�^�w�y          @ջ�Kb��ٱ{��J��*�ǌM�4	           �^�V���N�g�}���J�}��          �i�����cӦM�z�U������U>D          �O�W�^�w�yq��V��VY]ޥK��۷o           �{��?�|�^��������??           �M���1f̘7n\��g��%%%q�	'           �k������OǊ+*���$p?�s          �ܖ�����w�qG��_��{��nݺ           ��_�~ѩS�X�dI��W����}           ��ԁ�3&n��
��J����           T}��Ν;ǢE�*�~*-p7�          ��:��s㦛n������}���Ѿ}�           ��9���{��1o޼
��J	����Mo          ���?������+��WJ�>x��8�c          ��k׮q�	'�|P!_�R�Q�F           ���ѣ�o�޳g�h߾}           P����+k�W�XQ�_��w��          j��O?=&L�P�_�B�T嗔�           5�����G��?��\�n��G�����           ��(,,��#Gf�{�~ݨ M�6�           5ϩ��O=�T�����׬�����OϪ|           j����6lXL�:�ܾf����ՋSN9%           ���8�x�����\�^��#F�����           5W�-���1cƌr�z���ȑ#          ��o��ѹ����y��          @�שS��ܹs,Z�訿V�rJ           P{��<���-[�	'�           ����z(�m�vT_�\�#FD^^^           P{ԩS'/���Q}�r����c�С          @�3|���	����M�4	           j��;F�bٲeG�5�-p?�S          ��+Mq�ӟ�tğ_.�{��ͣ��$           ���&M����#��r	�������           ���_�~0 ^{�#����S�~��'           >���޽{GӦM           �t��ڵ�U�V��u�>lذ           �}N>��x����*p/..��={           �3p���4iR�ݻ��>��~��Ea�Q�          �i֬Yt��9.\xX�wTuz��          ���޼���FIII           �?K��C=eee��9G����?


           �Y�ƍ�k׮1o޼C��#�SM           3`����5jݻw           8��?��QVVvHD�{�����           ���7\}�ܹ���G�80           �������&M�D׮]           �H�������={�|��v�>`�����           �"6�����={�~�a����           8T�{�.���~��ѵk�           �C���'~��V�ޫW�(((           8T-[��֭[ǚ5k>��+pO�<           ��={�_�����Mp���m۶^߾}{�ݻ�S�N)**��z�YV�^�          *_�ѧM���sȁ{�Ν�A� Gc׮]�iӦ���c��ͱe˖غuk��p}�J����Ǝ;b��ݱs����={����N�:�J�{��������ׯ���o�{�q��ѨQ������u 
         �w��{�%<�C.�N<�� �ϓ��6dk�����/jO�zUK?���I��*E�M�4ɂ�f͚E��ͳ۴Z�h�ݦ8         �?u�֍nݺŜ9s�1w K��?����裏b͚5ܦi���)�W�>��4l�0Z�j�[�>���c��y         ��z��u�{
�:v� �7n��U�Vp{�S�k�-[�dk��şz_��޶m�l�k�n�m�         j��={~��)p/))���� �fJ1��e�b�ҥ��%KbӦMA�HS�Ӛ;w�oO�{�P֡C���{Zyyy       �^�v������ۣ��4{yϞ=��;w�ݻwǎ;����y��ԩ��}�ի�@�����������կ_?�ur= G�c���-[�ڵk?�������# �RX�����hѢ,hO7T���ͬY���O�F��S�Nq����_�       �����6d���͛��~��[�f�z��sɾ�=ui5l�0�6m��6n�8{9�k޼yR�@-�����⋟�>�;@VVV+V�����g1{Z�ׯ��t���{�e+I�����w��%�u�mڴ	        ���}͚5��裏�f#��7fa{��^]�&�ɻ����f͚e�{�-�պu�hժU�� ��Q��J�!@�KA����c���p�;wn����c�޽�z��l���k��҅`��޵k�())�:d!<       P�R�����=[+W��?�0��S�^ZZ�#�Ok�ҥ�z_�Ҕ��(��]�vѶm�l�	� �\�wK?R�Ͼ0p�޽{ ��V�Z��~̙3'�����I��f��V���J�{:���O�vA       G'M+_�lY6|0�i������5�[�.[i��'g�{��۷o��;��c���( ��4h�=Ƨb�L�P�lٲ%fϞ�E�i�c���6o�o��f��6m�d�{Z)|�[�n        �-E�i��%K��im۶-�<����O~~~�Aw�q�J'�w��Q�PMu��M�P]�ݾ��n���{1o޼سgO��Jǟ�5mڴ�S�Nv�K�޽����1_       P��ر#V�X���,�ŋg���=iZ��ի���odo����=MyO]D���� r[
�_x�O��s�F�E�֭�ʕ����}�̙YԞ�a��k׮���|����}�{��      ��n�ƍ1���+��ij;��'���ӧgo+..�B�N������[� ��!�n����b�����E�bƌ��[oŦM�*Zځ��SO=�Ms�ׯ_0 �t��9        5Bj0� �>� �׬Y�l۶m�Y�fe+)**�Z��D���C��#7n�Z������܏?�� ���޽;fϞ�E��	���������c�ԩ�jڴi�4H�      @��N7_�`A�ϝ;7�-[fB{-WZZs���֣�>��;w�b�����T��x|X�{� �W�`Z�pa���曱y��\��c{��լY��߿6�=�       �&�qi��{ｗ��i� L
������-[F�^��O�>ѽ{��S�N P9�@��ӧ��ѡC� �|�Z�*��׿fQ������u�d�c�=6C���w       �
eee�|���Q�ҥK��ڵk�Lq{ ػw�l`ӦM���Y���o�>�֭ ��۷�[o����ij;Tw+W��?�����#�dGt:4N:�$�       �p�v�9s��̙3��wߍm۶����l�t��z(�,�N�O}D��@�J�zQQQv��>�Ӄ2 �o�޽���^{-�y��I/�4������dS�O>���رc       @y�Ϙ1#�0v��PYR�hѢlM�4)ڶm�Mu8p`�2 G/???:t���������5�Óv�I�S�N͎-��"���wLWz�p�)�d�{�U       ����,>����>}z6���]�*�^�:��l�݇�Z�
 �\�N�-pO%< _l�ҥ���/gU��Sۥ~��4hP�92�=��       �ϓ&e/\�0����o��͛r�'c�4pȐ!Y+Ѹq� ��w�q����{aa��3 >G
�S�>mڴX�re JG¥�iu��=N;��۷ov�       �f͚��_���6TG�N�4)z��'�|r���'


�/�σ�?3po߾�V�ϰiӦx���^�-[����͛���-[ƈ#b���ѠA�       �vJ�g͚�M�;wn6�j�={�d��*..�ĩ������ �M�6Q�n�عsg��g�L�dɒ��_�o��v�D8|k׮�ɓ'ǓO>��TNS�[�j       ���H�g̘���5ٶm۲Miu��18dȐ(**
 ����{l,^�8{�3��P[-X� �y�lW%P>v��S�N�iӦE�޽c̘1ѩS�       ���7���矏��FK�.�֤I�bРA��|������{*�j�t��{�O<�D�s��{m߱\]�t���:+���       T�W�Φ�O�>=�o��?���Z��0 
��k߾���?�Q�m۶P��޽;^{�lb�ڵk�<i��m�ݖMr��W�}������       ��H���Ν��Ꝇ�ׁϖZ��z�8����N��M�@m��~�S�{z�,..��"��o��VL�2E�U,��0v��h׮]�y�1d��;      @�+--�7�x#���lr;p�6oޜ�L�?i �Q������&5c�~�;j������'�x"6l�@�X�jU�?>��K�����#???       ��q���˱m۶ �\j�f̘���ݻg�DϞ=j��F�F���?w��ٳgO���Yؾq�� r׾���瞋��;/۩      @�Z�v���}׮]��y��e��c��ѣG��c���>��m�6 j��{���o��<�H�Y�&��cŊq��gGp]p�QRR       T����4��7ވ��� *�ʕ+����=�X�~��q�)�Dݺu��J�g�mڴ	�����ߏI�&������/^���o�G�q�Fǎ      ���hѢxꩧ�����kݺu���f߇��zj�5*�ի 5�1���
܁-Ű?�p,X� ��#mZ�;wn0 �[�l       ��}a��Y��z�7o��<^x���,tj�V�Ze��EEEѨQ� ��6l�O<�D���+vC����z뭘9sf�;��sύ���       ��,\�0�L��rϖ-[����_�"������kݺuv[��o����ꪴ�4�}��x�gb׮]�|{�쉩S��믿g�yf�~��QXX       �U�Ve��3�}i���ɓ�^j���q�i�E�:u��jٲe������PݤI�/��r<��c�7��ٺukv��ꫯƥ�^�z�
       �غu�⩧��~�ZVV@��&��f�^���>;��� �Mz�j޼��'�T7K�.��'ƢE���?�[n�%����]vY��      �O۸qc<��Y؞N������ǽ��S�N�.� ��� �M���`@u��5�c��M��Mp��Y�fŜ9sbĈ�E[QQQ       �s�ά�x��'cǎ�,�V���o�=:w�_|qt��% ��Գ���� �.��.��L�۷o��ٽ{w�+��wމK/�4���       �U ���oǤI�bݺu�l�-�믿>N:餸袋A��Գ܁je����1:K�,	�C����;�O�>�}-Z�h       ��ܹs㡇�+VP{��-3f̈Y�f�g�g�uVԫW/ rէ�f͚@.JGc=�����s�e��D�XK�h3z��8�쳣��        j�6�#�<ӧO��ڵkW<��S��k�e�܇yyy�kRϾ?p/..�+�I��NL�81��8Z�6̼���o|#:u�       5��ݻ��_�G}4JKK ���c���1mڴ����u@�9`�{ӦM �l޼9~�a;��
�|����/Ç�K.�$���      �&H�[?���v�� �,K�,ɺ�4���/�F�@.HM���=�s�3f̈��?��*�޽{��_��s��UW]ݻw      ��j�ƍ1q�Ę9sf |��M��iS�E]�	�����TXX��{�&M��mڴ)��~�� �,}�Q�����i�      @�TVVӦM�G}4JKK�pl۶-���x�����_�z�m�6 ������@UKS���غuk T�}��?�����ꫣs��      ��-[���K�.��1����Og�qF�{�Q�N� �
��ƍ@UرcG<���YX
P�֬Y�_}�5*�?��(((      �\�&�����^x!�P����<�L���;q�UWE׮]��	܁*�dɒ��{�� W�����ڼy��k��֭[      @�HS����?�-�
���o~�>|x\r�%QTT �E�T��>��s�裏f�� r��ŋ��?�y\|��q�)�      @UڱcG�ZL�6��v�¥Ǚ�_~9�̙�Ms/))	�ʰ?poذa T�u�������� �.�ѽ����~|�߈���       �l�g��~w�~�� �L�������iH�i�@E��7h�  *ڌ3���m۶@u���D�k��&�u�       �a׮]1eʔx��gMm�Lz�y饗��6��ַ�K�.PQ�)M@����c���P]�I7�pC�92��կFaaa       T�իWǸq�bŊ��4����7q��gǘ1c"??? �[Ve�׭[7 *¢E��������K;��N��=�}�;߉-Z      @yJ��|�W����;w@.)++��<�̙�\sM�j�* �S�7k֬(/// ���/�'N�ݻw@M�dɒ�����ճg�       (�7o�	&�{� �,���~�_~y:4 �K�7mڴ^ ��]�v�������j �T[�n�[n�%F�^xa�0      �ٳg����شiS T;v����ǬY����F�����@9ٰaC�q��tc��.��3���ի�ꫯv�      �4Hp���1mڴ�w� �͌3b���q�5�D�n��hd�{qqq� (��͋��+;.�6I;�����;����h׮]       ��+W�=�ܓ�Tg�ׯ�n�!F�_��W���0 �D��QTT$p�J�=����#�<eeeP�Y�&~��_�UW]      �����/�ĉc���P��l�ԩ�lٲ��w�M�4	��%p�ڎ;b	���o@mWZZw�}w̝;7.���(((      �OڵkW����+P-X� ~�ӟƷ���8��p�ܝ�?�0Ǝ�W�j����hذa�۲iӦ�z��W�ݘP��I��߳�ȍ7      �dÆq�wĒ%K�&ۼys�x�q�ęg� �*��֭k�;p�f͚�ƍ˦S}իW/5j4H�X���!�ԩ��~�����y��׏���O}Ϳ��o�q�ƀ�n����_�"��_�5�;�       j�y���]wݕE� �AYYYL�<9V�XW^ye�|�;pD�d�?��O�rS~~�����mڴ��m�F˖-�U�VѢE�,lO�zyK�!p�H�������k�_�~      �>��g�}6y��P+����jժ��w���K �'��������<[��w��%N<���ڵk���ѡC��رc6q����}���C:�"18f̘8��s      �=v��&L���~; j�4��g?�Y\}�Ն�k_�� _`׮]����>�z� w����N�=zD�n�8�gԨQU�gJ�;p�}��D�+��"
      ��>���;vl�^�:�Q�F�Ջ�?�8��J�~Ґ�ѣGǅ^yy�U�Ӳ�����#�6o���v[,^�8�z��q�}���^�zEQQQ��;\:Yaݺuّ[���      �fJ�� �t�35Gf��֫Wo�˩�(((�n�`�t[\\4�VӦM�y����������?P��!��<�L���k��O ���yyy�pk֬�[n�%��j�m�v�ްa��Uw�|s�΍_���q�u�E�f�      �Y���x衇����!��-Z��V��4i���"���p=M`?�
�?�f͊_���o��oѦM� �'�����	��gZ�pa�~��e˖�j���={������:Hxig�����l�V��_����}/ڷo      @�WVV'N�_|1�=�e8��G�1��شiSt��)[�s�Q��"�yyy6?�������W���~��ѽ{� HLpꭷ�ʎ�ڵkWP�:v�'�tR�x��qV�M�q�|�� n�ƍq�7ĵ�^�"      ����Ҹ�����rG�WRR�E�)d/((�ޞB����4>�����[��M7�W^ye:4 ���IO=�T<��v�V�t�U��~��'W�cw�ph�m�7�|s|�[ߊ���      P�lذ!n���X�bEP�RD������7�t�?j�i����{��l�~�w��j�� �'S�L��<�<͚5�dۋ���&H�;ph�Iw�uW\u�U�/})      ��c�ʕq�-�d�;U'???�v��{��&���=W��b�(c}��'cݺuYC������~`��ᡇ��>��۷�aÆeV5mס�OYYYL�0!v��#G�       �͙3'�����|T�&M�dQ��A����M|��_=>�����w��������V�{��ꫯ+���|:4;��r1�/m4z���c�F�      @�z�W���˚*W��|�	'Ā���lѢE �o�ܹ��_�:���h֬Y ����?5x���A�IGa��ib{�֭��KO,

bϞ=��?��ñy��袋      �-�wz�'O�g�}6�\�5ʢ���GqqqTW�¡Y�jU\��Y�~�1�P{ܡ�KS�Ǎ3g�*F�%|�'�i��V�vঠ�y����Gp��y����/�v�      ��JC���?�k��T�v��Ő!C����G��7nEEEQZZ��[�n]��W�����N�:P;ܡ۹sg�;6�̙��4��W�^1bĈ��GK��w8r)r߾}{\q�"w      �bi���~���1cFP�Rw���/}�KѦM��iRK��S_l۶mq�7������ҥK 5��j�����o��s��+E��k�ȑѬY���Z�j��~ G^�����oֈI      P�����w�y'�Xi�y������I�&QS���w8ti@�M7��^{m���#��M��P��v�-�ĢE���չs�5jT�m�6�Z;���믿;v��|�;QX��      T�4�j�ر�U���СCc���Q�^���R���x|뭷Ʒ����ׯ_ 5�B
j�H��Z�.]������g��:u
�O����w�}7ƍ�E�&�     @�H�����A�ٴ�!C�D�:u��04�L:Q㮻�o}�[1`�� j&�;�";w��v����O�ƍ���O�>}�D^^^p�t1����ݻ7��7s�̘0aB|����      l۶mq�M7Œ%K��W[��}Lp�#�gϞlH`�:lذ j�;�i��w�����^��JX#F���u�����(5j�6m
�|L�>=


��+��     @I����c�ʕA�*..�SN9%���7_KC���eee�����?�1��ӀR�f����I;���Θ={vptRLڻw�8�3���|���X����W_�z��ť�^      @�Z�~}�����5k��'<xp><�}gm���&M�Ć82{��|0�o��sN 5��j��Sm���1k֬�褝�g�}vt��%8t)p_�hQ �����&�@     ��v�ڸ��ȝ�N�0`@�1"6l���T���M�2%��P@�!p�,�P�����7��\�:ubذa���|4֑Jc@�Hh�1��3�      ��lܸ1��.n/?�;w���:+Z�n|Zj*�ϟ��KEj��cP�)5�{���W^	�\III|�+_Ɏ���ܡb���Ύ�;��S      82�7o�o�1����K�@�խ[���Z�h@�IE���8� �7�;�P�'O����/��iРA�=:����;T�tZ���ߟ]���&      �óm۶���c����ѩ_�~�92������T@�KCaӠ��ÇP}	ܡz����g�	�LϞ=����"w�^�F����(JKK�)r���{���E      ��ٱcG�t�M�lٲ�����E�>}�a�z�C'p�����/k(@�$p��W^�)S���q��q�9�D��݃�.b��ʕ+�8eee���.6l%%%      |�]�v�m��K�,	�\�6mb̘1ѡC�����I�i�P~RC1~��,rO�o��G�5��ٳ��g�4�=]l�O��cϞ=q�wď~��h׮]       �m�������͛��u��ȑ#cȐ!�����T�X�"���;�3��_�%kÀ�E�5ĪU�����v�q��.�Q�Fŀ��ӢE� *���۳)?�񏳓)      ��;�o�[pd:v��w�����w��63]w�uѭ[� ��;� 7n��o�9�9t�;w�.�@ Z	�nc��]�6n�����~��      ��޽{c���1cƌ���$x�I'E^^^p�4P�v�ܙ5������9@� p�jnǎ��6�&�5bĈ8��S]lUcP��.]�ƍ�k���q�      ���w�}��o����$ƌ�5
ʏ�*^j�� ����Ѷm� r����td�=��˗/M�&M��/��;.�<�8�ئ��@�5kVL�<9{�     ����'���_~98<���ѣGǀ��'p�ʱe˖��[�'?�I4n�8��&p�j���EM�=��΋������� �5k�֭�r=��s�&��#G      �Vo��V<��c��I/���h޼yP1�[C�r�v��[o����� w	ܡ�z���^�X���:�4hPPuҎc�;T�|0�G��}�      �6��Ϗ����޽{�CSXX_��cذa���T�Ե4m�4֯_@�[�ti�7.����ls	���P͘1#y�����d.��lG1U+�|�A �/��Ogir�N�      j��>�(���ؽ{wphZ�j_|q�i�&����C�5kVL�4)�ʀ�$p�jf���v��;fOB6lT�t1T��;w�رc�?��?���      P�mݺ5n���ؼysphҩ�cƌ��u��'5�������/ɾ�F�@��C5�.�Ү�]�v���:�����Ow�L�C�۸qc�v�m��(�ԩ      PS��"�nl͚5�KA�9�}��	*���ƃ>͛7�6� �E��DYYY�u�]�aÆ��
��s���#�#̀��lٲ���{�ꫯ      �������b��kӦM\z�ѢE��jܡj�&oܸq���?�?�� r����I�&9��4j�(.��h߾}�{�ի6�-[�P��O��:ur�      5��ɓ�7��X�޽�A�i�;U���:;wc�Ə�cߋ�C�P̜93������9昸��ˣI�&A�J;���1[�ڵ�N8!      ��x饗��g�>_~~~�v�i1|���5h� ���c۶mT��?�8n����я~�����	�!ǭZ�*Ə���g�ѣG\t�EQ�N� ���}ɒ%T�t���w���_�͚5      ��.\'N>_�F��K.�:�#M��C�I��]w������M@@��C۱cG�C���4�lC��3�<3������-�7o�;�3~��Fa���      T_i�n��מ={��k۶m|�k_�&M��%\�|y UgΜ9��c��\@�R2A�J������ի�OKA�駟j�U�V�ŋ��ɓ��K/      ��RԞ�ȝ��ٳgm֩S'�=�Bnx�駣}��1p�� ���r�SO=3g�>-MN\�z�
�����=�?�|t��%      P�L�81,X|�4Dpذa� ��2�IS�a�`�֭[G��w�A��~L�2%��z���W\��C5��8K;�w��@n�0aB�k�.;�      ���^{-^z�೥��_t�EѣG� �	�!w����;������P��c6n�w�}w���JO����8�c��)�OGj��� ����Ƹq��'?��#	     �V�X���ي���k_��!��D�f͢�� ���@�[�vm��]w�u���@��CIǛ�?>�n�(M��ꪫ�8��-�8�CnJ� 8iҤ��       ���b�ر�s���Ӛ7o_���u�H��S䞢Z 7�������O��g�@��Cy��b�ܹ��R�&��ȝ�ϑZ�ۦM�%%%ѯ_�      �\��s�=B��h߾}\~��ѠA��zIM��א[{��ԩS�x�T�;��˗ǣ�>�M�6��v]5��r߄	�c
�T      �5���={��c�>��:�Ï_��Җ����e�K�jX�l��j�؊�=��˼�8�E�v��$��E�U�UHt$$!�*zG4�����h�([���g�_$v{�9�>�뺃ˍ3&����:����򣩀ғ��~��_����0`@ �C�%���1~��_GSSS�aÆeq{�޽��p��w����p����,*++      J����c�����&L��=�XTUU婶�6��s�ԩ�������Gt�;����~:���|j������XܞC)pO/z---��>� ���C=      P
N�8��F���r�3fd��UTT���@(][�n�^x!}�� :���؆��^>5bĈ,n�իW�?ݺu��������(m�`���}-F�      ЕR���_�:Μ9\쮻�o~�A��Ci�7o^|��_�q��б�Ѕ��%&�/6l�0q{���J_�i!����?�yTWW      t����\�[��V�y�A>�^���� ������W��_��ѯ_� :���H��Kq�ɓ'��?��O����>� ��w���x����'�      �
�w��>�TEEE���1{�� _RS!p�ҕz�������}�w1�1��E/^��np^mmm���w��A��R�˒%K���.Ə      ЙΝ;���MMM�y)�|��b֬YA���f׮]��6d��}��@��Cؿ̝;78o��Y�ާO���P^ҭ#����㗿��A$      :��O?��:�y)n��c�̙A>i*�<<��s1f̘���hw�d)���~���AD߾}�?�i�ScP~�?�<�L��'?	      �iC�e˂�R�������Ӄ��T@yH7����g���kTWWо���,X۶m"z��?�яb���A����d[�Ϟ=@�X�bEL�6-���      :ҩS��7��M�H����o�����6��o߾x������}	ܡ<x0^x� �����1lذ��ҁL����C��̆�      �#��=��'O�λ����;��/-��֭[�(}/��r�(�_�j �G��$�~���Fccc]eee<���/})(�t���ݻ(/G���s�fCJ      �/^��npޜ9s����!u5)r?|�p ��m(����e�Ў��I��k�֭A��?�ƍ�m�����W_}5�M�f�     �vw���l��͚5+��ޠX��@�;��#G�ĳ�>?�яhw�Ǐ�?���A�]wݕE�P[[@yJ�ǿ��������      �������o���A������'�@yY�lYL�:��Wh'w�O=�T444D�}�k_���/ q��6g������|'      �=���+�u�� bԨQ��c�EEEEP<�B�ICZ��������ߢG���;t���z+֯_E7bĈx���������[�n���@y�7o^L�>=�      p#�9�?�|p����~�}�N1Y���ѣ��?�9����pc�A����?��Qt���GQ]]Ц��2�
�<��?�����       �-m���o~Qt�{��Xt��=(.�;��ŋǔ)S��n��	ܡ����ǏG��W�*���	�T:�	ܡ�mٲ%֬Y�g�      �˖-˾w*�^�z��C�ѳg��ӧO�>}:�򒆶~����/~�7q��:Ⱦ}�bɒ%Qdi�>C��ǐ�<�LL�81z��      p-N�<s�΍���������G��gA�����1����w����CHSXO=�T���D�}��_�������`�p�ԩx���_�     ���ӟ�gϞ�"Ky�5jT@��T�ܹ3��4o޼�>}z6,�k'p��v���_�5v��,p��#p��H���q�q��7      \��7�믿E7gΜ�4iR��4Pޚ����C��g?���k#p�vV__�=�\Ymmm<���>��B�0�~Nҭ@yK����K������      |��������7n\�s�=�J�P�Ғ�5k���ٳ�6whg/��R�8q"��{����OF�=�H�y�۷o�<y2��u��X�n]v�      |��W>|8�lذa�lp�|x�gb	QSS���C;:x�`,^�8����!C�\����!G��l�ĉ�       \ɡC�b�Qd�{���^��2`���֭[455P�N�:�?�|��?��	ܡ=�쳅~��1cFL�4)�Z���m۶�Ǐ�~��      �J���?�������}�{1p���ϒ6����f7����k��]w���rK WG��d˖-�~��(�#F����p�\�����/g����      \(�6l�"�ַ��F�
�"���C�kii���z*����9^����Akkk<��3QT麬'�x"�	�U�6򥡡!�^��?�q      @�����}ERWW�g���
ȏm۶�ڵkc֬Y|15*�����k׮(��~�n���ȧ+V�׿�����[      �ġC���R���#�\-M�˳�>�&M��={���p�������dq�Ѕ�կ_�쥭��>��H��<��s���      'N�����GQu��=�|���ѣG���C�|��G�g�c�=����Z�dI;v,�hРA&�iiJ}�޽��{ｗ=�ƍ      ����s444DQ}�;߉!C�\��STTTdƀ|X�hQ�}��ٟo�	��|��ǅ�.����'�x�d1�"M�!��Νcǎ�~�     @1�ٳ'V�^E5y��8qb��J]N߾}��ɓ�Cccc6�����|6�;܀ę3g�����7��\���k׮x��cʔ)     @1=��3���E4hРx���W��,p�|Y�vm�{�1r�� �L���ԩS�x��(��Çǜ9sڋ��-mq�4iRv�      �����{�ETUUO<�D���Wj*v��@~���������������rw�N/��R���G�t��-{���E��v������;�#      (�����瞋���7�7�|s���T@>m߾=֯_�'O�rw�ǎ�e˖E}�߈�C���t%[�hnn �^|�Ř9sf6(     @1�%H���"���g��Qwȯ46q�Ĩ���b
#���͋���(��n�)n���������Ƒ#Gȧ�G�ƪU����      �/u/��RQϞ=�G�����U[[@><x0֬Y�Ƀ+��5:~�x�\�2�&ȏ>��i1:L�8�C���/�e��     ��k��V��z��߿@{H?K������@����1c�-\�F���/���9s�Đ!C:�+� ��;�]Cy�]w      ������͋";vlL�81���� ���?G��e˖�7�� >%p�k��GŊ+�h�*F�ùR�!mq�={��c     �{�W��ɓQ4}��Gy$�����wȯ�R�q�ѣG� �S�5H$E��2;|UUUt����i�x͚5q�w      �������~���ݻw@{K�;�_i(l�ҥq���p���R�)����ӧ�M7���Ơ8�ϟ��~{6D     @����gϞ����׾�ƍ�����ۂ�{������ҢE�
��=]�u��t��={f?s�O� �:o��f6D     @~�����ŋ�hz��=�P@G�4�/5S���j|���@�W%��-[E��<I�1t�t �C1̛7/�M�     @>���gΜ��y����n�Q����jkkk ����/�׿�u[�!�pU�dTѮ��җ��Ǐ�L)p߹sg ��gϞx���]�     �iy`
܋�+_�JL�4)�#u��=���}�Q ������k�o}+�������
w}VUUU|��ߵU�N�J-(�����     rbɒ%���ޭ[�x��:Cj*�,ȶ���(2�;|�U�Vŉ'�HfΜ)4�K���bI�ӭ#G�      �Wccc�&w�}w���t��Tl۶-�|;y�d�\�2�瞀"���hmm-��Y555�t�;ϢE������     ��|��,�+���y���0�cΜ9QYYPTw��6m����G��{�ѳgπ�п��z�s��P�֭�����_80      (?---�[�<��ѭ���ci Ǒ#G�7ވ�3g��,�E;�6,�L��U***����@��_x�����c�      ����_�ÇG�����m��Й�P,/��r̘1#멠���<�mp/���ߵ&t�t �C������=z      �e�Q$UUUq�}�t��}�fߩ644�{�쉍7�����H��!moomm����W��F�
�j&��xΞ=k֬�9s�      �#�w�w�"����cРA�-mq����}��Pi���������n���Q���{�(w(�ŋ��w��j-     �2��IMMM�u�]]E�Ųe˖صkW|�K_
(�;\��U�
u�ϤI�bذa�@�Ŵ������E      (}�M�6E��s�=ѳgπ�����Y�ti���?(�;\���ˣ(�u����7JE�6������� ���W_�     ��E�EkkkE
��N�Е�P<k׮��<���P$w���͛u��̙3����"]0 �;@����[q�ĉ��       J�ٳgc͚5Q$�������*�+	ܡx���������w�D��HE�B��o�=�Ԥ-�w(����X�jU<���     @�Z�lY444DQ�9�MĔ��STVVFKKK ő��x ����B�8y�d����Q3f̈�}������|@���kq���g��     �����H�+**���P
�2�~��e7c�q�ԩX�n]̞=;�(�p�+Vd�c���vJY�8�)�ްiӦ?~|      Pz6l�G����4iR�1"�T��_���
(-�S$w�?����r��(�iӦe�P��a(�4p&p     (ME�ޞ��{��$5[�n�X�m��w�[n�%���ҋߡC�����;�(Uw(�w�y'�^�o߾     @�h���(,�i*���-[?���@���H�ۧL�� FI����޽{�ٳg(����x���m�      (1i{{KKK�偔���� �i�����ODϞ=�N�����!�|��(���*0�B�8���(��˗�     JHZRdy t=ܡ�R�v�ژ3gN@�	�����Q__E�`(uw(��{���ݻ�[n	      �������ɓQ�R����mo.J�\,-�Sw�_�V��"p ���8��'�|2      �zE��>y�d�)i�����0�xv��{�쉛o�9 ������c�֭Q'N����;�����������      �Ή'bӦMQiy�]w�P�RS!p��J}SOy&p��֮]���Q�g�(w�ԩS�y��7n\      �uV�^---Q�R�w��R����G�n`��O7���"=zt:4�\����KXSSS ŕ>��      ]+�tE�n���r`i ۙ3g��wߍ)S����Bۿ�ٳ'�`֬Y�$�� M<x0��z��7�?�aTWW      �o۶mq���(����flʁ�X�r���\�Shk֬�"H��o��r�dw(����l�x�ԩ     @�[�zu��픓A�e?�---ӆ�ԩSѷo߀<�Sh���zA�ޞ^j�ܘ8��y-p     �|���ٍ�E0v�X�QS6�u�-�<v�X Ŕ\֭[��sO@	�)�]�vő#G"�w��*ʖ�߀$M744D�=     �γq��8}�t���PN�@���--��Ww
뭷ފ"�<yr���3����s��e�<��     �s�]�6�ছn�[n�%����b˖-׶m���ѣ���Kw
��{EEE̘1#�\��X�9nmm���՗w     �Γn�}�w��㎀r#hRS���?��y#p����������(Wݻw�~���G}@����������     @�{���=��ƍ(7ii �����SHil̚5+�ܥ��������{/&N�      t�7�x#�`�̙QYYPn�@�gϞؿ>< O�R�2λt�J�����QUUP�ҁl۶m��[o	�     :A���K�O�<9����D�^���?��RO!p'o����ǳ���kii�g�y&���ƦM�(7&��6��n���FEEE      �q�y�hll������޽{���T�޽;�b{��7㡇
��;��~��,�+�ӧO����cŊ1jԨ,t7n��(w�ͩS�bǎ1z��      ��M�E0cƌ�rV[[+p��>���;����Q���oߞ=}���I�&e�����2�;p��9.p     �8is��"�7�tS@9�T m�pڷ��퀼�S(�Ν�-[�Dѥ���S.�@FϞ=���> R��裏      c�ƍ���y�������M>E��m�|�M�;���By���ȝ�.��>hР�:ujL�2%jjjJI:��ٳ' ҵZG�ͮ�     ������Q)ܴiS�����ٳc�������@��;wƉ'b��y p�P��W��رc�hѢX�dI�;6�Ꞷ�WTTt5�;p��5dΜ9     @�J���w1E�n_�n]��F"������
(i�e�ymnn���g��⮻�
��;��6����o:��'Eœ'O�6����;���8.�6i�     �ߎ;��ɓQ4)
ܾ}{����7&M�ӧO�������s�n�H������8t�P9r$�z�?���}�ҥ1f̘lRy�����Up��6o�---QYY      ���ݩS�b���bŊO���7�wS����R�$ipcccTWW�;�;����r}���>��B�4�<eʔ�޽{@gH�1�6gϞ��;w�     hg��Npޅ[�S�N�Z�����R����$���!�l�uuu�N�Na��$n��Çc޼y�x��?~|̘1#�Б�]���� I�\�     ���Ǐ�޽{��;v,-ZK�.�1c�d[�}WE�����6�6�;y p�ZZZ��$�O��Z�n]��1";�M�8��&t�����ȑ#�����      �ǆ���|����ظqc���ٓ'O�z�^�zt����&��7P���Ν;��ٳA�طo_�,\�0���5kV2$�=���h��������={      7nӦM��K�_���˖-����ǌ3bذa�m����&}>����N�N!l޼9�x)4�p�{
��!.m߆��Pssslݺ5��     �ƴ��h+�SCC�E�D��>q�Ĩ�����޽{[�	|"�͙3'��	�)�>� �\i��ܹs���mWr80�z	܁K��w�;     ������̙3��I�DzR+QWW�-2dH@GKME�s����{wʞ���KS�۶m���ӧc���bŊ5jT��7.*++�����6     ���6��~���?��~뭷f��رc���*�#܁����Y7�ѣ�	�ɽ��t����ؾ}{����7&M�3f̈���\�����v�ܙ]�أG�      ���M�t�ԭ��O�>1y��>}z0 �=���@��g�fM��ѣʕ���۲eKPZN�:�mu_�re�9�Vw�J
X�pD��H���cǎٶ      �Ϲs�eut�ӧOg�Ċ+bԨQZ	�U��p���]�N9��{|�AP��5(m[�S�N�)S�DMMM������P���     \���}SSS�9Z[[��;�;p�����
(Wwr-
�m���cǎŢE�bɒ%Y��&���rEEE@�t Kۚ�lݺ5      �~v��e���ѭ[7�*�'� UsssTUU�#�;�v���8s�LP>҇�ƍ�'�̓'OΦ�{��`���Ν;�A\�     p}҆W�֕Z�����+�j��KS�Z)����!>���lp
ʑ��\KSH��#G�d��K�.�1c�d��ѣG�%p.U__��n�)      �6i۳[�K˅�D]]]̞=;��ERS!p.����+�;����@�6�<bĈ,t�0aBt��=(�;p%i�M�     p�RW������J�_�>{�Z��'Fuuu�������>�������ʑ��\��Ͼ}��g��1~���1cF6,(�~��e��Ν�6�����      ��֭[����J,\�0��>k֬2dH��,.�>�[[[���"���ɭ4a�w�� �bݺu�cR�8��V�8޿ �1�     p}�m������OZ�[o�5�ǎUUUw�R�q�Y��ʍ���ڽ{wv]�gR�XҁL�\(���~�׳g�      ���ܹ3(O~�a����'&O�ӧO��%p�$-�S���֮]��b�pR9}(��}���&�sƁ�T�NkϞ=�|%      �:��S�N����ӱ|��X�bE�5*�M��ƍ���ʠX�B�4�~& ڤ���;�(7wr+mp���F��s�f[�Ӥr:�80(w�J���     ��m߾=ȏ�*�w��~���ԩScƌQSSGmm�����{ʕ���J�0�I���Wb�     �ڤ����ɓ'c�ҥ�lٲ;vl�J�f���"ȷ�T�ڵ+ ڤE�����-PN��RSSS�߿?�ͅ��}���I�&e������K�6N
---��`     ��ٹsg�o��ͱq���I���ɓ�ؽW�^A>Y\*us�3?<A9��K)nO�;\ɩS����+W���#G��ٳ��n3�\&�u��cǎ@�����w      �/��{��	��ȑ#�hѢl�{]]]�J><��;p%�f�;�FD.�޽;����m[�S�N�)S�DMMMP�ҁL�\����[n�%      �|�{���Ơx��j�ׯϞ#Fd�'L�ݻw�_mmm \JOI9��K{���)�n�T3fLv�5j���%*�[�l	��۷O�     p>��À��Zz.\�mu�5kV2$(_�n�N� m|�S���R�4��^�7nܘ=)��<yr����+(�����?     �ձɕ���Ǻu�'muO����㣪�*(/i��A��СC�&�����=z�(wr)M�:r��e[�G�t=�;p%>�     ����ϒ�s�;wn��=-�>}z0 (���jmm�={�ė���r!p'wҤщ'�˅[�Ӥr
�'L�ݻw�����     �X���|�ӧO����cŊ1jԨ��7n\TVV�MS\I���SN��N�$M�1���+=,Ȯ�1cF6,�\�{�Ξ�g�@�ÇGcccTWW      W�n3������پ}{����/�N���555Ai����K��PN���t�tS��u벧m��ĉE��h����k׮ h�~�v�����[     �+KK��z�<y2�.]˖-��c�f�D��^QQ�܁+�URn��N
۠3�mu_�pa���ŬY�bȐ!A�J2�;p)�;     ���q����c�ƍٓ���<yr����+�z鿓4t���1�F���;�
�
�
�����zk���媪����R��Ç      �M�N{:r�H,Z�(��>f̘�={��T]�G�ѧO�8u�T �9{�l|��Gѿ��r p'w�m��?�0{���S�L�&��ܸt�َ;b�޽�?\�{      �������>��>bĈ���0aBt��=�|i����TzаQ.��J�ZG�F)I���^{-�/_��v[v�K������;v,�y�x�������y��     ��RW�{W:ھ}��g�QWW�f͊!C��'��J7�;6��ɕt�FCCC@�iii�͛7gπb�ԩٓ���r�*�?�U�VŮ]��j	�     >�ѣGut����X�n]����)t?~|TUU���6 .�ʉ��\���rp�ĉX�xq����D\��>j�([��|ؾiӦX�dI9r$ ��ɓ'�_����3      �����B�<w��l���ɓc���ق@:F��p)K)'wrE�N9inn��7fO��M�{:����;�(f_z�ػwo ܈4 s��7      �U��N�>˗/��+W�m�ݖ��_��W,l'�q��yǎp)���;�r�ر�r���[�`A�ٽ��.��o���(�������իWGKKK ܨ�w��     �r�6JE�6oޜ=�:�)S�DMMMpm�����~l۶-8���p%��lll����R'p'W{�_�>{��M*O�81z��y��,?����0@{9~�x      p�C�����ޢE�bɒ%1nܸ��9rd��Μ9o��F֗襀��`R�5|���R'p'Wm����㥗^��_~9ƌ�f���V�49���OG}}} �'��     �2�)e��ͱaÆ�<xp�O�4)z�����G�k�����i�"��J�wʁ��\��G�@�q���馛���������u��e�~�r��	�     .׶��A
0�͛���J�H�VbĈQT�t��x��ׅ��1�F���+w�n�޽�3��� 7s��:th����z+^|���' ��      �������ƀrr�ܹx��7�'/K��{���_�ԩSp���;�q��٨��(�4�����'M(O�6-&N�X���?����v�C��     p9ߡP���Z�����~����^,�\�ɍ4iE�o߾�I��)S�d���A��Լ����v�S�w��wMEEE      p����h[
����92��>v�ب����H���ٴ�;���;�!p���-+V���+WƨQ��нTp{��^xA�t������Ě��      �<[ɛ� �ر#{�����R�D9���������<ڛ�ʅ���8u�T �p۷oϞt��<yr6��U�3g�ğ���,8�,'O��     \@�F��>}:�-[˗/�d)�q㢲�2�I���z�8w�\ t��Y��c�w�P���F
ـ��\:����]q�K��s�=��'��ҁl���     �yǎȻ��E���H��ӂ�R�u��ls{SSS t�4�6t�ЀR&p'7lp���U�%K�Ķm����     �؉'�$�̿��+�t��;vl�J��Qj����ӟ��@��S�䆐�N�.���v[̚5�Cp��6�t�      �ST��ͱq��쩭��N�:5z���������SOŹs��3|��G�N�Nn��צ��%6oޜ=�}�K��͛����     �������ѣ�hѢl���1c���G��?��x����:���r p'7Μ9��i�����cǎ�U�      |��ٳ����yMMM�lu1bD�IL�0!�w�ީ�>R��k׮ �L'O�(uwr#ƀs�n�С1}���8qb�����5���c�Е�      |ʦV�l���˞�:L�4)k%���w7o��V�
��潀r p'7�lо</��R����QWW�gώ�Ç�?o͚56']��?      γ��XZ藚���muOK������VCCC������ ��{�@�Nnܡc����ׯϞ/��+]i�v�� �j�      >eS+\����K�,�ɓ'g������_�ҥ�\]��?��;������ �`��?~|̜93������7ް�(	w     �O�>}:�k���,_�<V�X�F��B�q��Eee�u�k>|��@�K	�)wrA��+]��nݺ�i��^WW�W��R��      �S���imm��۷gO߾}cҤI1cƌ�߿�5�k��/���� �*�
ʁ��\����k�mu�?�������      ����O�|����Z�*ƎӧO��#GFEE��s�n�;v�����������m����¹s��Z�v��455e[��H      ygS+����}�ƍ�S[[S�L��S�F�޽?�bŊ �j��H�o555�J�N.����X��޽{      ��б�=�-��K�Ƙ1cbڴi1z���w���g{;P2����R&p'� ������      �̙3t�t�t�V��Ç����c	���+W��R�vJ���\� ��~      p�������/��B,\�0���bӦMP*�P��䂀 �Tccc      ���@ר���u��@)�n@���w �R�      ��	 p!��:�;����  ��     �< p!��:�;����  jmm      Dl �żP��䂀 �Tsss      ��[ �bwJ���\�� ���     ����&ߛ  �S��䂃 p)�      6 �rnw��	�� p)�      �3 .���P���� p)�      �3 .���P���BEEE  \��     �� ���:�;�PYY  �~      `C+ p9p�:�;� ` .��      ��V �rwJ���\� ����
     ��� ��~@���w �R       ��Z[[J���\� ���     @S \���N�N.� �K9�     �� ����R'p'�u� \�{��     Pt6 �R�(u�`rA� \��     �� ���J���\� ����     ��� ��~@���w �R�      l �媪�J���\� ��~      ѭ�< ����R��\� J�H�      "��� �B�KJ���\�ѣG  ��ٳg      p~1P�����  ���R'p'z��  m�      |*Elw ����R'p'��4q���  w     �O����ٳ ��)uwr���"z��gΜ	  �;     ��Dl �����J����H!�� H��      �	��y7��	���Z�6�      >e9 p!]�N�Nn8� m�      |J� \HWA���}�� ��_�~     �y"6 �B��(uwrC� �1�     �) p!��:�;�!d �|     ��� hӭ[��޽{@)��B6 ���7     �O���+  ���;�!d �|     �TMMM  $nv���! ЦO�>     �y�
 �M���J�����. ��I����      ༾}� @⽀r p'7R�^YY--- נA�     �O�� ��^@9��)nO����� (.�;     ��Ҧ֊��hmm ��lp��ɕ�
����      ����޽{Ǚ3g (6�)wr%m۷o ����      K1�� ���r p'Wm ��     ��0 ��� @��*(wr�_� ��     ��� ����y��u�����0�0�30ð�"��b�7�D��W�TJ��m;��{�U7�][��ʹ�̫�l�i'��Ina*����2��,2���t��PYf�.��9�3�R�����|>���xO@>�SP (n���     �_�իW  ŭ[�nQSS���A ����l{M      ��i� @z?PRR����������  �O�{      ��� ���B�NAi�ںq��  ���\      vM� x?@��Sp���#p�"%p     �5[ ��w
N
����? P|�      �VYY555�y��  ����|!p��� (NMMM     ����B� �K_I��Sp��� @q�>      �ͥ���V�
 �8	��w
�� �SUUU���      ��w �8UTTDMMM@>�Spz�oݺ5 ��a�     �[3� �WZ�VRR����ܷo�xꩧ (���      ޜ� ���\�'w
R��*p��b�;     �[K������  ����|"p� ��
 �ǅ     �[�������ظqc  �EWA>�S���� (.��      o/�@�18�|"p� 4( ��&����      o-Mo}�� (�������/�����,tkii	 ��80      x{)p �KCCC�����;+Mq�@q�     ��; ������;+�n<�@  �O�     �{R�VRR��� �;�F�N��@�H;�      ��z����/ P����;k��� �����ݻw      �{R�&p��ap �F�N��իW���EKKK  �k�С�6�      ���w�} ���J��;w
Z
�V�X @�J�{      v�)� P<�y��@����&p��'p     �3w (�7w
�� 
[Za�|     �gjjj���.ZZZ (lw����6dȐ(--��;w Px���UUU     ��IM��~��  
����#�;�{��1`��X�fM  ��E     ��I�Y� P��������|#p���9R� *��     �sÆ ���m%%%�F�N�K��w� @�5jT      ������s��  
S
�!	�)x)pO+�Z[[ (������      칊���߿�]�6 ��d�����WSS}���u�� P8Lo     �7i��� 
S<dȐ�|$p�(�)�w (,��     ��1bD�� ��������H�NQH^�_ P8�      ��� (\���|%p�(�3&�n���5 ��WWW��4     `����;;^|��  
��l�3�;Ea�������X�fM  �o�ر     ��K�� 
���|&p�h�)�w (w     �����˗ P8���uuu�J�N�H!��� @~+))�ѣG      ��tW (<���;�;EcĈQ^^۷o  577GMMM      ���	�--- ����? �	�))nO��ʕ+ �_iW      �Ϙ1c�W��U  ����$F��������� ϥ�9      �G� �c��ѳgπ|&p��p�q�7 ��z��Ç      �O�A7M{mmm  ���k�������hjj��> ��������      ��&���v��  ���B p��L�81~� �&L�      ��4�]� ����<F������	� ����f�     h)p���� �_#F���ݻ�;�;E'�N����-[� �?����     @�5jT���#^}��  �S �@�N�i����_�: ��1q��      �c���Ř1c���  ?	�)w���,p�<���      t��	� ?���/���P��q��EEEElݺ5 ��7hРhhh      :N
�KJJ���5 ��bz;�D�NQ�޽{�[u ���v     ��WSSC��'�x" ��"p���)Z)��@~8蠃     ��7q�D�; 䙪��>|x@��S��Yyyyl߾= ��5`���۷o      �����[n�% ��q�DYYY@��S�***bܸq���. �ܕn�     �9����_�~�nݺ  򃶂B#p��r�!w �qS�L	      :O��~�� ��*++c̘1�D�NQK�r���#^}��  r�СC�O�>     @��@��0aB����;E-����}��� 䞴�
      ����9B�~��  r[Z��F�Nћ2e�� rPIIIL�4)      �|tP�v�m ��ݻǸq�
����7f̘����M�6 �;F�uuu     @�K;�
� �p�QQQPh�������?�i  �c�ԩ     @�8p`���?�}��  rӔ)S
����a�&p��V|��     @�I���� �{���b�ر�H��k��1hРx�� �z�'O��     @KSao���hmm  ����[70��o6���ӧ� G��U      �Z1t��x�' �-i�(Tw�?i����Ŏ; �:MMM1lذ      �륞B� ����>F�P������������ t���JIII      ����3m�4mM�o0c��; t�����"     �ܐN�81��  r���B'p�7=zt455���? @�;�����.      �i^�; 䆑#GF߾}
��� m�q���M7� @�{�;�      �q��E}}}lܸ1 ����A����8����[o��۷ �yc���      rKiiiL�2%n��  �NEEE|���N����:&M�˗/ ����i7      rOx��Gkkk  ]c���QYYP��)��@�)//��     @kjj�Q�F����  ��GP�Æ�!C���ի �xiK˴�
      �+Euw ����Y��@�o��|g|��_ ���.      ������hii	 �s͜93�X��ML�<9n��fe ��ƌ��2      ���������G?�Q  ����29䐀b!p�7�.���Z��zk  ��v     ���Z���Ǳs��  :ǴiӲ�����B�(�����ؾ}{  �O�>1a       ?���g�w���  :Gj����-���Ĕ)S⮻�
 �����%%%     @�H�x� �9ƌ(&wx�gώ��;Z[[ h?���1}��       ��=:���c�ڵ t�#�<2����m455Ł+V� �������       ��)��^{m  �O�>1~���b#p�����w hG)l�9sf      ���N���rKlڴ) ��������;�!C�ĨQ���G `�͘1#���     ��ԭ[�����  �_UUUz��H��)Mq���+++�V     ��Ҏ���~{l߾= ����UTT#�;즱c����c͚5 콴]e�^�     ��V[[�M���/~ @�I;�H1��n*))��s��W���  �Niii�+
      �a���q�w�Ν; hӧO��={+�;�<0���c�ڵ �iӦESSS      P����{�7 �}��}���L�{ Mq�7o�)� �Lo     (L�z׻ⷿ�m��� �o�±>}�3�;�!S�`�L�2��v     ��:�ѣG�ʕ+ �7�sL@���JS��ΝW\qE  �'Mo�3gN      P��=�X�; �������������A�5k� ���M�fz;     @>|x�5*}��  ����'w�i������K_�R  o�[�n��'      �4��s��\  {nܸqق1@�{-mb�1 ��#�8"     �:
- ����/���K.�$ �]����w��]     @qH;�
�`ό;6F����a��@&L�>�`  ��#�����      �8�=:F��=�X  �g޼y����Q����CEkkk  Q]]�sL      P\�?����K x{'N̆�!p�}����zh�}�� �EZ]ܣG�      ���Ho	��� ��JJJ���~w M���㎋�����u��  "�#�      �S����CEkkk  �v�!�����kwhuuuq��G�~��  "N<�����[M     �b5`���<yr��7�	 ��ű���SA;�={v�u�]�q�� �b6jԨ8��     ��6��X�bE�ر# ��v�a�E�>}�{wh'ݻw�VS]{� Ū��$.\      ����~x���? �/***b�ܹ���ѡ��]�=��� �(�      �̛7/��x��W ��c�9&����5�;�����X�hQ\r�%��� PL*++�m&     �MMMM��]o�9 ������>:�7'p�v6lذ�:uj,_�< �����={      �ёG���/�^ (vix`EEE oN�`��q����^��ѯ_��9sf      ���֭[w�qq�UW ��ƴi�xkw� ���1gΜ�馛 ��I'�eee      �2y����OO>�d @�:�����$��&p���׺��cݺu �,݌;vl      ��I1ߢE��3��L��� �I�&�������CISl/^����\�P�*++���      �vӧO���+ �����ǂ�=w�@#G�ta@A;��㣮�.      `w��K+V��-[� �9s�D�޽�=w�`i��<�7o ($C��#�8"      `w���ļy����n @1hhh���>:��'p�V]].����: �P���Ʃ���}     �=1k֬���c�ڵ ���O���� v��:�ԩS�W��U<��# �ਣ���      �4DiѢEq饗Fkkk @�?~|L�81�=#p�NPRR��vZ�˿�Klݺ5  ����Ҷ�      ��F��vX�y� ��{��ق.`�	ܡ����;�ϟ7�pC @�J���8㌨��      �'�pB����y�� �Bs�q�eC�='p�N4k֬����� �G3gΌ�#G      ����X�pa\}�� ����9���#p�N���.Y�$>��O���� �I�n$      �^�M�˗/��+W ��	.^�8����;w�dMMM��w�;n�� �|�v�UYY      О���d��m� �����aÆ�����:�x���� �3f̈q��      ��>}��q�7�xc @>�ݻw̟??�}#p�.PZZg�}v���klٲ%  �544Ă      :ʑG+V���<  ���Ē%K���"�}#p�.R__��̮�� �\ն(���2      ���(��N�O~�}�� �|3cƌ3fL �N�]�����S��=�� ���̙Æ      �hMMM1o޼����� �|RWW�| �C�]lѢE�jժذaC @.4hP�     @g9�cbŊ�z�� �|�v!Y�dITUU�>���z��g�uV\z饱s�� �\PQQK�.����      ��RZZ�=������k�� ��f̘�Ǐ���!><�����   �r�)��      ��c��o}+  �544Ăh_w�s�΍������O t�I�&����      �J����#�Ľ�� ��Ү#g�}vTVVо�#�Nv���'m�@�I+��,Y      ��/^�V���7 �9s�İa�hw�!)*<���k�	 �lm��z��      �ժ�����O�/|���� �+��@��C��>}z���=�� Й�?�x+�     �)cƌ���:*~� 䂊��l�`YYY C�9hɒ%�nݺx�� :�ĉ�裏      �5���φ�Y�& ����=�� :��rPyyy��}�O}�S��+� t�޽{�g�%%%      ��[�n٤�O�ӱm۶ ��2y��6mZ K�9*ņ�sN|�_��;w t��EU���      ��_�~�`������ �cɒ%t<�;�1c�Ĝ9s�?�A @G8�SbРA      ���xG<����� t���HX[YY@��C��7o^<��S��� ���;,?��      �|PRRg�yf|�ӟ�^x! ���x�1x�� :��r\�8;묳�3��L�_�> �=6,���      䓪��x������gc۶m m���1s�� :����/ζn� �/jkk��s�Ͷ�     �|�����zj|��_ �HMMM�dɒ :��	�Ā��UW] ����ʲ����>       _M�:5�x���� �***������t.�;�C9$�8��; �ƢE�b�ȑ      ���O�5k�ĪU� ���ŋ���t>�;䙅Ƴ�>�<�H ���5kV̘1#      �t��-����O}*ZZZ ��QG��t�;䙲��8��ⳟ�l���7n\�t�I      ����6�=�������رcG ��=zt,X� ��#p�<TYY\pA�ۿ�[l޼9 ����/�9�(--      (4Ç�N8!���� �޽{�ҥK5���m�.��2+�xS��_�(�G�      ���#��5k�į~�� ��Q^^�}�{���&��%p�<6bĈX�xq\s�5 +]x-[�,      
ݢE���}�ڵ {���$N?��<xp ]O�yn�����K/����� �6��묳Ί�C�      ����x������g���% `w͛7/9� r��
@:�n޼9~�� $'�tR|��      Ť��.�?�����Kc۶m ogҤI1w�� r��
��'�7n���? (n�gώw��      �h���q�gƕW^��� ofȐ!q�gDIII �C����4�.]�]vY<��@qJ�e��      �,�v|��ƭ�� �+�{��.� �w�@n�CI'ڴ�ֿ������? �1c�XU      �gΜ9�~��X�|y �UUUŲeˢ��6��#p�SSS����K/�6 �aذaq�y�E�n��     @�C�v�i�y��x�� ��V���������PP����㢋.�"���� ��80����GEEE       QVV�{n|�s����~: (nm��F�@��C�jll�}�CY�iӦ �0555�>��l�,      ��UVVf��.��X�~} P�.\S�N �	ܡ�����/�V!oٲ% (,}��/�8jkk      xs555ٮ�)r߼ys P|fΜGuT �O����9�@���?[�n 
C}}}\t�Eѳg�       �^ �lٲ�����^ �G��~�)���P��~\~��}��  ���)n�ݻw       �oȐ!�| ���/P$<��8�3���$�� p�"1z��,r��;v� �SUUU\x�ѷo�       ���������j( 
ۘ1c�sΉ��� ����رcc�ҥq�W�Ν;��RYY�Mn8p`       {�-x��+4 �mAS�nRY�7��B�9蠃���O�k���@Iq{�*q���      �<0�8㌸�ꫣ��5 (C��:���� ���дiӲUi_������_ r[UUU����aÆ      �~�N����^{���@477g�E&�'�;�ɓ'g'�~���}��  7����E]�]|      �o�����k��7� �>}�ą^����/�;����g۰|��_�.� �-={�������      �q���wƖ-[����~ ��z��u����7�;�Q�F�?��������J �z�>766   �-�رc��}�{���  @~�7o^l߾=~�� ����..��⬷ ���!C�d+׾��/��/� t��}�f�����  @�Ν;�)z)"O1y�ұu���{���j�1}���g?���?���f?�>�}�~����+�L:v���RRR��<�����]}��������O����ʲ�����\^^���+**������ا寧m�Zڞ9}���
   �����]��v�m@~HQ{�,(w 3hР�������?---@�8p`\x�QSS   �b۶m�y��?��)VOQz:R�����������):o;
͞��)�o���t�ħ�-�O1|����6��G�QYY�}La|:z�����  ���p�	����o�9 �m)j��?(n���3�g������q�e�ņ�Εv���>��,  �Ui�?��Y���+�d��H�-To��S��>���s���.$H�wW����I��c[���t��b����/�ӑ�  ��fϞ�����|ǵ-@�J�[��^WW@a�%�d��⋳�}���@�5jT\p���  �Ζ"��7f��7mڔ}�"�4a�m��`�]i�}H��ۤߛ��65>M�O�H���t�§k����,�����~  �+̜93[�{�u׹�1��/�0���;�wz��Mr����㩧�
 :�Ag�}v�0  �=�����HS�����i�)H��UڦƧ�����V�b�tݜ�����)�Oӹ��� ��2cƌ��ꫯ���F�˖-�& �I��Rz8�&����g���@ǘ5kV�|����  `w�M]O�_z�l�z�����q�6�7���w<���J���"�4>�'555ّ�u655Euuu   �C9$�ָ��+�]� �:�F��.���(pw�M������}q�-��m�� ���ϝ;7�=��   �[)�}��c���Y̛&��p�m�q���ߋt��'iǂ�������S߽{���g������eccc���  ���8qb�w�y�|E��E&L��}�{�!@a�o)m�{�	'dx����lR ��[�nq��ǔ)S  (^)T߰aC��	�i{[��A9�����?�n�����#�<��_�L������uuuY ��ܜ��  @q7n\\x�q��g�� t�ɓ'�Yg��ݿ
���-3f�Ȧ]u�U�m۶ `龜�iw��e  P�^~��l
{���D��y
kS��	���o����Y����{���o߾��  ��0r�ȸ袋�K_�R�� ����ŋg�Z�� pv���G���i� {&톱lٲ��7  P8R��nݺ,do�طnݚM��C�x��==\M�{eee���D}}}455e���  Px���ǲ���� :��ٳ��㏏��� ����#i+ޏ~���E�ڵk��3|��8���  @~j�ƞ\��5}�B���-�Ȑ��#-tI�N|���{m����o�l�{�>}b���Y  �4�*	��W��=�X о�@�E��G@��{,=����?W^ye<����[�>}z�UV�n�z @>x�����"���]
ٷmۖ� {ꍓ�7l��?�x�}���C�4ݽ��*jkk��}����W   ?TWW�E]���7�7��M �>***b�ҥ1q�� ���
�+i�������w◿�e ��҃�M�1�  @nI�z�ľnݺ,dO�_}��,d��u(E��H�C�W�ξ��'���)|�ٳg444D������>  �ܓ�\�}���{��o�= �7i�\C�	�x	܁��.�N=��l;���ر# ��4�!�&;vl   ]+E�)f_�vm����iӦؾ}{���@�I�{Zp�����O<��雷��!occc6�}РAv� �PRR,��}��u�]�����K���-[�{�����	�3fdo.��կf��]�q�v�hjj
  �s������3�ĳ�>�MD~�W���bv��;6lȎ�+Wf_K�{Zh��E�E�555  t��;,z���i�& v_ x��F�=@����Ç�'>��"��'��b5q��l����   :N�p�~��x����---ٴ��u�b�v������W��_���QZZ�ݛ�������)~O_  :֘1c������/����Ҁ�E�EYYY $w�ݤ�%_|q|��ߎ��+ �Iz@<��8�c�- ���&�=��ӱnݺظqc6�=M1`��b�-[�dG��"I�+***���6��{���!z ����k�E�k׮ v-ݗ8餓b֬Y�Fw�]����i���F��믿>�n� �.m�����i  ��IQ�3�<�=�}�bӦM�}��hmm �^zM�ґv�X�re��{�)zoll�"��  �������h|�[ߊ�˗ ���:�9���Kw�CL�6-W\qE6]�P�92���ٳg   {��_�5k����?---ٴa1;@�H��iG�6dG�������l�Φ��>|x��  �siA�g�����[n�%[�@Dsss�w�y��� �"p:L�~�������7��{��B�&��-�.\eee  �������g��B�W^yŃ]��^���u:����+�{��_6�2�9C���ݻ  ���s�ٳgg1�UW]���(f�'O��N;-***��܁�&����&L�뮻.����Բ�O?={m  v-��<�L�]�6�ξiӦx���Mg�C�����cv�^�:����֭[���fS��i�;  �k�ƍˆ~�+_�u��@�I��ϟ�sL���܁N1mڴ<xp|�k_�n�ѣGǙg��m�  �EKKK�Z�*���H��
ێ;⥗^ʎ�+Wf�{��My4hP6̔w  �i��'>�����w�uW �4H�Ί�c������_�~�},n����; ����s�̉y��YI  ���_�'�x"�8����۷{�P��[�lɎ��i���Q^^�MyO������a6  ��>���N�Q�Fŷ����
@!9rd,]�� A`�܁N�.�N>��1bDv��v ����8��c�С  ��瞋'�|2��&����� o%�:iAT:~��(++�"�4�r����=  (VӦM�����W\6l�B��̚5+.\�� �w�KL�4)[�w�5��C= �*�XZ�hQTVV  ��;w��ի㩧��^x!^~��l2/ �tٱcGlܸ1;y��Awuuu���7���=i=  (������o|#x�� (UUUq�g� {C�t��5�e���;�o�1�n� �"M[�d��-  ��k�����O?�t6e7�&h���sMZD���gG
�{���{�����l�{�ne P�Ң���??k'n��l'$�|6t��X�ti444��rW�R�Ō3bĈq��Wg��ڸq����O��={  �m۶ţ�>�]����K�� ��R�Y�c͚5�|��lW����6lX6�҄w  
Q[;�y~�k_�g�}6 �Mz-�5kV,\�0���`_܁�Я_���G>?�я��?�q�U-@gK[d�x�1}��  �B�s��X�zu�Z�*^x�x��W r]
��9+�0����<M��۷o�92���  
I������x�|��q�w@�������>;�^hw g��{�{lL�4)�����;@g?~|�z��E  ��{.{�X�n]����Y$ �,���9���ώ4�}����>}�Ę1c�w��  ����<N>��l����_���J ��z-^�8[��^�@�I+��4����gq�-��&�Pij�	'��m�  ����%�׮]��9Mm�B��u�6mʎ��gϞ1`��;vlv�  ���ɓcԨQq��ƃ> ����2.\�� :���I�AđG�=���7��m����M�SN9%jjj  ��k����|O=�T��⋱}�� �b����7f�C=�M�L��<8�"�{��  ����6.������;��o��[�@.H�L�y���� A��~��Ň?���{�������v����-����  �;vd�W�^��h�[K��֯_���{o6ѽO�>1bĈl�;  䃒��l:rZ�y��Wg�� �JZL>��lpiz}�(w �7CӦM˦��t�M�|�� �iw��3gf[  ����%��Ӕ�M�6Ekkk  {.�C� �'�|2;��ʲi�)tOCҶ�  �������G�g?�Y|�{�3� �tÆ��N;-X
���@�H��6ӧO�뮻.��� �]��SO=5ے  r�Ν;�)\�V�ʮ{�m�&j�����ƍ�㡇���7���  �4�+MM�8qb\{��裏@GKSۏ=��8�裳�!�� p���������w�qG���?�*xK���1w�ܘ5k�-  r�k��+W�����	����q:�#�C����&Ӎ92�w�  �KҢ�}�Cq�wƍ7ި� :̈#���MMMЙ�@^J+gϞS�L�[n�%�/_ o�Dv�a1���o��  r�s�=�E��֭�W_}5 �ܑvTy�����{�=zD���c�رѫW�  �\PRR3f̈ѣG���_������TUUł��"�� t6�;����3�<3=�и���g��Q���;}������Ir��@¾( ⾡�(�-ڷ��u{z��{k��<�5U��>������wf����]^���Kk7����l�����dO���"\�n[� Y^/�S�sN�]b��������]���/bٲe  S���H�2��ѣq� `�K;���Ç�TTT��ʕ+�;�c   7]js������O���������C<��C���Q__ 7��;0#������x�w�W^�7��g������<_l �ͦ� f����hooϓ������˗�]wݕ��  �f���{c͚5���/��o��k|)s�w�w��fpf�Ԝ�e˖x����^�m۶��̗n��_�U���?����  ����ɓq���8w�\ 0s��Pooo�۷/O�X�%K��}�ݗw �-�7M;]�_�>������� �&�,�y�x��d.�)C��q�[jp~����׿�u�޽��d���Л6m������5  7���D?~<:�C�Z��522��Z[[s!KKKKn�[�ti  ���z���?���Ď;b�֭��� �w���?��X�hQ L%����`���������/⥗^�#G�03���Ń>���.  ��R�=]k<x0:::,� �&������ӧ�{SSS�~��  7B���aÆ��{����w�ɟk$)W������{�7 �"w`ƻ��������y���q�ĉ ���z����+W�  �QR#�}������^�v ���^��������X�vm��:�P  �S]]]����a�_��q��� f����x��b˖-yA6�T�;0k�P���_�+v��������`����[�g?�Y�[�.  �FH[7��q������ �*5fvvv�����>����X�jU�y�Q,  ��T �?����O>�$����3!0{�]}�������FCCC Lu����N�z衸�����W_}�ELq��rK������y  p�uww��Z[[��ŋ p��a��0�q�ݻ77k.[�,o_[[  p=��ʹ���wߍ������ f�T
���ݿ�ל Ӆ�;0+�����?7n�?�0^y���0Ť��-փ>��  ��r�,;u�T��� �����i�����s�=5�����  L����x���G�!���{/����Y�,Y���w�uW L7������6l�[��޽;~��Ĺs��y�/_?��O� �������>�� L9)��O>���<W��iS� ��T__���>�l�������>&&&�ޚ��r��M��P(�t$�P�B�=�PԦ�������8�W�������7�  �zHA�O>�D� �V�¼49�~��w��M  ����������ǹ�=�����2gΜ�`%��\YY әO� �"�S�6��Ç㷿�m? �G�o.m��V�z�  �mdd$���G����^7� �i-��|��Ǳw��ܶy���wܡ� �I�dɒ������Yگ��8t�P S_]]]<��39�^UU 3��;�7X�fM��G��믿�oB��H+�7nܘ/�,X  0�FGGs�i����  3M��:��?����裏���1֮]��v��;  ?X�}��������lꩧ�駟���� �I��E����������.�{ｼ%,�ݥ-�7oޜ/���X  0Y&&&�/�����7���"�uvv����cǎ9�~��w�1 ��J1`*�x���a�lfw�k4������=�\n�y��7��ٳ|��˗Ǐ~��ذaCno ����P{
u��  �ٕ������������sO,^�8  ��J�������Y�?��?������R�`
�?��Q]] 3��;�w�N�x�x��������o�>��GR�������  L����ػwo���� |����8}�t��Y݊+���"  ��m������?�{�7b�Ν>�� �r���?�y�b� ���;��TVV��w_����x��r+N___�l�Z����{,���  &C�ٳ'Z[[cxx8  �v���q�ȑ<i��U�V����n ��-[�,���/���ױm۶��H���J��=��3��#�D�P��ħV �`޼y���?�i\���C�iug�H7��b��Zxݺuy  �P��)mw|������u� 0	��>�;��϶��޸��[  ���*��_�"g%R!�R@��R�⮻�-[��w� ���;�$J!߇~8OWWWގ�w��]ttt�D�/��7jk `R�<y2>��hoo��1 �u��ϱS����}��ʡw  �.���ڵ+�x�hkk�ڥ������'?�I,Y�$ f;w�뤱�1�t>��q�������w�-�^]]]��jӦM�|��  ����ߟw�jmm����  ��ˋ�TWWǚ5kr�{�X  �V)��aÆ<iWƷ�z+>��S%�455œO>�?�x�c p��;�u��Z�n]�����sn!����������Aeee��*}q�}��&  ����F_|񅭋 ���������yZjsO�m�~��  �ŕ�Dwww�ر#�~���/Y�'�x"x��(
��I��@)$��xM��}�Q�ܹ3�=�����$������֞ښ���  &CjM�ϝ;�Z `�J�i)��}�����c��9x���  p�Ңɟ��'��3�䅔��=���\�٨��!6n��7o���� �L��&����[�I7	҅\
x���Y���S������O `2����ȷ��-��� ��#���>}:OMMM�^�:�X,  �Ej�N�i�����C^L�>7��,�ݿ����������o'�0466�m��������w
�sݥ�P�b���{�'���  &Kڱj�޽q�  `��E-����m�i��e˖  \��;��~���������������H�L�p��x��cӦM��� |7� SLڎ(mE�fxx8��S�{
���;L����JS{
�WUU  L����سgO�kk ��.]��w'}��7���2V�\�<�Vw  �YYYY�q�y����s��������|��9s������Q��
��O�`
K��+[t����]9r$>���܎s�ԩ�k������[sC{�J  \�� f����8|�p�[�;  �G]]]<��Sy�B��螚�O�80���)׳aÆ\4XQ!�	0|7�&R@���n����<����СC�����{�����?����ijkk  &��v  ��� �dhll���~:O[[[�ڵ+>��hoo�
�5�]wݕ��w�}�y �w�i���>�(�I7R���r�=5�\�x1�]�E�ڵk�"��*���9  �z�� �_�ǭ�>�`,_�<  �H;����~�O��A���}kkk����r��ӹ������: �~�f�����u[�l�x��/��{{{��%5�_	��cz  ד�v  ��+��۶m�� ��dɒ<���Ν�ݻw�'�|ǎ��0��{��-�h0]� pc��@_�?��S�����8q�D��I�S��CUUU���n��I�v�  �(�� �_muoii�͇.  ���y�O��<i����}
����/^��{o�իW� 7��;�,���M�N��t#!��Ӷ]'O�̏Ϝ9����͕��R�=mכ��[oͫ��B  �����w�ؑ�\'  0�R�f{{{���Q]]�=x��� �����œi�g�i��������?����_2gΜX�n]nh�뮻r���O�`�J�&���i��ӧO��4)�����/��mjjʫ�.]���)؞V��� �͒�v��n�  p�ŧ�~�}�Y��tÆ���  �}����r����/����{
�wuu�[EEE�Y�&��<+V���0	�pU:�O'�i�*m�B.W�Y������٩����i��4�-ʓ��͚���  ��mbb"��I��t�  7ZZ\�>~��s�}����Y5  |W�������I����ȑ#9�~��ᜃ`f+��p�J�=S���M��o���J[Ħ���I!�+��4.\������3+�
�EUccc477�c
�/X� �׬� `*Ja��;w������=  LiWѷ�z��N��<�]/ ����C=�'I��ʡ��G�ƩS�|V:ͥ���zk�Z�*�\V�\��^|��{K7�4��9ccc9�~%����J�nN\y�&�j�T>���������;�ܹscΜ9W�ijj�Gv  ��Ԍ�k׮���ٰ( ��itt48�;bnذ!�U  `���G}4O2<<���q�رxO� )��Ԕ�멝=گ���ϟ L� \7�B"5���9�~�&�䇆�b||���tA��U��k�&կ���ɍ�W�UUUy;������+�^ ��$�?�ݻ7o��έ `�H�2�"�_|1�ׯ_+V�  �l)+�v��<W�C:M��'N��ٳg���`)ױt���Ⱦdɒ���[n��0C����q%\~��x  �ۥ�v�ܙ��l� �t�v}뭷���2V�^�<�Hޑ  ���cX�fM�+R1ߙ3gr���Ǵý�����-�b�r�%�]�   f�tCe׮]����
  3���h8p <��.6l���  p#������R�=���?>O{{�������ei���������㦦�(++ f7w   �"5��޽;}ҍ  ���bδ���_�y��Ń>+V�  �R�}�ʕy�XZ��
I�����4�q
��݊Ҏ��]
�ϙ3'�9z:���tL��t�;wn �_"�   0ͥ#��=�W���  �F)��[oE�X�;�3���(
  SA
~�݇�|���n___�������ϡ����̏�1=ʏ��I�'###1666)������\���:�s��~z�����D]]]>���_�\O� ~(w   �i*x>����X��+ �����?�8>��X�fM�_�>**� `�+//ϭ�i�/_����|O�}&�%�_��W� {�g ���'9    ��ٳgc�Νy;[�v  ��R{��СC�hѢشiSn� ��L�: 3��;   �4q�ر�裏�ִ  ��I�iף�[�Fssslܸ1�ϟ    LM�    SX
��ݻ7>���  �����W^y%����G�e˖    S��;   �422���:ccc  L�K�.Eooo���Q]]�֭���?    ��   �����رcG?~<��  ����P|��Ǳo߾X�zunu/
   ��#�   0\�p!v���O�΍�  ��3::�;(�X�"6lؐ��   ���   n����������'  ��+�vSJ��/��7F}}}    p��   �ǎ������   ����R�]��_����x�Ǣ��9    ���   n��ƞ={��ŋ  Lm)����/��r466ƦM�b���   ��#�   p� ��������J����ƍc���   ��p   ��R�}׮]144  ����{{{㷿�m444�   \�    �lbb"����}�Y���  0��믿uuu�aÆX�lY    ��	�   L�+��O?�4FGG  ��R�{l۶-jjjb����jժ    ��p   ��R����>�������X   �K
���~��عsg<��ñz��    �p   ��R���?��;  ���P���{9�~�}�ŝw�    \;w   ��hdd$7�<x�jc{YYY   \��҂ؽ{��{
�   ���   �Q
�l߾=�9��  �&�:��?�����<�֭    ���;   ��Ha��ؾo߾���   �E
��ر#7��_�>V�^    �)w   �o���)|�F�  �CCC����Ǯ]���G�[n�%    ��    �g�}�w��-�   �-��}�ݼ[�ƍcɒ%   ��;   ��8p 7)��	  �����o��f�����?.   ��L�   ��/���;w���`   �H�.]�A��^{-cӦM���    ���;   0��8q"�o�}}}  p�uuu�+��MMM��}޼y   0��   �R[[[|����ӓ�  ��t�������ob���y�樫�   ��@�   �U�������}�   Lu��^�E��F����    ���  �Y���#��Qc;  0��k�3g�į~��X�ti<��Q,   `&p   f����x��w���-   ��tO�6���/cժU��c�E�P   ��D�   �������C|��� �%]�9r$Z[[��;�3    f
w   `�ٳgO�ݻ7��  f�t���Ƨ�~7n�+V   �t'�   ���}ǎ144   �E�z�w���.6o�---   0]	�   ���ӧ��ދ���   ��.]�����ꫯ�{
���;   �t#�   L[������o����  ��A����x�b�ҥ��OD�X   ��B�   �v���rc��'rx  ��K�Jmmm�����w�>�`
�    ���  �icbb"v����y~  �_���������z(n���    ���  �i��>�]�v���X   �݌���|�|�I<���x��    ���  �)�ȑ#�}��
   ~����x��ף��16o����   ��D�   ��.\�۶m����   `ruuu�o~�X�|ynt/�   0�   S���H����q���   ��:y�d��?�c�}��q���   ��&�   L{�쉏?�8���  �#]��ݻ7<�6m�e˖   ��"�   �t�O��w�y'  ��chh(�m������SOE]]]    �h�   �M��ߟ���Ν�K�.   7_ggg����bŊؼys
�    �Q�  �nbb"v�����l  ��ҵZkkk�򗿌����ڵk   �Fp   n��?�<v�����  �Ԗ�ݶo��~�insoii	   ��I�   �!.\�o��Vtww   �K��꫱hѢx��'�X,   �� �   \W###���Ɖ'��   LO��̙3�����w��ׯ   ��&�   \7{�쉏?�8���  ��abb"���G���{,�/_    �E�   �tmmm���.  ��ihh(�z�hll���z*���   ��p   &M
7���q���   `v��ꊗ^z)V�Z���B    |_�   ��سgO��U=   �˥K��ȑ#yG��<�-[    ߇�;   ������%���@   0�Ƕmۢ��9�l����   �]�   ����X�������   �U����u�ָ����{�   �k%�   |g��y�ر#��  �ϙ���={������'�����    �6�   �5����[�www ���(�]��,.Ey���𤋮����ңKQ(���2��~OMMM��}��先�?�ߚ�T�.]��|hh0.��/���h��\�M�cc1<2W�9���c� �����x��WcѢE9�^,   ���   �*�������-� 7B
�� z��cDMU1j�����*��������X�������ʊ�����b1��K�����beeT/?���,���4�QV������(��,��f�ti"�FF�>�A��O��������q������X����p������|�q�}�C�������qpp(.�fpx$�t�zKגgΜ��[���?k׮   �?G�   ���;��^��� |_��2�����p9�^S,Ɯ9�QW[uu�cMm���Du���zu�Kϋ��L�Sz^(��l������W|��dI�F��r ~xx$7��c鵡��.�P����?0�}��S������o |ccc�}��طo_lٲ%���   ��  �?��ŋ��o���� ��Ԭ^,/��,*J�k�����>�룮�&���Ŝ�ڨ)=����buMT��U�c��:7�s�
��.�{J�]������P^,�;���`i��b�_����x1zK_��틾�{�@���/��R�Z�*{���    q�    �{��ɓ]�}�eQ����XQ�ڪb4��ż��Q?gN�ח�nN���Eu����%-R�-��H3����?>1C�����w9��ן���7:�����?�zz�b�= �|i�ӑ#G��ɓ��OĲe�   @�   ���ٳ��[o��U f�BYD��<������be4ϛ��^���������S��)�\QY��򨫛�g�_x���H���F�Ł��닞��|����=�q��+�GF��a��}۶m���[�l����    f/w    ���r��ĉ��V^V��<5�Q_SM�Rp}^�K����������!���(+�����X��������DoOO���EWww\(M�����s��14< L/����[�n�x ���    f'w   ��Z[[�wމ�Q-� �EE�J��<���PW-�͹����1�4̍چ����vf����<-��_����N�����t���������	 ������裏�������F}}}    ���;   �Ri������ L-eeeQU��W����ǂbol����b�ܹ1�a^�WVU�uUUձpѢ<lhh0߻.tEǅ�����;�t��� n����x饗��;����   0{�  �,���o�ccc�͓zի*ʣ����幕}������%�����)7��k�U5�L���X�(͟���GggG�?��:���s��8���.]
 n��}w߾}q�رx�駣��)   ��O�   f����x��7�ܹsZ 7P��,��s������X�2?̟s���~^c4�+�P(��)VU��%K�|U
�w]茎��8{�|�>{.N�k����w^p]��/��W���{�t�T   `�p  �Y�O>��>�(����룼P��QWY5��+VDKsS,X� �5��ܦ�h(M]}}��	f�t���/�s�W^����=5����S9�~.�/��;��:r�H���ŏ~��X�xq    3��;   �p�����oDggg 0y*R���<�)VDS}],Y�(���4�DCSS���f�bUu,]�2��J�.��F���ўB���ƉSg�����{�!����5�ҥK㩧���   3�;+   0��ٳ'���D ��e9�>�X���X��%ZZ�������9j��@RV�5�an�[V������pt�?gϵ��3g�ę�q��#F���%�w�k��g�&��>�x�X�lY    3��;   �@]]]���G___ p�
eeQ]Q�f�,����X���Fc˂<��GyEe |W�UU�xي<|����htu���z?{6�N��ֳ�h4ƅ������ضm[,X� �~��(�   L�   0�|����'�h�)�^[Y����^U��2�9���7�,��M�R��~����EK��u�����;ݝq�T[�:s6ZO��g����� �����غuklذ!V�^   ��&�   3D����o���@ 𧊅�h���2�^����/\��_ifof��B��ۤ���˯ƅ�sq�̙hm;�J�����@���X��������3�<UUU   LO�   0ͥ��w�y'�;���K�B�I��U�cE4��Ăŋ�y�hZ�8�,��� �.����+n��ࣗ_����Ϟ��S��h�8q�\����D �V���������o�=   ��G�   ����������P �V兲��,�9iR;{�����/�����ļ��(+��I�����u�x����h�\舳�ڢ�d[n=�}�d<&,�f��������������Fuuu    Ӈ�;   LS۷o�}���l�����1��27�ϫM��K�)��/X�[�+�U0�TTV��.�s׃ǥү����8w&�N���'�TGg���؄�;0�uuu�/�7n�U�V   0=�  �4�nп��kq��� ����hHa�bE��sr�}��%_��/�B� |]ڹbn��<��'~Tzmhp :Μ�S�Nű�q�ԙ���q�w`f���{/��?���Q,   ���  `����O>�K�������<7�7�c^Ue�k��2̞Z��ļ���໫���e�n���Ãq��\�=}*�;G�NG��h���L���[�n�'�x"V�X   ��%�   �@������ 3͜b��v��U����e�}i�,^����QUS�Wޚ灍���{Ǚ�q�T[o='Ξ�����8:a�%0�6���~;�-[O=��]�   `�p  �).5��ڵ+&&&`&�/Vļ���[]����0wn,X�<O��e�]��#ޗ�Z�g�C�q�T[�i;G�����=2���������矏'�|2/^   ��"�   S���@�������� �Ϊ+�s�=Oue���F��e�p��XP�����Ԕ-_�6�#OF\�뉎3g�ܙSq���8}�;��Fcx�bL`z�7�x#V�X�7o��   S��;   LA��۷������BYngO���h����%KsC{
��76EY� �OZ��f��u���~=���v2N�8_k���C�72��`��t�R���Ư~��زeK455   p�	�  ���^��8w�\��0�ʢ�x��}^Ue4��y��h_�tY4-Xee1f��Xi^sK���=O��EǙ�q���8z�X����ޑ���q��688/��r�~��aÆ    n.w   �">����v`�+��E}UE��2Ԟϩo��V����ce�* �]��+�π4�=�9����q��X9v4��^������(�v�ԩx��g���>   ��C�   n����ضm[�8qBk;0eUʢ15�����TUV��ũ�}EnjolY �U�5��r�</MDwGG��:'����'�kh4���bd|" �����x饗��{���?   �O�   n��'O�[o����0����E]e!������U�Q����E�WFEe1 �Z���b�4���P���q��h=z,:�rؽw�nF�͗��ݻ7�;?��O���6   �G�   n��������_|���2*
e����4M���*��e+r�=Mm}C �d���������x��j�3�����cq��B\����p��<�����/ģ�>k׮   ��p  ����;^}�ոx�b �l����\S��U1��2�kkr�}��[��pC
�WS=���q��'���9��#�32�#�p���۷o��Ǐǖ-[J߳
   \_�   p�۷/v�ؑo���ee�PU�[���������@����b^KK��~��RW?7��}�G����8}�H?v,.E��Xt��rw�F:s�L��?�c�ϟ??   ��G�   n�h����ԩSq�$pcU�rK{
����ʊʘ�xq�/�uM���	 ����kb��uy����q��X�;g�z�sh4���b�96p�+��w�yg<���   \�   p��;w.��Ӎp�%5�7�TFSM1�UWFuuM��Y�lETTV L'��W�=�ēq���8}�h����sp4:��bd�nI�����hkk��{.���   �\�   pm߾=�������幩���"�VUFM]],�eu,�uu�,Yee� �� �L[�ty��6m�������#q*��ϵ�f����v .�  ��IDAT������կ~�6m�[n�%   ��#�   ����@޶���' �������,�P��Ҥ�{��h_��X�d�P; 3^Y�Wc˂<w=�1.��ę�c�v�p�8y2������`2���Ż�Ǐ�͛7G���   &��;   L�Ç�{����p=4TU�@{K]UeQW�KnY�V�M� �Vu�sc�����j����S�98]C��3<�X&Kkkklݺ5�}��hll   ��p  �I211۶m�7�&S�,����5��T��B!�6��M��V����� &���H\����xi"�FF�����t���/�����<^��x��cc��mtx�k�/�~��|��+�7)��GEŵ}��vq��,���ߓ~oR����g����/�^Q,�]"���+K�w**��+K���ǅ���π��a����h;�Ei�����04�����d��_~9x����{   ���  `ttt�k���ohL��Ծ��*Zj�Q^(����X�zmin�9s��R}���xdd8FGFJ3c�#9t�B�iF���|<r��ޛ�c�D��+/��BEy�U��9_���)9_����=�yeUuا���b�ZX�"��\���y�{{.�ݏ|���5<v��]���.]��w���S�{�X   �p  �h׮]�w��|#��Hm����_S�uUQY(�a�h_�f��vf��A���H��xh����/�P���3.ޫ.�߿r����TU�DUMm�X���t,��ǜ������yz�.��#����Cq��+�h�������[�n���z*�,Y   �w#�   ����H���q��� �!j+�cAm1Ω�b�,j���@{jkolY0SLL����`ib(����p�8<4�/�K����.)$�f���OZ�B�Ś�|��������{u
�פ�5QS[�)�?���)�Z�!υ��rн�ȡ���C�����266o��F�\�2�|��    ���;   |i���~;߰�>R����X����(���Ukr��y��(+���bbb"�.�������+K�����_̡�^O�0��"��/L\��򊨙3'�k뢦�.k��DUm�׎�����Բ0Ͻ��3���������1�;Gcpl" �U����^�����Q[�9   |;w   ���o�����*|gU�XPW�QSQ����޺:��,Yee���&��^�X��+=���)Ȟ����S㺟�L��c��ӝ�/�,�nW��W��7D]CC>
��li�Y��yx�Gq��8q�`�>v4���s����h��߮�t���/��͛cŊ   �e�   p�FFF��_���� �V�BY����9Ŋ(
�p��X�v],^ykn��)~SX�b_OiJ��t�-��{��f���y��ȅ�����I;o��{m}×���W�5u���=3C�P�f���#_D�r�{ϗ����؄�>�7�;��\�2�|��    ���g   pN�>o��F�����)��ESMe,����ұ��ZCSs��m]������itx8�sp�4����@�qOOne׾�]Z������?���Kǜz��C��q�c}Cng���,�-��ʓv�8u�p;�?�:�G��x��ą���m�&�����K/�s�=U��   ��p  �o�}��ؿ�����cAmUnl�,�EMݜ�Ծ�u���p�\�4�ep�;������+�z�s� ;�iaI���<,�ޑC�s�E��ƨO��ω�yM9���~ί���<Ο����Ç���@t�������?�[:oۺuk��G?��˗   �u�   �R[�?��?������T�r�}aij*
��u٪5��ۣe�2�L����ׯ��{R��+�'&&���Ǣ��B�?VUS�E͙�)�^z\?o���)��ea�{7>gO��C�Ǚұh$�ӌ��>�����x뭷bݺu�裏   �/�  ��hoo��^{-FFF���ʢ��2�V�cY�����s[��[WGyEe��511�C�}]]��}��0{O��t���h 3���`�<�O��������˶�yM�ϻ<�kL�B!�ܲ*���@�8|(��=:�{x,�/�f����8�O�����U��    �  �O�޽;�����N��H!��bynjo�-Fy�yjӽ��;Jsg�Ω�.R�=��s�sg>� djc�3�c�����|��J?�jJ?�����mj�y�[r|�P�<U5�q�=���:�������Pt|���;< ����u��زeK,\�0   `����݇wTס����M�����@�M��N��o��%\�Yy�ɻlc�m c�cS%��*H��4}Fq�QT�|?���b��،�>���&�    �7
��z{{599) x��4����v�Ô�phs[��־iK���S��/��>�^���� ��� &_�����[�wk�UM4�H}�"u��QB������^��{�ɑ{Jds�N<
�g��^�\N��v�ڥ_��W    ��p    �hffF~���� �4E}.m
x���jcuڶc��tu���
�!�Ĳ�g5,/���!����� ֝���_����з�{|>��?�jc����ُC�m����sniﲇ�(a��n]�B[B-d�Jd�0�?5��d}v߸q�^x�ꫯ��v    �jD�    P���ǟ�9�C v[��Ծ)��4�r��ұ][�w*��$ౕ��K�Z��f�5��Ѱ� P��ɤ��F�����DU��-�Vۻ�6������h��~c7�[����=2�+z��hr9�4��@U����;Ｃ?��Ojhh     Ն�;    �j
?~\���ہ*��m�Vȯ��Y�v�Rs{�N�U�\6���3���������̞�� ��:^,~�YC��~�
�[A�hCc�Ѿg��g��[��ܦ��G�nZ݁*�-�~��G��/~��{�
    �j��9    @U���Woo��� T'�ӴC�߶�{<�ڽK��(T�S>������4�`�ne_Z�g!��d�J11<d�ǂ5��44*Z�h߇c�r�\³ki�ԍ������Vw��YǠW�\����x���)     �w    @չy�>��s��@u��v��L۾s�Z;�	�U�������v�}~fھ�`J�|^ ����`��;��s+��D����ZM�ֽi:�'
GT�=j�����mvvV�����^{M�pX     T:�    ��r�����@u��v�é��Nu����<��_���ķavk��9 ���.l��1��~�j�#�56�n�f;��Ddo�aV��͟�?F�;P��鴎=����C     T2�    ����d��sssPC���`{�����hL���m�9]n�r��	�NNhvjB���P{.� `�Y;%=�ݺn���x�oP�q�bMM�54�s�hi���K��k�mu/��TN��i���Zt �2Y���}������;     ���;    ����̨�����|VC���nۭ�v����vm۵[ͭ��V�������v#���};��{H� JH6���ب=,Vy(��彾i���U��⟅5�?���ud�:��4���T"�\���@���u���kr�Y�    �<�    ����:{�,!G�
]5��j�e�|��:��Ӷ�����ʑͤ5;5���1;eڧ�˲�	 ʉu|��-�P��6ہ�ئ&; _M����O���߼Sm5^���$3�XJ+�+@�v�{��w�{$     ���;    �b�9sF���P�b>���E�.�y]S�:��S��)���f����� *�r|������n���?�Ge�U������?fR��m��LN��&�PY���;��������     ���;    ��Xx�=j���L.�Ц���{��Z;��s�
���R�Y���531nߧ�	 �O&����=,�áh}�wB�V�R�F�
G�_�yL��i�TMAS�M%2�X(T�B�`�\7==�    �J@�    PQfff���k��T��ˡ��W~�LÐ��W���صW��c�������F5U&ƔN& �+�󚙼o�>]�_�j�вE�-�jl�"�ǣr��ީ[W.����:L��x�Z<�z��hb)�D�  �a``�>'��k���v    �rF�    P1nݺ�s��ie�6B����)�Q��_��7�s�~���4M�|�������};�>=>j7� �,���u�F�!\W���V5���-��./夥�k��c�F�����&�3�Mf��Y;ٽ��v�=�    �rU^g�     �gΜQ� T�i�)�-��S�á֎.;�n�Q�@���=Ӄ�q�L�W.�. ��g-t�{0m�����p{lS��7����EцFFi/����)X������_��i�T���匦��
,ʙ���ѣGu��uvv
    �rD�    P�_��Z� T��a�ڭa��.���إ�/�(_ (�������Fih l�|>g��ƍ�*S�kܤ��-�k�\�����N���Һ���ijk�W[j��Jdt)�t��;P��?gϞ����t    ��p    ��������!w �/�v�9�S��m?��jԱk��w���JW:���٧�P���E Pjr��7?�F���"�Xc�xohnU��^F��Z:��=���Y��o
���x<�0���RZKټ �������k��&��-     �w    @Y�u�Ν;g��(_�a(�u�9�Q��e��kP����ҵ�$[U!�sY�LM�-�V+���>� e'��|'����T�Ԣ��m�\.��,����kia^�x����e��LN��2v�@��v�{��w�{$     倀;    ��9sF���P�L�P�߭-5^��;�n�ɶ���Ꚛ�Ҳ�R�܃i; 8=>�٩I� *K:�����=�Ex����ukq��{�{��]��RP�v�&�T"W��g��(/��wG�Ձ���)     Jw    @��f�:r���7����q���n����.>6�vt�{��T�
�#�J���1;�>1<�TbY  Tkg���	{ܸx^�O��[��ҪM[�������w�L��1��TWا-!�&�3�Jd�+uʅ��v��Y����7���     (e�    e!����T*% ���0���WNӐ��U��Աk�<>���V����)M�kr����n�`  ���_�������ݭ�{��������g5�B5Z�/��X�um5^���Y��S�t�F__�r�7d����    �j!�    (y���:~����� ���۩�W�~���s�ϯ��{յw�\n���2锦�Gii �)X���`ָu墜.��m۪���[s{�����Re���p����l*��xZ�s6�������ӡC���0/    ��    ��v��5}���e&�q��Ƨ��e?�#�~�EmپC��6-�  ��\6k/���6Vg��7�mS�q�3���tt�t��1�0T�s�����tN�񴖲݁R����w�yG�������    @)!�    (YgΜQ� ���ץ�Z�B�G���u����K;�e��XoV�njlD��jr�ҩ�  ��Y���G�����|jڲ��7�l��ޟT��A�P��E��0+Zc1���bZ�{ �+����?��~�;utt    �RA�    Pr
��>�����@y���j��~l�۴��oj�J�}��	M���M�VS�r  �/�L�^�M{8N�55�a��m���?���1T�|���MM�pw����_��a�c�TY;:}��g�9��_~Y     ��    ���H$������ J�������֧��a���Ҫ]���b�M��Z�/؁���w4;5aU  @���s���ճgT��i�Vm�ڮh�\���Y��Ǭ�{Mԩx&��4Aw��ݾ}[�ӟ�$�4    �F"�    (����裏�-��.+���V��尟�tti��_�6V'�����f&����A{,�  ����Y{�]�,�F�۶�i�6�7�|.���V�{ryI�,�vhGԯD���xJ�I��@)�����Çu��!��n    �Q�    JB__�Ξ=�B�  ��0�z�G[j��9�[;�k�/)�k/��jr��h�V&�  (����\��.�[�Z۴yk�}o��_��J�w�����F��� ����%���;z�7�    �F �    �p�}��p_YY��c��������B���Z6������hjtD�<�\  Pɲ��F���jr�C�4Vн+�Skȣ�xZӉ���#����ѣz�W�u�V    ���    6���~��q���	@�q���n����v�v��y[�v����k,�N�j��؈
��  @���LK��T��1fGا�G�iM.tJ�����'�h~~^���     뉀;    `C$�I9r���@i��훃^;h�"ؾn2�&��j  U��4���W<�hl�Fw��@I�ꫯ4;;�?��    `�p    ����رc�d2P:L�P�߭�Z��K:�����P��ݒ  P�<V�{�X��
�ǿ	��F�v�{����׿�UN'    ��c�	    XW������O�BP2C��{�V��3M�Ԗ�;���_+�VWryIc�w4^�S|  �;��w��L2�1����;���7�T(     k��;    `�\�r� J���󹴵�/��ߍ�{^����aa�d�i����'G��  x�1jWا�G��f�Y�8���jr�ӟ����&    �V�    �ũS�488( �!�s��֧��a?oli�����±zau��9M��j�������   O��4��+�i|)��)���F)
:y����G۶m     k��;    `MY>�?���1�x����S��贐l�����o�_�������>>tW�,�+  ��*��:���i4��B:' ��:�s����q�۷O     �6�    �5��dt��-,,�ƪ�����Zϣ�A�MM����75�g�x{85����ӧt2)   ���S�cNͧs^Li9�N9�F���/�s>���     XM�    kbiiI���R�� l��rK�OQ��~mh��~���-�󙝚���~��P*�   �W��T�>���tO*�+������/�i�    `5p    �������(��
���j���ﶟ�D��������)�xóI./id�OC�ohia^   �x�SaOPS9��SJt�����>�������I    ���]    V��ȈN�<�B�@�<S[j}j��e��5����ߪ���`�3�e3�;�{��5;y_+++  @i��}c>��^�������䙗�eaaA���:$��/     �w    ���q�>��s�p��ZB^5�|*>���U��_�k�~��Cx:+��éI�뻥�;}ʱ#  @Y0����b�:�K�����i噣�"�J����z����F    ��"�    X�Νӭ[����Q�ǣ��>��N�:������\n��t�jlp��'�  @yr������\v��T"# k/�˩��G�����,     �w    �s�׿����AX_u~�l�92C[������ˤS����ۚ��/   T��TGا�A�F�i�&ٙXk�BA���?���/���[     <-�    �gf]�<r�fgg`��x��V��-�������[�?)��krdHC�ojjt�~  ��e-
�����ix1��l^ ֎�������E��׿     O��;    ���R)���{J$�>�.��j|vs�%ڰI{�;�7����ZZ��ȝ>ݺ���   P]j=N��M���R9:k�֭[������      �w    �S�.L>|X�tZ�a��r9L����\�߸P8�ݿ����;���;�s���&��4t뺦���&A   T��ϥ�ש�DV#�)�9F���ؘzzz����4M    �s�    ����z{{�ϳ�;�����A�Zk�r|��$�Ш���d�~��̴�nߴ۳�   ��d���n��\_J�~qs����]�p��!��n    �S�    ��ݻwu��i
l��%+ʾ)�Q[�_.���v�!�������h��u�=�   �s��c��n��}&��շ�����{O����+��/     ~w    ��u�Ξ=��m�T�ǩ�H@��{���r���K�>+�n��G��)�%�  ���u���ks �������\��L&���_o���jkk    �!�    �YW�\��˗`�x����j���V�-�]r�����l:�{}7�`{|~N   �j��[�L*�{Ie,�VS.�ӱc��ꫯ���^     �7�    ��t��y]�~] ֆ�0�R�UK�'���_�u�.��v   �=�x�^�s)�uj,���rFv4VM>��G}�����jmm     ���;    �G�>}Zw����������?'�(��I�*��ibxH׮jvrB   �z����x��wih!��tN V��ʊ}�������     �p    ���ǏkxxX V_��T{دZϓ���ڽK�U���yݾ��[7�I�   l�ӡ]��p����\^ ��r?{����v�b�2    �#�    �Q(t��1MMM	��r�������>��F�뺺U-VV
�֝�W5=>f   �R�8��>��DF#���U��p��%�R)���    ��;    �[V�������ܜ ��w�1���Z�\󩿾�m�|��*]*����ۺ{�k%��   J�Q<�o
�U�sid1��d�E��*�~��������V    ��F�    `�f�z�w���$ �'�q�=�W��x�ﱵ���i�{0m����  @�p��:�>m
�5��T<���300`7�<xP    ��E�    �d2�w�}׾�:|N���^�w?�����ڴe�*M����{���K�NM
   (W�bֽuA=Hf5��R&_�g7::�?�P����     Չ�;    T�x<�Ç�[@x~�!��������ںw�4MU�T2��[vc{ryY   @�����85Oib9# ����:z���|�͊�    �w    �b������Q.���W�q�3���X��ٶ}�*��̴�޼��������  @er���������|RKټ <���99rD���I�    �	�@    �Rccc���U(�u:��S푀��U���MM��DU�V����{v[��ب   �j�w��[ЃdVË)e+���<��[o��^�97    �tp   �*t��]�>}�p;��Ц�G�a��Ըڶu�R9�f����Tb).   �Z��\
{���� ����L&��_��W    *w    �2�n��ٳg��B{�<Bn�:#�<ksz��r��c��I|a�����V>�    �e�������bJ��́��N�u�����
��    T6�    PE���k]�pA ���4�V�SsȻ�����e����܃iݹ~U#},�   ~D�ǩꂚLd4O���3�Tr��zzz���+�
    P��   @��z��.^�( �.�s�+��a��{m۱[�l�x����W/ivrB    ~�aHM��V��BJ�iv>�F>�Woo�^{�5���	    P��   @�r�= <�ˡ�H@��4���E7�
y����//*>?'    O��0�3��\*��Ť�y�܁'U(��G����    �<�   ��}���ꫯ�陆��oq�����jo7�~��$�Ʉ�޼��׿V:�   ���:U�j|9��Kis��r?q����?���I    ��B�    *؅���_�ӳ��;����u}_�0���[�biqAw���[ו��   `u9�� �Q����bJK�� �<+�~��I<xP---    T�    P�Ο?��ׯ��q����}j
z7���ڶ��h��NM���eMie�I   `�\��5����bJÁ�e�WO�:�����jmm    �2p   �
�駟���O �N��VW4 ��ܰ�ö����`��//��v    ���ѩ��V����BR�ivQ~�r?}������jkk    ��p   �
��'����_ ���4������߇��Wc��_�_)�&���֕/�pzJ    6��ahgԯߴ��s~�r?s�8���    �w    � 'O������Ө�[��A;��ںw�4ׯ=�
�����K�8�P    JK�ϥZ�CC�)=L���+�~��Y�1!w    (o�   �B�8qB����'�q��*�u�Tl�޵.�S(�5zg�nl_Z�   ���.�]�#~�&����Y�Ν+�{���    �<p   �
p��q��i
z���al|k�cu�6+���{�Y�뻡����\^   �����=N��ӚJd��YM��ϟW.��Ν;    (?�   �����j||\ ~���PW$�p	��?�u�ڵ�g�)ݹ���\��~   �<9MC�^E�N.$������K�.�a�]��g�4    ��!�    e�p;�d������j}2K���1�˭����:=�L�m�C�����    *C���uA�.�5���!^ �e���B���|��^    �|p   �2T(t��QMOO�O�ꎅt;T�Z;��t�^�|:�P��_ڭ��\N    *��4��ƫ�ץ�I%s��������߿_    ��@�    ʌn�������q�!��������l���;Vg�t��   @�	��W��RF����]V��ڵk�9�_|Q    ��G�    ʈu!������� ���۩�h@Aw���#�6nz��A�   �n�a�-�Q����\R�<m���B�ׯ_�i�4�   @(���     ���v������ڭ���Z��(�v�.�����J�   �
�z�>�1��}9c�z����n�^x�    Jw    (���z��� �0�ӡ�j=.�����O�u�   �k��87r��|Ri�܁oY�>���k{>�o�>    Jw    (===�������=��,����6om����_O�   ���u;��.��xZS�� <b�ܯ^�*�ө]�v	    Pz�   @�����߿/ ��u:��̈́�hk��]H�������ו�l   �d����Z��V��BR� <r��e���;�~g5    ��*ϫ�    P%N�<���q��:�[ۣA;�Q����M[�~���Yݽ�n]�X|L�"   �g�:r5����TV 5����cB�    PZ�   @���?����!�.�i�+���l�]2��Y>����v�=�L
    ��5���4�tjp1E�;���/��r���C    ��@�    Jп��/
�w��=���r�*wm�w~�B��ᾛ�y�����   ���t;uw>��LN@����Ϟ=+�0���.    ��#�    %��O?�ݻw�ߜ��ma���^U���f�o��o�wt��9--.    ֒�ahW̯�DF�S���r7MS[�n    `cp   �b]H�����x]��S��m۱˾�����t��y-��    �S�߭�ǩ���♼�jf5�[�N�S---    l�    P"Ν;�[�n�� H��5xد͡�hm��r�y[���G�����   ��b-&�hl)��xZ@5��˝:uJ$�    ��;    ���/�ƍ����Ю��.�*M(�g~���q   @)0��5�Q��T�\R�|A@��B�O�֟��g566
    ���   ��t钮^�* �4<��0U"�   ���ˡ}u-�4��
�V�BAǏ�_��544    ���   ��ꫯ��p9Lm��    �N�PWا�ǩ���
+�����8�^__/    ��!�    �
�_�xѾXT�Z�S;�Br;L    6^��e7��'����FV�����_]�XL    ��A�    6��k���_�vFql��iK�O�a    P:|NS{c�/�5��a�>����o��p8,    ��#�    �l``@.\P�<�nm��pz    J���%�����'�)rG���r����[o��`0(    ���
2    ����}��'4��������i�    ���ǩꃺ3��\:'����y;vLo���<�     k��;    ����I�8q�p;���4�	�!��`    (7��nGԯ�匆S��M&�ё#G����Mn�[    ��A�    ���̌z{{U(T��ǩѠ|.�     �)����Jd��I*�ROO��z�-��L    k��;    ����e{�bkc�����W[�~    T��Ԟ�_��)M'��I<�C�    `�p   �5d5:���{�f�Ћ��r��*�u	    PY���Z�"��.$�+��sss:~��^}�U    Vw    X#�LF���r�Q�ǩu!yl�    �,�u���>�D��P=&''u��)<xP    ��C�    �@�P��Ç�H$T��W��C    �*�s��hh1��;١z����ܹs:p��     ���;    �������E��i����    �����������BJ����Ν;�x<��/)    ��#�    ����W>Pm�n�vՅ�u:    �^�>��.���J�
��͛7���={    x>�   `?~\�MSЫ��_�a     ���޺��Χ4��
�t+++�r��~����    xv�   `��={V������0��!�     �ɚ3n��4�p��bZ�����>���VKK�     φ�;    ��˗/�����thw}H~�C     ��F�[A�S}s	�������z��W���     ��#�    ��ƍ���/T���jn���     �9��}u�]H�a*'��
�8qBo�����     O��;    <����?^+l��*aRg$�MA�     x�⤲;���rF��8��J�����ӣ��zK�`P    �'G�    ���ȈΜ9C�U��rhg,����	    �g�p+P�c�%�)p^��q���ߖ��    ��pE    ���̌N�<io7T��ϥ��ݶ    ��q;�B}P�sI-dr*U:��|�����2MS    ��G�    �R"�бc��&�������'� �    X=�"�1�F�i�/�T*�|���~��!    ~w    x
�\N�V6�P����hPu~��    �k)���G~���)VVT���9�:uJ    �p   �'T(�p�ոT:�ˡ��!��    ���|���T�\R�|A@%Յ���/    ���   ���������J���[�    �^.����?��B&'�������F;w�    ��p   �'p��MLL�t�5>m���0�    ֟��zg̯�xZ�Ki�feeE�.]R Ж-[    �>�    �3�\����>��a�U�w    ��d-�����4uw!��ʊ�Jb�ܭB��^{Muuu    |w    �	w�ܱ�@%��]���     ����*�UM��%��T�B���Ǐ뭷޲��    �F�    ~���>���Q	�T1�[ݱ��<     �&�rh_]@�sI-dr*I.�ӱc����o��fW=    x��;    ����E����MJ@�j��ik�O�A�    P��E�;c~���_J�$�tZ===v��i�    p   ���d2z������T"�i�;T��f0    @y��fo	y�w�\H)ώ{� �x\'N��_��    �   �wX�����ݜT"�ˡ��5�9i    ��:�˞�ޞK*�g�=T���)}��z�W    Վ�;    ��#G�؍I@%�x]�Y���    e,�rh_]@�&��e>T���!�B!�߿_    P��   �7>��#����DMA�:#�     ({.���X@�I=HfT�k׮)���S    P��   @����5::*�uDjy    @%1�3��ij4�P	VVVt��9;�i�&   @5"�   ��Y�Hׯ_Pi����!E�.    P�Z�����̧TXYP	N�<���zK�PH    Pm�   �jccc�pႀJ�s:��!d�    P�b^�<1S�&�-rG�+
����?��9�D;    TfA    �V<׉'�m�JR�qiW]P.�)     �E���޺���Z����L&�cǎ�o��    ��p   P�r���9b��dSЫΈ_�a    �j�q���B�	ͥ9�򷸸�S�N����   �jA�   @U����L&T��Z_q�    @53iGԯ�xZ�Ki�nllLW�^����    Հ�;   ��s��	���
��Pw4�:�[     ��-!��NSC)VV������׮]SMM����    ���;   ��b5ݻwO@�p[[�ׇr3�    �5�\��η����|Y!��g�*+�
    *W�   T���!]�tI@��B�V��
�    �r;��.���J��ʕr�裏����]^�W    P��   �
sss:u�}��~��cA��     ���:L���7��b��;�W.�SOO��~�m�&�    *w    /����ѣ��x����=�A�    �'�4��uw!��dV@�Z^^�ɓ'�ꫯ
    *w    �P(�ȑ#J��*���_�5>    ��g���>���F�/B�����_|��^zI    Pi�   �h������;�|w,�z�G     ���=r���ZP�n߾�h4���N   @%!�   �b]�xQcccʝ������z��    �Z�.{�}g>��
1w����ϫ��V���   �J��q    ��ݻ�ꫯ�;��Ԟ��]    ���:�+�׭��rB�(?+++:~���~�m��~   @% �   �������������\�m���a
     ����8����Ä����r���u��1����ir	   @�#�   ���R)����P�b$�[��Ү���!     ���S�c��%��������_]    P��   �V������d2�Yc���Ѡ��     ��ihgį����R9����:{��~���	    �w    ���WKKK�Yk�O��~    ��g�#���BJS	JP~U__��۷    �w    ���˚��ٻ�/����㯻�]f�aeSDC�|�6mOlN�tM��&��6�Q������ *"3,�,�ܹ��&]�����<�|��0?���~���ʕ@7{tC_��   ���C����\�=�&�V+'N��ƍ�iӦ   t#�;  ��>����W�
t��:��M�X�	   ���UR.$ߞN������^�O~�T*�   t�;  �����s����C�F�R1On�@�+:   t�ͽ��|���������Di4���~���~:   ���9  е��f����m���Q�\ʁ-��W�   �i�ZΓ#}936�FS�N�h��=z4O=�T   ���  �Z�=�\&''ݨ^.��[S-��  �����v�>:��;]�ټys��   t�;  Е�z�\�r%Ѝ�+��<0�9   ��7�}mS;r���\3�-N�<�M�6�?   �@�  t��>�,��կ�h�֓'7�T,   �.��ڑ�ٱ�L���A��ʡC���3Ϥ\��   �ϛ  �U�����/��@��W��@��   нz�z�bco޿1���;�avv6?��O���O  ��	� ���l6�a�F��l�汑�h�  �����<9җnLelz6���!ǎ�w��   t2�;  �5�{�LLL�̓�����+n  �5����؆z>��|9%r�;�?>�6m��?  �N%p  ��[o��+W��͎�zv�   X{ڑ���zz��|>q7�N�<9��  �N$p  :�g�}�_��W�n�gC_�   X���\L>���Z�V:�g�y&�l  �<�T  ��6>>�_|q���E�P�c����   `}x���R�����}ˢ����������/��/  �4w  �c5�����?M��t�R�������^	   ��<�ۓr!���T$�t�۷o�رc��w�  �N"p  :�s�=����@�(�yrS�j=   ֧M�����|pc*MK�t����g���ٷo_   :��  �Ho��V�\��=�b��e0}=�    �ۆj9�o����ij��p���/�#��7  �� ��s�ҥ��W�
t��b!_�< n   ��P��'6����̩��`�V+�3�<�rYF  �>o&  @G���ɋ/�8�ݠ����^q;   �TJyrcoΌM�!r������СC����   �6�;  �Q����m�0�A��q{]�   ����o���c�����������5���o  `5	� ��q���ܸq#�j�RlH�,n   ~��_G���t��n|��lݺ5   �E�  t�O>�$�Νt��,����    ܋����FzszԒ;��^�O~�T*�   ��;  �ꦦ�r���Z��|���?�:�JI�   ܟ�w�'G���g暁N�h4r�����?�s   V��  Xu?��O�M�����r`��   X�z��'6����d���P7n�ȉ'��o;   +M�  ���_~9�n�
t�v��uq;   �ڑ��#�9=*r�s�;w.=�P�o�  ��$p  V�G}��?�8���+��<�q;   �D��v�ޗ3c�n���LG�ɏ���j�   ��;  �*����ꫯ��j:Y��[�S,   `)UK�<��7g�&3%r���������я~  ��"p  V\����~�����d���r�`J�v   `�T~��>:�I�;�֭[y�������  X	w  `Ž�����Ɇj=��恔
�v   `y�o�{b�/g�&31k����f۶mٹsg   ���  XQ|�A>��@'����M�v   `��G�{sF�N�:v�X�lْ���   ,'�;  �bnܸ��G�:�`��'-�   �������щL5��N�l6�����_��_  ���  ��h~<��s�?�ST�9�yP�   ��v���H_N���@w�ܙ1yꩧ  �\�  ��8x�`&''����oL�(n   VW�ȝv�<��Cٽ{w   ���  Xv�O�ΥK�����4����   @�hG�O����wrw��$���Z6oޜ���   ,5�;  �������o:UoO)_�:4h   �I*�K���K�w�,��9������?��O  ���  ��ir<����?��˥|}ˠ�   �X�R!Ol읏�g�������9v�X���  `)	� �es���LLL:Q��?��J�   �NV+�䦾�w}"�"w:����cǎ<��#  X*w  `Y�6.^��D�C�v�^�   ]�V*�ɑ��%w�;����m۶T*�   ,�;  �䦧�s�ȑ�Z��<���[���   @ש��ٿ�7g�&E�t���������~  �� p  �ܿ�����h:�|ܾup~�   �����#�3c�i���cccy���o|#   �%p  ��ɓ's�ƍ@��)���z�   �n��#�9�;��w�͎;222  ���  K����9u�T�������-�v   `��oG�zs���D�W��ʳ�>�b��  ��	� �%�l6���|�:I;n�������  ��e�R���#ro�.G���ɑ#G�W�W  X(�;  �$���LOO:I�Xȓ��W��   �M����G'"q�|��g��㏳gϞ   ,�~  `����\�|9�I��B��4���W_   `m���w���nM�a�����g۶m���  ��r�  ,ʝ;w��k�:;��l��   `=�T��\���ܲ��k6�9t�P~��  �~	� �E���~����@'yl�?�{�   XO��V2;��gw�Vۭ[��_�"��  ��!p  ��ѣ�}�v����З���   ���}�:�����L`��;w.;w�̖-[  p��  ��|���y������z��   ��=2XK��ʵ���jj�Zy饗��3Ϥ\��   ���  p�fgg��/:ɶ�Zv�   �d�p=s�dtZ���jO>|�p����.   �B�  ܷ������)��V�w��   ��;\�܍Vn�mV�_|��g�f���  �C�  �}9u���at���<6ҟB�    �K�P�c�9;6���ji�Zy뭷�cǎ���  ���  ��Ν;y��7�b�Z���k   ��J�B�Л�F'2�hVK��̡C����O  ���  ��g?���!t���R��y0���   ��)ybc;r���9��X=����#*��ַ  �� �{Ҿ>���ہNP�)������Y    ��J�8���̌ȝUt�̙�ݻ7���  �m�  �t�ƍ���ہN�>�������    ܻZ���7�sfl2�f+�Z:�g�y&   ���  ��~��ٴ���k/������   `A�zJٷ���c�Ѹ�Z�����������  �	� ����ѣ�����b��'6���    n�R�ޡz>�5�VK�������{��lݺ5   ���  ���]��s��:�c�2\�	    �7R��L��������_γ�>�bэ�  ��  �U�����-8�vo�͖�j    X:��*�;�̕���j�����E����n   ~C�  �V�����&V�C�l�   ���s���f+קf��O>ɥK��}��   �	� ���}�p��j��[����    �|��2;�ʭ�F`5���y��gS.�X   �;  �4�ͼ��K��6T-��
   `�<����c������F��W^y%����   p  ���fff&����R��<���   `E���<ގ�G'sw�Xi��y>����ٳ'  ��&p  �Ӆr�ҥ�j���9�e`�P   ��S-�#r�L��
��'Ndǎ�T*  �/�;  0ovv6G�	��R���mH�\
    +�����6����T�-�;+��h��_�?��?  X��  ���~>r��R($OlHū*   �j���g��oNV���hΝ;�}��  X�T  ��a�իW�����P�	    �oS�'�s�|6~7��Z�VN�<�;v���7  ��#p �unzz:���Z`5�����    �9��W3;���ə�Jj6�y�����0  ��#p �u��K����v���`=    t�]C��4�����u��ͼ��9p�@  ��E�  ��ٳg3::X-j=ytc    �\���щL��VҩS��gϞ���  X?�  �N����7���ޞR�o�O!    t�b!y|co޽>���f`�4��>|8?��  �w  X�<�Fõ¬��b!OnH�X    ��R,���9=:��V+�Rnܸ�s��e߾}  ��;  �C}�Q�^�X�B�����{J   �{���g��nLVJ���ɓ'�k׮T*�   k��  ֙���ǎ����2T�:
   ЍFj=�1��g�w+��]��������   k��   ֙�fvv6�vֳ��    ����j��\�򝑕s�ڵ\�pa~�  X��  ��\�t)�/_����Jv�   ��g���F3wf�+���_ώ;R.�]  `-�?  ���µ�jVZ���#�   `m(�}�yot"w�|sde4�9r$�7  `�� �:��K/��ݻ��V)��恔ڧ�    ���>�7���щ�5E�-���J�o�  `m� �:p�ڵ|��'���n��q{�T    kO�\�c������cǎ��g�M��#  �Ew  X��f:�V˂+ﱑ�T�z   �e��r���Ӂ�0333���_�e  ��Ge   k\�#���$V�#C�l�   �����J��|19X	/^̾}��u��   k��  ְ���|�ᇁ�����G�z   ���k����\n��V�+���g�y&�b1  ��!p �5�^H�����J)���   ���PH�m��{��j�.��{�nN�<�o��  ��;  �Qo��F���+�Z*�k�Sj�f   ����Pϻ��i���>Ⱦ}�2<<  `m� ���O�>XI�B!OlH��:`   ���^.���z>�9�VK���j�����K��  `m� ����ϧ�t0+kT�f   �l���P_%���,����������/  @�S  �s�ԩܼy3�����j    �7��W2٘��t#��ڷ��۷/}}}  ���  ֐������[��4X-g�po    ��3T�Tc�Ǎ�,�V���_~9?��  t7�;  �!/��b���+�R*f����    ��V*��p=��&�h���ƍ��㏳gϞ   �K�  k��˗���VJ;j����TK�    ��R/��?�9=��˥��u�ĉ�ڵ+Ţ�  Э�  �F���+�XQ{7�e��   �?lC����*�t�n`95�?~<O=�T  ��D  �5��^���d`�<8P˶�    �W��+�l�el�XN/^�O<����   �G�  ]nbb"gϞ���j9{6�    �מ�Z��_=��ri�v�ꫯ�駟  �}�  ��<�f�a+�R*�̓)
   ��U*��p=��&�h��e||<gΜ�_r  ���  ��G}�����JhG�_�<�j�    X�z��݃�|xkz~i��/���ݻ7�J%  @�� @�j��;v�+fT�F   �xk�<����;3�����~�ȑ����m  ��L  �.��+�dvv6��e�@-    �T��U21;��w���ʕ+�϶m�  t�;  t�7n����0T��ލ�   ��T(�w���F'3=�,��G���g�  ��  Ѕ^xᅴZ��r���yb�@
�    ��+ylC=�G'3�'�dzz:o��f���o  �|w  �2��Nn߾Xn��}#��;    ,��r1;����t`��={6���O___  ��&p �.2;;;�2+ᑡz6�+   �嶹ޓ�ٹ\��,�������J����  �lw  �"����\`�m�U��Po    `���eb����(�ctt4/^�Ν;  t.�;  t�+W����ˁ�V)����    �J*�G��ywt"s�V`9����y��S,  t&�;  t��^z)��
_=�7�G�    ��j�Bv���ͩ�r���������SO  �Lw  ��E��):,�]�2\�	    ���Z9��=�bj6�.\��dxx8  @�� @�k��gΜ	,������    V�ΡZ�4����,�#G��G?�Q  ��#p ���K/��l�S�\��    ������p=�Nd��
,�۷o��?Ξ={  t�;  t��W��ʕ+��T($�7��X    t�j��=C��c2��Z�VN�<�]�v�X,  �w  �`/��r`���П���C    :�p��m}�\��	,����������v  �Ρ`  �u���ܹs'��6�V��@-    Щ����\�g�K�>ȁ���  �3� �5����XN�r1�F    ���ճw��wG'�h�K��j��ѣ�����   �A�  �W^���l`���Sj�    �Z*���ZΎM�ڵk�r���<��  V��  :���xΟ?XN{7����   ��1T)硾J.O��R{��رc��O~  `��  �ü����a�l�f[-    �m�Ts{f.�s��499�w�}7  ���  �A.\������ri_���H    ��z�P�;�'�h
ai������\��  �j�9  t����\
�B�4�r�    �V�b!�����t`)5�?~<���w  ��;  t�7�x#��dX>��3\�	    t��ZOn�����l`)}�駹u�V���  ��;  t�����9s&�\�j=yd�7    �V�����\���Ri�Z9r�H~��  Xw  � /��b���ˡ\,f���    �ZR,${��9=6�f�X*�����g���  V��  Vٵk�����ˣ�R-    kM_O1��+�t�n`��W�O�8��;w�X�m  V��  V��Ç�?��r��_˖�j    `���ۓ[w�5�L����l�z��ɟ�I  ��%p �U��{�e||<��=����    X�
�B�������6���tΝ;����V��  �J� �*i6�y��7ˡPH�����    ָ�b!{�jy��T`����9r$�w  `�� `�=zt��SX���2P��   ��1\-�ޞ\��ݕ�s���\�~=�6m
  �2�  �
�����G���z%��   ����Zn��e��,��Ǐ�G?�Q  ��!p �U���/�_m
K��T̾��    �zT��yt���F'3�j���۷s����ܹ3  ��� �
�y�f._�X�R*    ֫z���*�p�n`)�Z��<yR�  +D�  +쥗^
,�����+   ��nko%�f�26�,�������{��׾  `y	� `]�t)ccc����Sʮ��     �a�`-�3�m�K�ԩSy�'R,�E  ���  V�ѣGK��ճo�?�B!    �(�5X�7�Kann.���/�g�g  ���  V�ٳgs�Ν�R{x�7�՞     ���Z9��z�O7Kᣏ>�7���j�   �C�  +��lί��R믔��`=    �o�s���ىܝk������^�_��_  Xw  X'N����L`)�<>�?�    ����Bv�r��T`)\�t)7o����p  ��'p �e��Ϟ=Xj��{�W�Z    �P����=�br6��?����  ��  �ّ#G277XJ��r��    ܛ���uw.�s��b�����իy��  ,-�;  ,�;w��O>	,�R���7    �w�B!{�j9=6X
�����  ���  ���Ç�j�Ki�p_��b    ��3P)塾J.O�kbb"~�a}��   KG�  ��ڵk��/KiC�'�j    f{57g��m��7�̞={R,% ��"p �er�ȑ�R*�ٷi     ��
�ޡz��H��,���lN�:�o~�  ���  ���r�֭�Rڻ�/Ւ     X�z�8�������b�>}:H�,� ���?k  XǏO�e��������}�     Kc[oOn�m���\`1��f^��<��S  O�  K������T`����ytc_    ��S(�g��S�'ҴW�"]�x1������   �#p �%�^ii����R*    XZ�R1��r��t`1ڷ����k����  `q�  ���|������ʖ�jF�     �ckoOF�gs{f.�W�\���x  ,��  �H{��̙3���S*fφ�     �k�P=�\�H��
,T{���������   'p �%���[ogI��ЗJ�    `y�J�l����Ÿv�Zn޼����   #p �%�h4r�ܹ�R�W���    `el�dt���ٹ�b�Wܿ���  X�;  ,�cǎenΡK�T,�ё�     +��ճg��wG'�jlttt�	  p��  �H333���Keφ�TK�     +��\̃��\��	,F{���?�a  ��'p �E:r�H��f`)�z���    `ul�f�n#S�}Y��7o�/��֭[  ��;  ,���T>����R(
ylc    ��S���3T�{����x�����O  �?w  X�W_}�z;Kf�po�=�     �����m}�\��	,���x.]���۷  �ww  X�;w�����0P-g�`=    @g��_ɍ�F�猜�p'N�� �}� ����+��Y�B!�F    t�R��]C՜�
,���d>����ٳ'  ��� �ܾ};��y
�B`�����    ��U���ۓk������/)p �� p �x��K��RΎ�z    ���p57��ef΍�,���tΝ;�}��  ���  p��_��/��"�X� �؟��     �c������܍��B����w  �Gw  �O���j`)<4P�`�k    t��rFj=��,���LΞ=����  ���  p�����Ū���9�    �;����L#�f+��N��_q/�  ~7�;  ܇#G���rx��=:ҟR�    �;���_���w1;;�w�}7�G  �w� �=���Os����bm�W2��    t����\�j���\`!Μ9�Xq ��C�  ����_,V{�}�H    ��S(�k��wG'�h4�� � p �{����֭[���9ܛj�2    t���b�������B�>}ڊ;  �w  ����Z`��zJyh�    ��=�_͍�Ff����������  ���  �\�v-7n�,֣#�)    t�R���k���T`!�  �	� �8v�XZ-+<,ζ�Z��=    ֆM�r���rkf.p�fggs����߿?  ��$p ������,FO��]C�    ֖]C��s�N�6RX�w�yG�  ���  ~��G�Zog�vo�OO�    `m��
y���Kw�����LΝ;�}��  �/w  �n޼�/��2�C��<�_    �6=�_���l����j��� �� ���ꫯ�������     kW�;�#ռc*p��������G  ��  �[����/�,Ǝ�����    �m��rFj�N7��ԩSw  �o�  �[���[�V`�j�b�    Xv�rkf"��o�ܟ����?>�w�   p ��cbb"��y`1�n�O�X    �>���_���Ӂ����o� ���  �9r�z;�2R��?    ���@oO������\�~��w>���ر#  ��	� �i_z����B����    `}�9P�����:y��  "p ����W_��΢l��^.    X�*�l��s}����+W�d۶m ��L�  �6===�',T�T�Ã�     ���Ռ�m�iO��t�ĉ�˿�K  `=� ��;v,�f3�P�7��T,    X��c�U�ٝ����իW��  �+�;  |eff&/^,�`���}�     �=�_͗S���3�����/~���� ��J�  _9~���v�P(d���     �F��Ǉk���T�~ܾ};_~�e6o�  X��  �{�����z������+    ��X-g�����F�^�Z������ ��H� ��w�ĉ����T,d�Po     ~�G��5�H��g7n����x  �� �u�ܹs��j��R1     �M�\��z%W'g����������  Xo�  �k��^ff*�0�=�<4P    �ﳽ���ӳi4͸s�^�:�Q�T  �� �u���,Ԟ})    �{�����������j����������  �z"p `ݺp�B&''1R�dc�j    po��˹6U��l3p��g�g�b�  X/�  �['O�,D�PȞ�}    �W�B!;k9=jx�{�l6��;����F  `�� �.]�~=7o�,���z��R     ��@O)#�rF��{u��Y�;  �� �u���ぅ�)��`=     ��@57�6�l�I��ȇ~�G}4  �� Xw&''s�ڵ�B��؟R�    �����y���Kw���;�#p `�� ��=z4��i�_��-��     ,ƃ}�|19�Y3�ܣ�x��˗��C  �:�;  ����l>���B��M�`�    X��%�;�9k:p��z�-�;  �� �u�7������Sg~��_��g8
IX>���wk�)W���S�����ڿ|�U�hW�lY�@� 3�l�ȑ% �������K��t�G�;��n�i]��.    ��p�V���vl�{f�ɼx�"���brr2  `�	� ȍ,l���	8�l�=[o    8K��VㇵV�I]�~=����=  `�	� ȍ�7o���^�i]��c���	    8[�B������ĳg�bgg'��j  ��Rh  ��}�]�i�Iį&    p>��w��������;�����o�  0��  �������	��ǣ���     8�R!.U
�|g?�$?~�n7�Գk  ��� �\�������*��d�     ���F+���6�9�l���o��/��2  `	� z������pZ��ע�&    p�*�4>���ik/�$��k����ي;  CI� ���ӟ�pZ�b!��T    �"|4R�������q�x���q�������  ��� �����+++����z���v    �bd�I~8R�ٍ����s�� ��$p `����G�z�n8��J)��+    p��k�Xj����g{{;���bzz:  `�� Z�n7fggN���     �h٩��Vbf};�8��ύ7��c  �0� 0�n޼�N'�4.��1^-    ��p�Z���B4�<��x+++�����SI w  �֝;wN#������    �ٯF+q{�pׯ_����:  `X� JO�<�V��N��h-�%�I    ��5Z.�d�k���y��qt��H�4  `(7  J��N#M">�    @?�d���N�z����t:q�������  ��� ���-������G��(��     ��^�V���cŝ�ݾ}[� ��� 0t���?Y��T
i�Yo    ��ߍVbmg?<��8;;;������  �N� �P�v���ѣ����z;    Ї��4.�J����6��ύ7��c  ��� 0Tn޼�N'ऊi�V    �}<R��;��ur)�XYY���ݨT*  �L� �P�s�N�i|2V���v    �OU
i\�c�eŝ�]�~=����  �A&p `h,,,D��
8�,l�h�     �죑J,o[q�x�?�n�ij� ��%p `h���g�i|:^�B�    @?+�IL�K��x�N�w�ލ�?�<  `P	� 
�r���J�Ie��^�    � ��Q�g���Xq��o�� 0��  �?��O��P�S�t���v    `@�$>h��ɖw�ngg'���bzz:  `	� x�n7=zpR�z�t�z;    0X>l�c���]�/-�q�F��  Dw  �_����t:'��Ɇ�v    `��$�5�1���6+++������  �� ��w��퀓��
q�z;    0���˱�lǞw�q������  �� ������V+���D#     U�D|8R�ٍ���y��q  � � 0в��^�J'3Z.��z9     �t�t�������������>  $w  ���~,--�ԯ&�    0�V��x���6�o�� 0p�  �o��6�]�4�L��~�f�    Wk�Xh�Yq�^�x�f3�F  ��� 0��ݻpR�Zo    �H�D\k��w�q�ƍ��o  �� ��������'�(b�z;    0dVܷ�����277  0H�  ��ׯG��='�	G�    �'�V�G*1��p�N���ߏ�>�,  `� 8�v;���N�^*�T�     �h�V����س��[ܾ}[� ��� 0p����;��n�I��x-�$	    �a����(���n�Q^�x�f3'� ���  �{���D�X���J     �j�x�lǾw��ƍ��7�  �;�;  eqq1���N�Ӊz�n    �]!M�z)��G���  w  ���ף׳@���4���    ������9B�Ӊ����g�}  ���  �v�KKK'�w��H��    @>�w��Iӊ;G�}��� ��'p ``ܸq#��n�q*�4��     ȓ�x�jG׈;Gx��E4��h4  �J� �����	8�O�k��   ��)�IL�J�p�lP�o�	  �Ww  ���b�Z���d/p��T     �>����~t{f�9���\  @?� 0�_�p��׭�    ����\��b��8L�Ӊ����g�}  Џ�  ��v�KKK��^�|h�    ȹk�R,��aÝ�ܾ}[� @�� ��nܸ�n7�8�ף�Zo    �RH�J��Z{���؈f��F#  ��� �{333�)�I|d�    ��G�J,����s�^�w00��7�  ��;  }�ٳg���p�Gk��    �W���T�+�V�9ܓ'O  ��� ���������$I�[o    xՇ����#������\|��'  �D� @��v����p��F%*�4     �?�b��b�h�����w  ��� ��u����t:��d�     ��Ñr�X�s�������45" @�� з��8ΥZ)�B     ��r!�B4���^�w�܉/��"  �_� �K�v;�����w���    ��Z�3�������  ��;  }��o�=X��-c�R
     �6U)�\!�ݎ��l\�F#  �� �K���8�'�     ��$�F%f7v��%��_�5  �� �;ϟ?�V��6�b!��+    ��֊1��D������w  ��� �����瓱j     p2�$��z)�������ӧO�ڵk  �� ����ɓ��)�IL7�     �q�Q��V;�F�9ĭ[��  ��;  }eff�`%�棱Z�$     8�l<�r��Z�������v���i  ��$p ��d� �6�1��Xo    x���X�ޏ^ό;?���w�ލ�?�<  �}� �7��v������H%J�1     �VLc�\������	� �w  ��_���1���Z     ��>l��jss3Z�V���  ��E� @߸w�^��\iT�V*     �n�\���][�N����׿�W_}  �� �kkk����6��    �Ƶz9^���c�;  �� �������h�c�0     g�R��B��n��vwwcii)���  �u  }a~~>�m>�     g#I"��J1���[�n	� xo�  �w>�v�p�R!�+�;    �Y����Is7����y��Yt��H�4  �	� x����p�i     ��b�ĥj)V��^��t�>��  ��&p ���?�8JvL���     ��Z�,p�Pw��� �^� x�~��ǃ8ʕz%*G�    ��F1��r!6۞��s���CEi�=  K� �{������G��     ��L�Jw������~���  \$�;  �M�����p��r1�*n[     ��T�s[���t^u��=�;  N) �{s�Ν��8�G��     �|%I��Z���j}}=����X� pq|� ����R*�q�!p    ���R<i�F�.����|��  E� �{��}����Ñj�I     p�i���X��x�����  \(�;  ��_�������p��k�6j�    �"]k��ass3��v���  �� p མ��	8��z%*�4     �8�b��Bl�;/e�E�oߎ��
  �w  .\����ŋ��|4f�    �}�����ѣGw  .�� �w��̓�8�H��R     p�j���j�n��R�ٌ����V�  p��  \���Z     �~$���K1���R6\t�֭���/  Λ� ��j�bcc#�0�4���r     ��\��b~k7�ʫfgg�  \�;  ��͛G�n���$    ��SJ��,cuw?ढ़����܌���  ��$p �B=|�0�(�Fk    �����yU�׋۷o�W_}  p��  \�lգ�jf�Z�F�     ���BTi�t�/���	� 8ww  .̍7�=�0�F�    @��R+��V;ढ़��X__����  ��"p ��<~�8�0�4���r     �?���1�l��^u�֭��o  ΋� ����������Q�B�     ���&1Y.���~�K  �I� ���y�f�Q��V    ��3�(�������a����  �� p �B<y�$�0�R�K�     ����Q-����dz�^ܾ};����  �� p ��mmmE��
8̵��     ��J�s[퀗�>}  p^�  �����/�)�iL��    @��Z/�|��^�����������  ��&p ������F%
I     ��R��d����/ݹs'��_�%  �	� 8WقG��8̵�j     ���e�;?3??/p �\� 8W�n݊�3K9�D��R!     ���BTi�t��V�u0tT�� �l	� 8W>8̵�    ɕZ1���l��~�?��  gI� ����ߏ����ו�$.�+    ��Z/�|�n�G�	� 8sw  �͝;w��uT)o�nT#M    ����L���������<<*%H  ��. 87���8���v    �At�^��3?��c����}  �Y� p.�������׍��     �g�R<Xr���2<� p�T%  ��l�=���u�T    �����\+��f; ���~�N(M�  �� p �\d�Q��W�     `p]��^�w������&  �,� 8Ϟ=x�T�|pt-     ��^L�־�\�333w  Ό� �37;;�N'�u�#�     `�e+�����  ��"p ��ݹs'�u�4�K�R     0�.�J�xk7z���᣹����O  ~)�;  gnqq1�uӍj�I     �R��D�k����w�
� 8w  ����R����n�Q	     �ǕZI��O�={  p�  ��[�n��^*�h��    �0����&���t:��!����  �_Ba ��ZXXx�#�     `��IS�b,m;ٕ���?� ���  ��f�;;;�J�$�6*    ��R+	��ɳg�  ~)�;  g��x�D��B     ��r!��4Z�݀l��jE�^  xWw  ���Ǐ^��H5     ^�k�x����w�^��?�c  ��� p&��n������&q�^     ����We�Hw  ~	�;  g������^u�^�4I    ��UN���c}w?�ŋ�Hi�  ��;  g";n^7=R	     �_��.p'�"���ŧ�~  �.�  ������WU�i�WJ    ��"M"�{�o�߿/p ��	� �����boo/�UW���    �$1Y)��+�D,//  �+�;  ���۷���W]i�    ��r�$p�@�ݎ���  8-�;  ����|���B���n     ��x��4���Q"~�����/  NKq �/��v8�UW��    �N�$1Y)���^��'O�  ��;  ��ݻw�׳���	�    ��r�$p������PR��  �!p ����	x�h��b!     ȟ�r!Ji{]�8y�$=z�(~��_  ��� �_dyy9�UW���    ��R�K-+�Dܿ_� ��	� xg+++�����;    @�MUKw<�<  ��  ����.�U�RT
i     �_c������N7ȷ���X[[����  ��� ��^u�z;     s�R��-�;w�ލ���*  ��  ��v��f3�$I�J�     p�V���� �I  ��� �w����G��xi�R�r!     h�
Q-$���.!�Z�V���G�(S �d|s ��<x� �UW�     �����x�l��&�������  ��� �NVWW^J����;     ��r�(p����� �� pjϟ?�N��ҥj9Ji     �R�X�z��=��nmm-  ��  �������    8�TE�N���^lmm���H  �q�  ����B�Ki��T�     �Z9��333�?�!  �8w  N������F�K�b�$     �u�B�b��n�oO�<� p"w  Ne~~� r����+     G���e�=�^�x  pw  N�޽{�ʎ�    ��\���=�:�N<�<���  �F� ��,--�4^-E��     �Q*D���n�	�y�)	� 8�� ��v��l6^�R�     �R�O�V��nqq1  �8w  N,[���z/M��     Ǚ�܉���:TJS�� p4�;  '������F+Ũ=�    �x��4Ji{]C:y�)-,,��  p�;  '�����e��     �P�$q�Z��������  ��� ����9����J     �IMV
��
rnyy9  �m�  ��ݻw���L��F�T     8��r1
I�r��j���~��%  �"  '2;;�ҕF5     �4�$b�R��;�A�=|�0~���  F� ������4U+     ��T�$p�`XI� �Q�  kcc#���2�Bc�;     �7Q)F�Dt{A�=�<  �(w  �����G��I3��r�     �.��}�\��]+�y�+���D�Z  x�� �c����t�^	     xW��{�e�J333��_  �N� ��^�x�)�i�WJ     �j�Z�d#�ٱ��,	� 8�� ��Z\\�N�����"I     �Y)Mb�\����y���  p�;  o�	/M�+     ��d�(pϹl`��lF��  x�� ����!��g��    �/5Q)��f�c�^/�߿���  �*u
  o���������     �T�X�j!��N7ȯ���;  o� p��������L��     ge�R����=ϲwQ  �:�;  G�w�^�Kw     ��d�K�� ������nG��  �G� ���<y��Ҩ�
     ge�\�B�D�����Ç���.  �%�;  GZ[[�L�+     g)M�-b}w?ȯ��9�;  ?#p �P�V��XH�\��     ��d�(p�9�K  �N� ���ݻ�I�����    ��7^.�����n7�4  �� 8���|@f�Z�B�     ��j1�Z���� �z�^<~�8~��_  d�  �����K�r     �y�(������� ��;  o��ۋ����̥Z)     ༌��x����J  �Kw  �p����L�T88     ��d��ͽ����|��ގn�i�  � xCv$d�j�     ��$��������bqq1>���   �;  oX^^�L�J     �m���	r�ѣGw  � ������H($I�W�     ���#��_nF�P��   /	� ����كc ![oO��    p�j�R$흿������V  @F� ��<|�0 s�V     �(#�$��^$�Wr);e����155  �� ��YZZ
�LV�     \��F�Zތ��� �<x p @� ��5�̀Z��b     pQ��5��pA��c��  �� �������0Q+     \�4Ib�T���ݨT*A�lnn  � �Iv�#d&+w     .��1��E\�z5ȟ�����ىj�  �� ��<{�, I���
�    �xY�~s�iLMME�P�gvv6~���  �%p �'/^�)�TH     .�d��b!677cbb"ȟ���; @�	� 8�����`�    ��%;etz|$��������Z  �ow  <z�( #p    �}�6>�W�c{{;j�Z�/��;  �&p ����\@�$1^�    ��d��{u�݃����   ��  X^^���&     ��h�#�r4���t:Q(�|���� �� �[[[U��     �L�������܌��� _�={  �� ��P`R�    @�9�766�9���  �� �x��a�z� �
I��;     �_�����ۋ����jA~���F�ۍ4M ��� �����R$     �_�T��F-֚�+���y��i|��G @�� ���Հ���v     �����A��l6���D�P�cnnN� �Sw  ��jL
�    �#�&F㇅���z���A~���  �$p ȹgϞE���RH�^r{     @��:6i�D�׋���{�lmm  ��` ȹ��ـ	��     ��b!���z,o4coo/����V��������(�� @�� rnqq1`�"p    ��d+�Y���V����5����  �E� �skkk�    �GW�?���lF�ӉB�����  ��  9��vcww7ȷb�D��     ��+��H�$z������A>���  �#p ȱ�X��a0�6^)�     �~S.b�^�������i�Z @�� rl~~>`�Z
     �WW�?�{{{����j5~�i��j���h  �w �{��Y�X�m     ���X#~|����Y�,pϏ�D�/��"  �% @�e�ɷB��H�m     ������~��ڊ˗/G�$��3� �?J ��ʎt̎�$�F+�H�      ���ʥ�Vbsg����G�ٌ���`����  �"p ȩ'O�D���m�Z
     �wW�?��Z�{>���  �"p ȩ,p���[     ��ձF<x���ϭV+:�N
�`�e��Y�^�V �|P�  ����r�o�߮��w     �ߕ�7�ڳ����`�e'����o~�   �  9�����h��4	     �wc�J�ʥ�n�����=?�  9"p ȩ��N�m��v     ��qe������s�ݎ��ݨT*�p[[[  �C� �C����9�o�R     ���2���=���܇_��  �C� �Csssc�;     �cz|�ϲ�}jj*�$	����^t��H�4  ~w �Z\\�^*D)��    ��1Q�F�X��~�ϲ��jE������R\�v-  ~w �Z__�m�j�    �����_m�����>�V���o~~^� �w �j6�A����
     0x.���ܳ��N'
�B0�VWW �|P�  ������C^�m�b�    ���-�fkk+��ǃᵱ�  ��  gfgg����UL���     �A35R?����M������  �A� �3O�>�m�\�$I     M�X��Z%6�;g�s�ݎr��l�i}}=&&& ��&p ș�ϟ�6Z)     �K#�7�L��>55���y�; @� rfkk+ȷ���      ���z<Z^{�����}�-//  �O� �#�n��xN�m��6     ��55R?�������ىj��/^  �O� �#O�<�^��W��F��     �K#�H�$�����V��ë�j  �O� �#Y�N��VJ     �,��'�x��f��/_�S�ӱ� �w �YYY	�m��     ��wy�~h������Q�Ղᴰ����� ��n ȑ��� ��*n     |S������d+��ᵼ�,p r� �Ɏl$�FJn     |S#�#��/_�$I�ᳶ�  7u @N�������k�\�B�a>     �o�V�r������v��j���h�'�  7�; @N<}�4ȷъ��     �l����桿�"h��p���  ���  '�|-��    ��x[��l6���E�8�t�d�����r9  N
 ��X]]�m�R
     S��#���Y�>22������O ��$p ����moIz���|�dI����K���Z ȓY�=c�߻�lk3�̮mI�DuU� �)e��BT������A��� �:      ?\�}������� �M� P��b��b2��    ���hg�qܯ7_����H۶QUU��_�5  ȗ� � ���v��u>��    ���?�}3p���qA^�u~  �r (�O?���|�?     ��>��~���w!��=?��2  ȗ� � w�Fu     @n���{�E4Mu�<'���ݫ��   ?w �|��1(W5�\�    @���揾���>޽{�c��?<�ۿ�[  ��; @>����ۻ�     rs6�d4��v������	�3���?� 2%p (�r��uf�    ��]�g��͗o�{���mۨ�*ȇ� �%p �\w`�^��r�O|�     _Wg������������˗   OJ ��Y��|�k?     �z6{�=���V�   OJ �����wP��Q     ���'��"��}� ����&㪪 ��� 2g��l���Q�`    �|]ΦQ����|O�w����Y��O�>ŏ?�  �E� ��ϟ?庘�     rVU���O����w�w/p��_��W�; @��  ��k)���     ����ٓ�n�}0y�� ȏ�  s��:(��H�    @���G�Ӷm�V���/i���	  �#p ������	庘�     r���i�z��D����  ȏ�  c��_�r�*&u     ����E������?y�n� @~�  ���cP��q     P�Q]��tw��w��4����t:���d���b8�@ �ķ; ��}��9(����}     �q=�=�w�w�{�������  �x �ؗ/_�r	�    (���,��G���>|� p ȏ�  c��"(�|X     ��j>{����ml6���A�nn��  �"p �Xw8K��#�;     �x7�<��݊��=n4 ȏ�  S���~��4�QW�     �R\L'QU�h�ǟ�t����u�>7 �G� ���~�I�^�ٰ
     (I��O�q�\?���z��.�C�L��h ��� 2���?�:��    @y.��'�n����2H[�4ѶmT�� �\�^  2�믿��     �Ҽ�M��?o����b!p�D�\�Ç @�  �����5�    (��|���.�����1��}��Q� ��; @����5��    @y�=#p���.r���A�~��   � �L���L�j��    �Ҽ�Mٻx�)����p�1 @^�  j�6��	�t6�5    �2�*�&��[m��~7���� �� @�>~���e�3�     �z7�>9p��v��lb<�r�1 @^�  ��矃r�-�    P���4�߯�O~��-pO[��
  �C� ��_~�%(�|T     ��r6y�������*HWw����]���  �� d����A��F��    P�w��޿\.�mۨ*2)�n8� �A� ������Lê�q�     �r]�=/p�t+���}��)��?�#  H��  C��*(�|$n    �l����x����?#pO���M  ��; @��ۧؒ�����     p9�>;p'm>C �|�_  2ӭ�����L�Q     P���$~�����o�&��uL&� M�� @�  ����SP���     �b6}��t��tm6�   w �����A�f�*     �t�����>����4u+�  �A� ������\ӡw     ��=�}�^?D�u�=U�
�|>  �&p ����]P�I]E5     ��l2��`���Y?��A�����  �� dF�^��Ȣ     t�A��x��ͳ~n�\
��������  �M� ���j�i6�    �o.��g�݂;麽�  �'p ��f�Z�1V     ���lq�i���Y�x<��c �<� 2���2M-�    ��:��/�K�{�,� �A� ���j��>(�l$p    ��\L'�\I_^^�q�1 @�  ��_�r�,�    ��:��w�ݠ�`0Ҳ�n ��	� 2"p/װ���r�     ������.n_��1�N��4M  �O� ��ϟ?e���      ��hX��o�����s��.pO�b���|  �K� ������L�Z�     ��|6���ų��������t7� �&p �Hw�J�f�:     �?��N����z���m��̤�������� �t	� 2�]�I��#�;     �����������Z�,�'�˗/ @��  �l6A�,�    �?��M��nXH������   mw ��4M�if�     ������}�Xć����  }w �Lt�d�m��b\     ��������n��ƅ���LJ��u  �6�; @&>~��i:�b0�    �?��GQWU4�uk����A:��m  �6�; @&>��iRW     |��d���V���q�1 @��  �����4
�    �[f����b�e���f���x  �I� ������L��     ����C��n��6F�Q�������� �4	� 2�Z��2Yp    �o����ӗ˥�=1���w ��	� 2��R��Ђ;     |���nd�ݻwA:�E  �.�; @&6�MP�qm�     �e>9~������  �� db��e��    �������n��e6��� �6߼ 2��R�z0�a5     ���&��j����� �� @��  �h�6(�dX     �m�aú�]s����r)pO�z�  �%p �@w�����L�U      �7��vyx�l<-n> H��  777A�Ƶ�     s6�o6�h�&��ͪ)� �M� ����۠L�;     <j6�;��u�����?F   ]w ����e�    ������r)pO�~���m��<G H��  �rM�f    �1g��ѿc�Z鸿�����   =w �,��L�a     �����/����e��`�����  Qw �X)פ��     �����{�w�df�Y�_�|	  �$p Ȁ��L�`ue%     s69~��#pO���]  �&�; @v�]P���z;     <Ũ�^ۦ9��,�˸���o�X  i� d`����w     x��x��q��[u�� H��  m���    ��M�]&�>�w���X��1�L�~�>'  �$p H\���4�     <�t�2��r��'��  �� $���&(Ӹ�     x���e2��j��v�  �$p H���]P&�     �t/��^���s2 @��  �[,A���*     ����F/�{v���k8�����  ]�i $�5���     O�R�n�]��o��>  H�o�  ���k\�     <�K��󙳳���,� ��78 ��	��e�     ���鿻�����
  �"p H��2ՃA�w     x��^p�����  Aw ��	��4���     ���0�jm�?�w����l61����  i� $�;<�<�     �y&�a,7��]����ߺw  �#p H�v�2���eTYp    �皎^.p���/..���� �&�; @⚦	�3V     <O���t�u+�  �G� ���n�gT	�    �&/�o6�h�6*g���}F  �G� ������k��     �\/������t���  Mw ��5M�gT     x���W����Ƕ�m  ��; @�,��iT�    �^:p_��A�v�   =w ���V�\�     �y&���N	� �$p H�b��T,�    �s��/; ��M�Dm����  i� $���>(Ө�    �s�^!D�V���΂�i�6  H��  a��2(�`0�Z�     �6�|*�^��=��� ��� �X,����     p�q]����w�ɂ; @��  	��^�Z�     뇛R_r�[��o��&��q  ��; @�V�UP�a���2     P�Q]�f׼��k���U�u�?�`��  -w ��u��gX�p    �C�������l6������  �!p H�n��c�     7z����z-p�)�Q  �� $L�^�ڀ;     �[pi]�N?m��   -w ���m�gd�     6~�w+��� H��  a��44�     �^'p���18���  �� $�i��<u�p     5z��N�O&��_F �G� ���m��*     �Ì�����k�{Yp H��  a'�Tp    ����;�#p H��  a��4��     {�w��` @z�  	��iX�p    �C�ւ�����  �� $L�^&�     p��+-�����n�1���h�&  H��  a�A)��     ��R���V���"p H��  a�2��    �p�+ޔ��l�~� �G� �0�{y�AT�;     jT�^��-��/w ���  !��    �8��Ҷm  ��; @���8���     �y��}��=,��u��  =w �D��L��     �RW��6$��n�=���  i� $j�Z���     p�nPf�J��f���t�w ��� ��R�     p���b�J�g8�"p H��  QG�T�p    ���A�_�wo��   'p H���LU      Ǫ��;q��_��}  ��; @������     G{��}��E۶QUfk���,  H��  Q��(�w     8ְ~���*�L&  <��  Q�&�$p    ��_y]}���{b��
 @r�  ����Ay*g�     p���;��� @z�  �j�&(Ome     �&p ��� @B*�;     �~�+S��m   �� $ʂ{�*};     m���]���c`��ڶ��?s  ^��  Qݡ(��     ǫO�(�E��$x{w ��� %p/Sm�     �Vׯ;o6�{Ot�;  �� $�i��<�    �x��4�;�`8
  -w �D9�+��     �w�=��v��( ��� %p/���;     �7�Zp��; @Z�  �j�6(��     �w�A��� @Z�  ���^*�;     ��{��E��(x[�� �E� �(Ke:Ţ     �:�y���<W H��  Q�&�$o    ��2p��5M  �C� �(�;     @�	����; @Z�  �rW�S-�     @�':o��v��3 ��; @��     ��N�[pi �t� e�     ����� @Z�  ���^��DW�    @�N4��Vw��u]o�s5 ��� � �T>w     8����2݊���mYp H��  Q�2Yp    ��:p�N���� �E�       @QN9'��  ��	� UUU      �|Չ�y[u]  �� $�Wg���     �6��p @Z�  ��     �����y� ��; @�,M��,     �7�6Mm�z���  �!p       �Wԭ�O&�   'p H���2���      �Ӟ��]����C� @J|{ H���Lw     H�n�ގ�j  i� @BZ�;     �����&  ��� $��D�ڶ     �8��1Ղ�۪�:  H��  Q�2�-�    ��N}�.p[w ��� 5��w     8���� H��  Q��Դm      �i���m�>�<�y��  �"p H���2�-�    @����x��?,  H��  Q��tq��e      Go1(#p;áD
  %�� $���,Mӄ�     ��{2]��۰� ��; @�,���;�~�E     ��[-�  �� $��Dy��     p��8m���n4�s5 ��� � �<]��
�    �h��a<  =w �Duk���7     ��V�  �%p HT]�AY,�    @��  �4w �DUU��;�v�&     �-eڶ}xy�  �'p H�p�\i���     ���jP�������   -�( �D�F���A{��w     H�����  �� $j2��x���f׶     gۼ�y{�sZw ��� %p/�o�w     8^�
�KQUU  ��; @�\_Y��ܛf     �q��� ��; @�,���w�     p�]�6�2�ӳ� ��; @�������~oѻw     x9��Q�u  ��; @��M���}��    �X����v���x� ��;  $��;     ���}�r�'p H��  a�� ���9����	��     p����w�{]��i��  =w ��u�������     �X����� H��  a݂;e�-pߺ�     ��ց;�3ʣ  R� @ºw������b?     m��K!p H�op  	s�b~�ݴ�      ��{�A��n���i  �� $̂{��[p    �c�堌�Ӳ� ���  fq��?�~�+S     o9(#p?��h  �E� �0�{����,�    �Q���]�~Zw ��� &p/����     p��ݿ����I��( ��� �0�{������     R�Xp/�x<  �"p H���������òL]     x>�{YF�Q  ��; @�\�X�<�����+�=     bۼm���t�6��1�S� �G �0W*��������Wy     8�f�{��g���Nc:�  i�M  a��$��?�]w��    �C���{g��	�Od6�  i�M  a'��]Qڽ~��     �����i  �� $́\��v�����;     ��C2��QUU  ��; @�\������C��֡7     �C2_;���u�;  �� $���,�����V]     �`������Ӱ� �&�; @���σ�}u�}'p    �C�a��1fsu]  �� $l:�y�z����     ��m�����OC� �&�; @ºk��C�|}�][p    ���aHƳ���F @z�  �A����?�߶�-    ��m,�C� �&�; @��F𜭯po-�    ��6۷_p�l�4�  i� $n8�v�����}-p    ��m[��� @z�  ��w�e�     ^�~���9���4&�I  �5 @�\����povw     8Ķ�GX.p?�; @��  �����M�~�`     ��mv�苦i������f�   =w �č�� _�Zp�O��|�    ���4�YN��_�t:  ң� H��=o���;     <W�ܿ���3�� ��(b  7�L�|}�p{�k�<     ����l���uvv  �G� ���l��{��mf      �M�כ�	^�t:  �#p H��=_�������l     x��?���_�`0��� ��� 'p����[V�    ���tC���uu�;  i� $n>�y����҂;     <�J�^��  �� $�ݻwA����7�me�     �m%p/�p(� H�or  ���fW,~/�&M�;�^	�    ��V�b� �� @�+��	����m      ϳ���|�x��L& @��  �(���n����     ����c��g5]�����i  �&�; @F�Q��� /�_p�    �s���^E�m۟�>G��<  H��  ��8���ٛ���n㡯�     �}��[pUggg @��0  ��fA~;����     �4��� ҥ� ��t:�����r��w��     �dݳ��m���\\\  i� d`>��y�`�o�     �g��ryy  �I� �yz�`{��     �4�r��� @��  ��鱃��F�     Oշ����\9\UU @��  p�b�]p���      ��o7�Zp=w ��	� 2��ݻ ?��[�;     <U����g4  �� d�[��^�����{��f     ���x3j�l������ @��  �����}��    �S�q8Ɗ��L& @��  ��(v��-�p���`a��     ��vMۿ�\��:��i  �.�; @&�C_�r�ءvw���b2��    ��,��[o︝�u���   ]J �L�f������Ֆ��F�     ���魨�_���y  �.% @&&�I�����ϭ�     ��,6�\p���; @��  �p�b~�r���+U    �O�=�۶^���e  �.�; @&,Q�婋-��^�
     }�<�,ggg @��  �x��]P�;�     �����?u���QUU  �.�; @&�����,zz�*     ���r�r( ���F �����?,RX���S?�Ū��3     �ݙ�b����s��7� ��	� 2�]�ؽ��	���+U    �/V�]�B�b�f�   mw ��tW.
����w�ӑ��     �5�M?��;�_�|>  Ҧ� ��d2��z��9�݊��     �n��o���;??  Ҧ� �H�Hq{{��;���     ����+�/���2  H��  #)���w     ���%y��}  �6�; @F...��,�     �M���_���u  �6�; @Fؕ��     |���PL)�ATU  �M� �W.��9�-�    ������[pY��(  H��  #WWW�C�r�^     �Ϻg&��.(�x<  �'p �Hw�b�j�&H۳���h�6jWn    �tg�mk���$  H��  3�Ջ��t1�b����C[     ��/�~߂�Vޗuvv  �O� ��n�b�Ze���     �G��MP����   }w ����󸹹	���Ŗ/�u�u      �c��,��� @��  �q�b��~@     o��yY��� ��	� 2��ݻ }-�     p��D�YpY�׮� ȁ�  3�)�0��~4     ������y9UU=�  H��  3>|�sg�     �`���v�D�=w��o��:  ȃ�  3�������,ˮmc���l<
      ��O�/g<  y� d����ߋ$|�!��A��     ��n�	�1�� �<� 24�Lb�Xe�[��O��     Hc���sqq  �A� ��n�B�����-�     �oR87?�y _wuu  �A� ��n��ӧOAY,�     ���n>�?��c  ��; @�����/�KP���*     ���[[p/ɇ �<� 2��?i;�@ۂ;     �ݮmc��e��*�C @.|� �п�˿�Yow��51�     %�[�1
c��e���   w ������~����n����<     �dw�MP��t  �C� ��n�b�Nc���#p    ��<��݂��8??  �!p ��l6��v�
     (���yyI��� �|� 2uvv�?�t�b���5     ��}������Ç   w �LuK��_�����2     �t����?  �� d�A^�n����_     (�r����	��=��� @>�  ��ӟ����@}׶q����t     P���:Ra��x��(  ȋ�  S�����ݚ7e�Y,�     �f�
�1{& ��; @Ɔ�al�� =�,�t�~     P��e:���㝟� ��ٻ���3��/ �)J")q�,K�▇�޻�\��]՗�T�S��$�'�<E�e��'� �igQ'qEX�y��w�<�������� ������sh�2     9��W������d  �_�  }l||<vww�lJ���v�����j     @^m[pϕ�g�  �E� �ǒŊ�ϟ�����w     ��lF� ;��
܏off&  �/w �>f�"ۊ�b�Z�#���f��clh0      O�*��I��x��'  ��� ������u�Ֆ��}�;     ��]�V�n��xJ���H  �	� ���=ێs���ۏS     y��d���x��� ��#p �c�bE�\�l6��9�Q{�R     ț�j-����񌏏  �G� ��FGG�\.�s��=cO�    �Iض��+gΜ	  ��� ��MNN
�3�8G�-�     �L�Պ��zd������� ��#p �sgϞ��O��s�gI�덨5�1<P
     ȃ�j-��vd�q������  ��� ����l�M�]nٮTc���     �<��ۏ,��~<� 066  ��; @�[XX�鸇�M�;     9��ųD�~<CCC @� �����(�J�l6�l9��     �"kw�d��w7>>  �'�; @���D�R	�币�Fe/      /6-�����T  П�  9p��)�{w�e�\�V�Er     �\����Fd���x��� ��$p ȁ3g����r�-�=l7[���ۏ���     �~�����q�n�nnn.  �Ow ��������:Ȗ�Xn٨T�     ������]��nbb"  �Ow �XXX��$ۛ彈ٳ     �l��Yc���  �K� �ɂEK��� ;N$p��b     �fe/�Ƃ��  ���  '���c?{�%yv�-����    �(�V��D�XpwSSS @�� �D��.pϖ�8l���;��ؐ�:    �O�k�Y|�V��� ��%p ȉd�buu5Ȏ�:lo��b���     �~��W�,������  �	� rbff&��� ;
��:�j,�    �S�l�R)8����s��  �K� �.\����+{     �j��Yd���  �M� ���Ӈ��V�dC�@�����c�:ɂ;     ��䆾���;���݌��  �M� �#CCC������J���f�X���~-�V��    �/���7�,������  ��	� rdllL��1'�'�5��j�L�     ����^d���ݜ;w.  �ow �9s�Llll�qR����/p    ��l�ewاT*G777  �7�; @��?>�߿d�I�ɂ;     ���޿���Gg� ��	� r�ҥK����qR��z�     �o�L����y3<<� @� rdbb���f�d�I.�7[�(9�    �'���_oD���ͩS� ��'p ș���(��A6�ԁ��j�F�3��     �`m7���&�D�ٳg ��'p ș��)�{�����nY�    @�X/�EVYp7��� @�� ����L<~�8ȆB�pb���nv�     ���|��]�Ʌ ��'p ș������d�I��v��T+     ��V���jd����J�R  �O� �3�����v;H��<p��עVo��?     �m[��h�Z�U��  �A� �3��tdd$��쮚��I��v+�p�t     @����E�%k����T  �w �����g��     ^�^�D�Yp?����  � p ȡ���XYY	��\�2�h     �5��  ��  �����޽{A�ub�     ���l�N�Y&p?�B��N�
  �A� �CKKKAv$G�f�y"�V�ވ��ZL�     d�zy/��vd���hFFF ��� ������O�^��$���NE�    @f���E�	܏���� @~� rj||<�����+�'��m����ٳ     Y�.pϝ���   ?�  9u��Y�{F���{u�     �U�l����[XX  �C� �S.\��w҇����l��t���     �i{�ß,���w �|�  �.]���y�~�ћ�vlU����X     @���f{�=a��h���N��  �M� �S���V��['����    ��Y/��&�N �|� ����X��� �:q�^�.�{s3     Y�����5�Gs���   _�  9v���{t��͕m��    ȖV��sgnn.  ��; @�%�G��։Cw�v���852     �k�{�l�#��o�P(���R  �/w ��v�Z��w�ҭS����S#��     ��uR�����K�  ���  �&&&���f3H�d�$�i�Ov�fe{7��
�    Ȇd�������d  �?w ������ ݒcw��8�_s�O�n     ���zy/��������  �#p ȹ���{t"p��ۏZ���     ����~4��EZ��ۻx�b  �?w ��[\\�����֩c���n,��
     H�~y��X,���
���P  �#p ȹ+W�į�� �:u�N��    �v�;��������h  �Ow ��:�988ҫs���x    @[�����ӧ �|� �������W���h4[1P�*     �S�E���``@����� �|� ������\�ޭv;Vw�175     �F�;������]�t)  �'�� ��/ƽ{����䓥+�w     �ke��B��v��EN�:  �O�  ���b
�h��A:u�ོ�?�7     ��U�{�  ��S3  Q,ctt4����tJ�u�?BX۩D�Պ�_~     H��A=v�k�/�o��ٳ @~�� ����)�{�%�q6��u�VlV�1=a    �tY��WH�ogaa!  �/�� 8t�x��i�^�ѻ�{be�,p     uVv*�O�1~���b  �_w  ]�z5���?��ɣ��v9n/�     H��>
ܓ!�B�������  �%p ��ٳg�X,F��
ҩ�ϖ&�{��vX     5j�fl��G��䝿�LLL  ��3  s�ԩ���	ҩ���F������x     @<��9g���3==  �O�  �M��.pO�N��m�
�    H��[��'��s�ҥ   �|r �o�~ҩ���[����     i�|[��7�B!fff �|�� ���r�J����{�N�>|/o�F�ՊR�     �K��A��k�O�lxx8���  �=�� �������a��_�~�t��v�ݑ_���_we�sS     ��lk7������;w.  �'g  ~fjj*����t*�J�h4:��?���    �sϷ��o�lii)  �'g  ~faaA��b�񻣁���_��B     @/=߶��GW�\	  �� ��y����C�N�>~o��Q�7bx�     ��ʋ[u?�����!��  8�S!  ?399��p�]�T���n�Wq.M�	     ��[������M  ��O�  ����ӱ���O7��6w�     ��3�{.���  $|z �%sss���J�އ_     ��v;Vw+�o�7�z�j  @B� �K�]�_|�E�>��w����b|x(     ��Vw*�h�����,��cll,   !p �%�ϟ�b��V����[O�>�܉�     ��y��2*p�ӧO  ��� �W������� }�Ƚ�ht��H�@�    �m�;��G�7�p�B  �_	� x�d�]��N�ܟm�     tS�ٌ��^��B�еZ���ի  ��3  ������ }����������FlV�qf|4     ��o���jG���Y�T����  ���	 �WZ\\<\i��u�:�'+�w     �ey��(������  ��� �W*���r�?��Y֭����v�^<     �O�v�	���  O� �k����S�[���N%��f�J     ��S���_~����ͮ\�  ���  �֥K����ҥ[��f�϶v�⹩     �Nz�ٟ��	���%/
���  �=�;  �u�������v;H�B��R)��f��'�w     :N��O���  �H� �k���HT�� ]�7���oG�     �F�����W�כ��	  �Gw  �hzz:=z�K��j���>Ճzl���쩱     �Nx���>}M6��'/��j�/_  �Gw  �hiiI��B�\{y��#p    �c�;t����zI����  ���  �����㷿�m��t9%��ŗny��\�     �	϶�y422�b1  �	� x��8<<���Azt3p_ݭD�ь�R     �IڬT�R�G�������  ^E� �/J�>ң��{�ޟ��_�=     p��l��z{B��zW�^  x�;  �������)�JQ(��nx��#p    ��=������5Y�|Ǳ��  �*>E ��nܸ���o�S�v�՗�����^ɂ{��?98    �I8h4c}w/���W;u�T  ��� �E�b1��ǣ\.�����Vo���^�L�     ��d�����:�k��/���  x�;  o%94~��wAzt{�%Yq�    pR����Yo��ׯ  ��� ��r��5�{�t�0�xc;>�<     p\�v;�m�F?
^��ڟ;w.  �u�  ���/F�X�V��C����^��bl�A    ��Y/��~��L��j���  o"p �%ǭ�� �P(��t˓͝�qa:     �8�n��z{B��jKKK  o"p �-,,�S$�ۓȽ^�w��|��%p    �؞llG���K�Yq���  �7� ��n޼_~�e��q�����͝�7�1X*     ��J� 6*��g����5���  ��'i  ������1��h�����f��6w���T     ��x�����CCC��Ξ=  �K�  ə3gbuu5H�^<o�����    �w�h}+�����.^�  �K�  Irx��G/���[�l��T,     �~���{���/+
q���  �_"p �Hnݺ����t�E�~�h��v9��L     ���h�����/���  �̧F  �d||�� Y�Ղ�K�N�cp����������    �#{��yЋ������	  xw  �lzz:�<y�Cr$�zྺ����a`     o��L^ݍ~����/�r�J  ��� pd�/_��Hr$�V�]�=��X�݋���     ���dc'��v��������ii)  �m� 8�7n���v����W+0�6�     ��Gۑ��_6>>�b1  �m� 8�dydtt4������ա�ǵ��立     ���nǳ����/���  x[w  ����\ܿ?�^����جT���h     ��<�܉z�y p�{�  ��  ��[�n	�S"yҳT*E�_$+�w     ~���ȋ^ӤU����L  ��� �Nb`` �F�{�L�Z������Vܽ4     �:�v;o�D
����ٳ  G!p ��%ɕ�����5�^j��kqjd8     �UVv*Q��c0G���+W�  �� �w�$���˃y��~{�|     ��<Zߎ����ڵk  G!p ��ݾ};~���>-Jo�4p_�    �z�7�"/���x��N�:�$  ��'H  ����`���G�\z+�wQ(z���T�zP�ѡ�     ���QދJ�y!p�����  ��� p,��7������j����IT�pm3n��     ��V7#Oz��j�$�<�n�
  8*�;  �r���{J$+��?��    xُ�ۑɝ�X,/�J����
  8*�;  �2==}x�����hZ�rfe���A�[�    �������8/���\�  ��;  ǖ(�={�V���3�w�     $�mF�?�z�j  ��� pl׮]��@����;     ���v���y2d��o
�B\�r%  �]� 8�[�n������X<00�F�'��zy/v��19:     ����r��{s���?����b�  �.�  [r���������u�^��W6���      ��l�=��$�ᅅ��  �w�5  'biiI��Iྷ�׳����M�;    @ε��x�����z��ݼy3  �]	� 8�oߎ/��2��v�;I��K�{��Y�ƙ��      ��n��A�y"p�I�]���D  ��� p"���bpp0���u���ae#�\��(    @^=\��z{"������	  8�;  'fvv6?~�N�T:�i6{�����F|$p    ȥF��7�#o,���ƍ  �!p �ļ��{�HVb��j�~���A��Vbzb<     ȗ'��h�"O
���+���g��` ��� pb�^���o��V��i��{�'~X��    ���խțdx&	��8}�t��  ��� pb�����Tlll���{������ʂ�>    @���x��y���|Z\�x1  ��  ��d�]��[��ý�K��A=V��q~j"     ȇG����+�###���~  �q	� 8Q|�A�����v�������~��_"|��!p    ȑV7#��0<��N��f ��� p�crr2�����I���j��׶�]��B!     �o�z#�wʑ7�BA���[\\  8	w  N��˗�����I��ܓ/3�n�����    @KFOZ�������s�N  �I� p�>���{���9����w    �x��y��{|�������X  �I� p����xT*��7�rP���F3�J    @��ۏ��^�Qv���  pR�  t�ŋ㫯�
z�X,���@4���u4[�x�����     �)���a��ܹ  pR�  t�ݻw�=��{�'��|]�    Ч��v���yT*�bpp0�nhh(N�>  pR�  t����᳜���Ao$�J��뿌Xۭ��^5N��     ���v9��G��_�p�B  �I� �1q����7�tX���_Y     �˃��ȫa�����?  �$	� �>�@��Cɂ{Z$_p|ty>
�B     ��f<^ߎ�J^�ͻ������  8Iw  :&9h&��z=�O��Z�'����A��Rb�vp�L���D     ��oE�Պ���133  p��  t���\���Ao�%pO�_^�    ����W��O�T���u�V  �I� �Q�o���P�S.�#�n����C�    �u��Z��V"���G��XXX  8i�  :��ŋ100�F#�4؛�V<\ۊ�    �l{��������H����{?  �!p ��fff�ٳgA�%O�
�h�ۑ���     }����ȳa�q���  �N� �q7o���Prd��ߏ4X�.��~-&F�    �*����"��a����b1�\�  �	w  :.Y���o~�V+辡�����q��\     �MV6"ϒ�{����ӧ#w  ��;  �8ϝ;���A��mE�����.^���     ��V<Zߎ<���v�Z  @�� �7n�{$m��J� V��q~j"     Ȗ׷��lF�����͛  �"p �+n߾���o��nݕ,�F�^�������     ��lDލ��F�MMM~�   �"p �+�C�����NU��pm+>�7bx�I     �b�Z;|�3ϒA�R�y���  ��& �knݺ%p���r9=_:4[�x���/�     ِ�Ιwɽ=�
�B���{  �$p �kn޼��y4�͠��xp��ٚ�     #Z�v|��y7::yv����W{ ���  tMr𜙙��ϟݕ<�:00�F#�b{�+;嘝<     �ۏk[Q�����+#9_pOƌ  ���  t��۷�=2<<���=����    ����ȻdLfpp0�*2�r�J  @�	� ��ׯ�o~�ԅ�y���T*�H���������G    ��ک�be�y7::y6==}� @��H  ����Ǔ'O��J�Ӧ�jŃ��xa6     H�/�d�����  ��;  ]�O��O�H�MM�UZ�V�ɷ���     )�j����� ��R).^�  �w  �nii�0����Aw%�2{{{�&�{�çmgO�
     ����V��Ȼd@fhh(�jff&  �[�  ����\���Aw�.pO|�lU�    �B^^^����۷  �E� @O|���H�4z���֗bx�Q     �b�Z;|��|�R)  �E= @O\�p��)σ���{���P(D�ݎ4i���`e#�_�     ���k�����Wɫ�  �Mw  zfqq1<xtW����G�|�lU�    ��v;�_��p8&�/�vï~��  �n� �3~�a|����[�w�3�iܷ�����=}*     譇k[Q�7��^Gͣ������	  �&�;  =3==}[W�ՠ{Ҽ2����    z���������W���  �&p ������K3i\����֗bx�U     ze�Z;|q����<J�K�s�N  @��F  詏>�H��e�A:�����#m��v�_^�ۋ�    �����Z�BrS�k�>44�Ν  �6�;  =555ccc���tOr�Oc�����J��0{��     �Uo6���F�BrO/��G�+�  �w  z����q�޽�{Ҽ6S��㍝X:w:     �+q�h/���F^}��  � p ��>����ꫯ��n�1<<|�8�j�"��z�,p    �o��?�k���}OLL  �� ���ӧO���V�=I�^�V#��o��V�S����     ��m��N���Ť�E�N�v�Z  @�� H���?~���ݓ���5pO|�t%�ύK    @w|�t5�I^���B|��  �"p  �ܹ�����V+莴��<Xވ�./��?�     t�n�v���O��OMM����<  ���(  ��<�y���x��Y����Q*���lF5Z����z�Y<     tַ�ע�n?�k��� @/	� H��?�8��_�%�dŽR�DZ}�d%n/�>�
    @gԛ�x���$���I���\�  �Kw  Rcaa!����V�ݑ���R;��;�t�t     �I�~�H�k��266y4??  �kw  R�ҥK���ݑ��U�z�,p    �o��?���y'ܽ{7  ���  ��'�|�}�]����F�^�GZ=�ڍ�J5����e    @'=�܉���U�Q����3g�  ��� �T����S�N���n���:́{��+�n\
     N�7��_���/��|�r  @���8  �w���������;��=��A������B�#    �II�۟m��>�ccc�Gw��  Hu  �������h�ZA�%�{�5���^^�;��    ����h���ύ��F�LMM���P  @� H�b�333���t^��;9ZD�}�d%n/�F�P     ���lƃՍ�ey�oݺ  �w  R飏>����#9֧=p�����v,��
     ����F���熇��a�$���v�Z  @Z� H��/���`�����FFFb{{;��ޓ�;    �1������Z𲱱�ț����.�  ��  �V�߿?輿.ҴZ�H���Xۭ���x     �n~\ߎ�j-xY��B�w��  H�;  ���'�ܻ$9`'+�{{{�v_>Z�����     ��|�t5xY2����dhh(fff  �D� @jMMMũS��\.�7::��������e����     �h��ˇ/e򲼭�'.]�  �6w  R�ƍ��?�1�$pςv��/���q1     8�{OV�W�c�~���  ��� �j�a������f:�T*>Ezppi��嵸{y>F��    �m�Tk�lk7x���122  �6j  R-	�gggcyy9�d�=�{�Վo����Ks    �����A��HB�d&On߾  �Fw  R��O?��>�,�$p��ގ,���J�Y<�b     �fՃz����Z��ۓ��ƍ  i$p  ������j�t���p��h�Z�v�z#�/�����     �;~�-����}qq1   ��  dµk��/�:/��	*�Jd����Ǎ��(
    ��՛����z�jɚy2 �'}�Q  @Z	� ȄO?�4�ݻ��e��R�^�?�Gk[qi�L     �j~�~��jy[o�������  ��� �	���133���Ag%�{�|�xY�    ��V;�y�����x���۷  �L� @f$+�}�Y�Y�b��)�Z�Y��[��[�qa��    �?�am3*�z�zY~9�R�׮]  H3�;  �1??###���tVr��J������    ��~j��M�{x2��������  ��  d�����/�:+9�ommEV<�؎����	     ^x����j�zccc�'}�Q  @�	� ȔO?�4�ݻ�V+蜡���gJ��fdŗ����s�r     �½'+���)p���8� ��� �)���133���Ag%+��r9�������|�    @�m��by;;7�^8|ɋ;w�  d�� ��IV�?�쳠���7[���x9>��     y��cC1�d||<�"y��ڵk  Y p  s���cdd$�����I�
�h�ۑ�>[�;Kblh0     �j{o?o�o666y����b1   �  dҍ7�O�S�9ɡ;�ܫ�jdE�Վ�/�'W     ���G�35^���K�i^|���  Y!p  �>�����/��j����d)pO|�l5~�t!��q    ȟ��~<Z��l||�0rσ����  �
�  �444333���tN�k�V�{�]�    ���ӣe��o!	������  Y"p  �>�����ς�)�J1<<�Z-���+q{a֊;    �+����qm+x�d�=y�4�;����  �D� @f������H��������������%+�    @~|�x%Z��Q�zi�X�<XXX���+  �C� @�ݸq#���?����5_?]�ۋ�c�T
    �~W�����������G^|���  Y#p  �����9���h[�阁������ȒZ��<]�_-]    �~�������R^�����  ��;  �688�����ɓ�s����//ǭ��(y~   ���ޝ>�Yh�>��-�؀1�;lll�l�Kg��d:==�n*5U���n:@��8x��]�*˖dk�۷�3�tX$Y����qT��*��`]��9/(�����>/��ͩ���?�y�  @%� P�������]X>E�>44�JS�����'}(     eu���L�Xo�����T��e�'�x"  P��  T����tvv����ayK�������J�)Vܷ?�&u�V�   ����ʩ�7���.�@� @%� P
�v��|�Oq�_�"(��-.w��    �l������������]ʮ��f��  *�� �Rعsg>���LLL��Q��{����e]�w    �TƧ���/@[[[���u����  �Tw  Jc˖-9r�HXŲM]]]���SiF�'r�ʍl[o�    (����f��l�j܋���{.  P��  ����?�cǎe�S�˦XqN%��lYכښ�     T�"l?y�z������X5oooOwww  ��	� (��p�xv���?,�J�G���Vܷ��    @�;r�j&����W5���~��  @�� P*�/~�<���R[[[�+�8?���Xq    *���T�Xo_�bټ슅�͛7  *�� �R���Igggn߾�^MMMZZZ2::�J426�׳��5    �T�/]ͤ��y����p)�'�x"  Pw  Jg׮]�����hmm����P��oYד���     T���9i�}A�a���)�G  ��  ��Ν;���gbb",�b����6333�D�����ky�ч    Pi��x%Sz>��TC�nݺ466  �@� @)mٲ%G�	K�X�)"�J^q���@���MC}]     *���DN]�毾�>���)��{.  Pw  J���ϱc�*ve|�kkk���}|j:G.]ɮ�    �R������Ά��������tww  �B� @)544�=�����^��^[[[� 8z�jv<�P���    ����z3,L5�O?�t  �L�  �ց�_�",���֌���RMLM����ٳ�     �t�����>MMM)�b�g��� �2� PZ===s�r�����Vс{�X���|dmZ    �R�˹�Caa�;��۲eK  �l�  �ڮ]�������ܜ���LOO�RMM�����o�     �T��d�z�������jjj�{��  @�� (�'�|2�|�I&&&��kmm����������1     +����\�q+,Lcc��W��_�>���  �ǿr (��y�#G������V����L�p�r�o},     +͗���}���w��  @	� (�����رc���	K���infjj*���������t�6    `��6<����yP��www�} @	� (�"�޸qcΜ9�^��~�Ve?�;;;�C�rpǦ     �_�W��444��jjj�o߾  @Y	� �
/��bΞ=;2��Z[[+>p/��v3?ذ.��Z    ���Wn���+�z{KKK֭[  (+�;  U���z�\�|9,���ƹ%����T���_���kOm    ������8eܟy�  @�	� �Ŋ�����Yq_mmmJ��pchn顮r_~     +[�����ݰp��ͩ�/oS��lݺ5  Pf��=  �'===����͛7��*K�^����yg��     <3�����H����;v8� ���  T��>��կ��*�p�՘���T��Gs���l\�*     �۱�k�S�����.O?�t  ���  T��{,����s�NXZŊ{�B�⾡�;�55    �_&��s�╰8����զM�R[[  (;�;  U��g��o~󛰴����7o�F�&r��Zv>�6     ��.\���Y�2�����d�޽ �j p ��<��S���2>�ץT__���挍����kW����M    ��+�7N\�S��K�e������1  P�  T��۷�СCai�e	��'��޳�     ,�/�dfv6,N��^[[��z���  �B� @U���Çgz�S�K��3[�K����d��k��d    X>7������a�:::RV===�^� ��L� @U*V\�x≜<y2,��	���֌����gf��������     ,�b��ū��OKKK�j߾} �j"p �j8p �N�*���JQ<[���p��`v>�6=�    Xjn���[�a�ʼ�^���Y�&  PM�  T����<��ùt�RX:��X˙��J�����y�m    XJ���W筷߫2�{��	  T�;  U�^�����3,����ܺu+eqyh8�7o��U�    X*���֝��x��JCCCʨ��6n�  �6w  �ڪU���ӓ7n��S<�Z����Y����=;SSS    �{55=�?\��M��۟z�  @5� P�^|����K���>MMMOY����+�ٲ�'     ���+�;1�$)Wʨ8g߱cG  �	� �z�֭�[xK��T(S�^���<�fU��j    �Xw&&s��Z�7mmm��-�y��͛K�� ��� ��ڿ���1,����fvv6eQ\:�x%�l\    ��:t�r��g½)�kʨ۟{�  @�� ��ڴi������hX�|���w����y]Oښ    �P��w�wu0ܛ����3�2�� @�� �������{/,�2~h`zf&�����;6    `�~�w�T/_>(e^o߳gO  ��	� ��mݺ5}�Q�޽�FKK�܊���t�����l[ߛ���y�    ,���n���r��<(e�7nܘ�F/� P��  �<��s�����)V�o߾�������ճ;RSS    ��353�/���{���T��8o޿  ��	� �?عsg>��3+�K��������ȝ��|=�֯	    ��9|�JF�'ý+�z{}��  ��  ��ݻw�w��]XsK:)�/����5����    �#c�9�5ܻb�V)���z���  � �/<�������3>>�Fq�088����ʡs����G    �m>?۟��p����RWW��y�G��b   �;  |�]�v�O>	K��o޼����]�뿚-�{���    �����p.ܸ�FgggʦXo?p�@  �#p �o�{��|��WVܗHq8_�ꌌ��lffg�ɩ�y�m    �����ߟ�K���>---)���ק�و
  ���  �œO>�/��",����R�[`ʆ��     �щ����FWWW�h���  �D�  �b�޽���399�]cc�����D���������    `bj:__��F�Rh1�R6�֭�{  ��;  |���ڹ����*,���������s���`ú     |q�?�S�aix]]]ʤ��8  ��	� �;�۷/����T�wE�~�����Φ�������!    @��9z7���s��A���L٬Y�f��  �sw  �Ŋ�����"w�]�FS�쌌�����g���Kyi��    ��gg.�v��A���OKKK�f���  ���  �G�<���ǭ�/�����+7�m]o�vY�   �jt���\�U�3����+e���[ʟ  ���  �G��e˖;v,ܻ��ƹ�����է}����s��    @���W���*�S��?�a  �o&p �yx�r���LOO�{W\Fܸq#eucx4'�g��k    T�C�rgb2,������եLV�Z����   �L�  �P__�'�xb.r��������MY}~�R6�v���!    @�����������J�8p   ��� �<�������jjj�"��������t~�w1wl
    P~�������z<��LKKK��z;  |?�;  �Sccc�mۖ�G��{���Q���p��`�X�:��.��    �'���ȵۣai�q���^  ���  � Ŋ�ɓ'355�M��kbb"eV�6�������    (���|yn ,�b(�L֬Y�իW  �nw  X�����ر#_�u�w��č7Rf�w��������p    ����̥�OEYjmmm���K�8p   ��� ��߿?'N�(����P\Pfvv6e��������jm    P�n����`Xz]]])�u�֕�g ��"p �*Vܟz�|��������E�###)����|r�|�|f[    �r(��>��^CCCZZZR&/��B  ��� �"�ݻ7����d�7�����C�9{mpn�    �|G/]��ѻa���e��#�̍�   �#p �E(Vܟ}��|��'��K<���K�}z�b^ՙ�z�   @%������W��Y����y�� �¨*  `�v�ڕC�UE���:::���xwb2_�Ⱦ�    T���.fjz&,�"n/Ff����y  �O�  �`߾}���½immM}}}���Rv���eӚ����-    T�����XeZo/B����  X�;  ܃;v����}�ܹ�M��~��͔���l>>}!���>�4-    P9�ff�Yߥ�<�1���ƔŦM�J��  ��"p �{T����?�s�7���������hN\����    �89��aytuu�,�������  X8�;  ܣ͛7�O>���HX��ֶ����=~q�?��v���!    ��74z7�������0��^[�lI}�,  ÿ� `	����?���T���r��쬚�}bj*����W�|"    ��V��~�w133΀�K������  `q�  �{�ttt����a񊅞��挍����~3��-�    +ױ��v{4,�����3��عs�ܫ�  ��� `����������{S\bTK�^����<�՞��   �J4:>�C���)^�,K^__�ݻw  X<  ,����g�������:w055�jpwb2�?s1/l{<    �������	˧���駟��v  �7w  XB�/����Ά�+V�o޼�jq��<�fu^U�K    (�SWnd`h8,�b����1eP�E�  ��;  ,��kצ��7׮]���ޞ��������N��}��4��    x����8��WWWW�b���  ��  �ث�������W��/^�|k[[[FFFR-F�'�����ۼ!    ����鋙��˧��an��ZZZ�cǎ   �N�  K���;6l������uvvVU�^8�-{WemW{    ������0x+,�2���߿?  ��� �2x���������LX�b����9ccc�����N��O�<��ښ     ����t>��WMMM:::RE�_�   KC�  ˠ��1۶m˱c������n�ˡ�y��    ���]���TX^�+����)�_|1  ��� �2)�O�>���ɰ8���sK���;<|�r��NO{k    �����휽v3,�b��z����  X:w  X&����ݻ�駟��+V|nܸ�j23;��?��zv��T    `�MM��Ӿ�a����ύ�T����<x0  ��� �2*����:w�����֖���LOO�����#����    X~_�����DX~eYoߴi��K�  ��� �2+�[���1���a������Ƚ�|y�?z����    `�\�=��W��%����%��ͩtuuuٿ  ��'p �e�q��tvv�֭[aq�����Uۇf�����sy{����    Xz�9�G�.�H����ݝ2xꩧR_/� ���_�  p����������8���ioo���p�M�u|�Zv<�6    �����@n�˯��1����t�ϱ{��   �C�NU�  ��IDAT�  �Aooo֭[�˗/��)V�1p/|�w)�;��Z���   �JRL����ٳ'  ��� �}��k��o��o<s�H�S�mmmM����ɇ����۵#��5    ����L>:uޙ�}RWW7�Rg�+~�m۶  X>w  �O�C�M�6���/,N��^��{����x%O?�.    �����K�}w<��z{MMex���  ,/�;  �G̹s�2==���1���K5��|^Ց���     �704�SWn���Ë�J�z��_�>  ��� �}T�O=�T:�����}ff6�9q.�����V��    <(�������p�tuu���6���_  ���  p��۷/Ǐ����o���e��FC�w�չ����H    ������ܙ��O�W�G}4  ���  �b����?��ð8Ŋ����S�_��GVw�.�)    �o�쵛��)������S�s�^x!  ��Q�A  @�ڹsg��⋌����kmmM]]]���S�fgg����_�>�����    �����puww��mݺ5���  ��;  < ̯~���p555s+�7oV�����x~�w1�o},    ����ԅ�OU�hƃR��466����ū�  ��#p �dÆY�vm�^����=�n����L���ky��+���
    ��N]��K7o�����{��Im��4 �~� ���o��?�yUGڋU\(�����})����_�>���   �7���g�����Ԕ���T�����ر#  ����  ��x�u�֭9~�xX����gvv6����d>9}!wl
    �犳�ߝ<����p�Z�*����&/��R  ��O�  Xq@~�̙LLL������[q/"�jv��`����5�}a    K����\�5���ƴ�����[�.k֬	  p�	� �����������������HU��>:u>k�����     �}w,_��_�����  �`� `ؾ}{����ܾ};,L��^,�{5���G'�絧6    ����l~s�\�gf�����0��f%{ꩧ���  ��� �
��(��n�/�/F��>::Z���7�r��Z�?��\    �ۗ�28z7����^���>�l  �G�  +Dooo}��\�p!,L}}���Y߅��jϪ��    @5α�k��+�j;::R����  ��� �
����g?�Y�����+��dzf6���O��L]mm    ���ON�w'��K�F����^�:�=�X  �K�  +Hccc�y�|��aa���>::�jw��X>뻘緸�   ��|t�B�NL������kjj��+�  x��  ��<��s9~�x�ܹ�Xq��������l��
    T�c��rq�Vx0����"�J���Wt�  e"p ���_ί~���0imm����g�=;���    (��U�/�����.����T����/  X�  �mذ!����~�zX�b�]��o�'����y����    �ezf6�9q�_�;�J_o߻wojkk  �w  X��x�����?2;;毱�1---�{�nH����+���u   �2�����u������H�jkkˎ;  �w  X�:::�e˖�<y2,L�$p��/��g]wGz;�    erq�VN]��J_o?x�`  ��E�  +��/���g�frr2̟�?73;����O��LC}]    ��NL棓�ÃS[[����T����g�ڵ  V�;  �`����������)�������x>>}!/m<    P�fgg���3>5�b��8ǮD��]��   +��  V�;v��/����p�����477gll,���+7�pwG�x�'    PɎ\��˷��>HE ^�T��۷ϝ#  +��  *�o��w�}wn���+.W��S���ٞ�7    T�#wr����`篕����ؘ�{�  X��  Pz{{����̙3a��w+�njz&;��wmOmmM    ���[�=q.33�@�"l���N%����K/�T�q>  T�;  T��_=?��O399毸d�|ٚ�t}x4_��ϳ�	    T��O_�����*�]+5_�vm}��   +��  *DqY��/�׿�ufg��WSSSZZZr����'�p9������    �'/_��k7ÃU�UwuU�b���k  V6�;  T��[��СC�W�		���oO��O��L[Sc    `%�9z7�?��U�VU�z�3�<��F�  ��	� �¼��[�ۿ����̄�).,Z[[s�Ν�'�S��Ѿ���m���)    �orz:�;�ig�\]]]Ů������  ��'p �
��ё;v�ȑ#a��w��_�~{4_���s�    �D�;y>#c���[�zujjjR�^}��   �A�  ���������X��������ett4��#��dmW{��    �$G���[������`�D7n��� �� p �
T[[;�6�_�*��W�gggß����j��_�   �����h�<�V�J]o������  T�;  T�6d����S,+�###��MNO���}y�����    <HS�������X�2+q�����΍�   �C�  �7��_��_gzz:�O��>::j�����O�.f���    Jqv����+C��^����[�  �,w  �`���ٻwo>��0?�s�����D����h��    �×�f`���J���8w�Zi����^{-  @�� @�۵kW�9����0?�jO������>:u>��[���    ����ɡ���Q���۶m��0  � @)���y��w��T[[����ܺu+������h_�yvG��    ����T~{�s����)mmm�4���o߾   �I�  %��ۛ�7��ٳa~��}xx8333�/ݺ3��N����    ˭�ڋ����dX9zzzRijjj��/��   �I�  %��(?��O39�h>���>44�ٙ��y��=�֯	    ,�C.g`h8����iiiI�Y�vm}��   �K�  %Q�����|��o߾m��;|z�Bz:����    X�7o��ūaeY�zu*MqN�ꫯ  �lw  (�;v����߯x����+7o��lzf6�r�t~�gg��		   ����oO����lX9Z[[+r��駟NSSS  �ʦN  ��y뭷���V�穣�#��Ù��
߬�d|�h_�xz�܇    `)L�����g2>�ln����I�iooϮ]�  T>�;  �Ll��?ȡC���+�����\�~=|����|q�?{6=    X
�;y!��w����ٙ���T�����_  Pw  (��>}}}	߯��mn�}||<|��/\����<�fu    �^�t5��+K��^]y�۶m�2  �A�  %���8���������ˏ+W���������Ҝ���    �b\�W���S����ե�477ύ�   �!p ��*Vv�՚cǎ��W\������]O"�陙�����ɞ�ij�'%    3:>�O����lXY���W�_{�   �F  �{��s���ܹs'|�U�V	�硸�|�h_�xz�ܓ�    0�x����d|r*�<�hJmmm*ɦM��f͚   �"p �+.#�|����̬E����А��������604�/��gϦG    ��ѩ10�g�����$���s#/  @�� ��֮];�b����_�������.gu{K_�:    �]�^����n�����'�楗^���y  `~�  P^{�\�t)������ե��+CCC����Ĺt�����%    �M.��saejnnN[[[*ɣ�>:�  ���  �@�b��������+�����t�nS�3���O�'{v�����    ����|x�\f���b����������_  P^�  �Ś͆r���jjj��ݝ7n��W\R��/o<�u�w    ��ټ�L�'�����ޞ���T�^xa.r  �˿� �����[��O�����݊��۷o�]��@�����<��    @��28r7�L�X��իSI֭[��<  @�	� ������W^�����7|�U�V��իa~�p�rV����5�   @u;r�j�������+�uuuy��W  ���  �̦M���C�ʕ+ỵ�����9ccca~~{�l�Z����%    T�?����U��tww�Rk����Kccc  ��� @z����,����+�a~��g��_��_�ٙ�r   T��w����3������Y��s�b�R��m�  T�  T�b��������w+~Wmmm�3:>���T~�k[�kk   @u���ο9=�_V����tuu�Rk��z  ��!p �*�s��=z47n�߭X�s�Nfgg����o���+;�    �733�����[pge��驨u�ݻw���5  @�� @{�����<333��O��FCCCa��]��C�yf��    Pn����˷�����Ғ���T������?  P]�  PŊ՛�{���O?߭�H���T��/�����)�֮    �t��՜�V����T�be�G?�Q  ��#p �*W<���ח7n�oW\��Z�*׮]����"�ގ�    P.�7o狳�a�+F<S)v�ڕ���   �G�  �w����s��ߣX�onn���X��陙�w�t�yvGښ*�   ��v��X><~6���ae�����Օ��bwww�y�   �I�  �E�/��B����݊K��~�Tuwbr.r{�����   ��6>9����ebj:�|Źf]]]*A���  ���  ��}���8q"�/_߮��a�Y����0�#w��3y��'RSS    *���l��h_F����W�ivuu�����{M  �^w  ��y���������d�v�󸣣����	s��P�8۟=�	    ��S�s��h�������Z��   �M�  �?Œ�+��������l�f��E�>88�����ܘm��   ��r��@�\u.V)���*f���.?�я   p  �̦M��裏���uttddd$a�>9}!�-�Y��    *���C9t�r�555���I�8p�@   p  ��[o�����g�nժU�r�JX�����������t�4   ��mp�n~{�\��+�ū����G�O<  ���  ����y��������577�=�{�Ν�p�S�y��鼽k[��y
   �Rݙ��{�Ogjf&T�����������W^	  �)  �o�裏f���9}�t�v�W��ݻw3;;nh�n�;җ7�ޚښ�    ��L#�O���d����sC&���_���  ��_  ��z��W���?p�͊%����ܺu+,Ε��|x�l�x<5"w   �cfv6�;����+I��d{{{*�ƍ��V   �#�;  𭊅���~;��������Օ���LMM��9{m0mM����,   ��⣓�304*K��^	�����  ���  �w*.Cv�ؑ�G��oV��www����a�_��֦��|dm    x�>?s)}WCe)^�ljj�JW�����ks#+   ���  �^/��R.^���akMߦ��-###��Y�Ŵ55���    �`���#����R��W�N%غuk֬Y  �o"p  �����/~���̄oV\dvv6,N���ؙ���֬�l    �ץ�����b�<===����J��ښ���  ��� �y�����ݻ��矇o���0��[���M��佯O���;���    ��w���3*PSS���d%x�7  �]�  ���ݻ7}}}
߬��+������
�7>5���d�yvg���
   �܆���ޑә���c%Z�fM*�~���1  ��   �w������df�E�7�����իs���poF�&�"�?�=�u�   `y�ON�ç36i���x���� {��	  ���  ��֖W^y%��^�f---imm͝;w½)����Ѿ�������   ��553��������Py���jժ�tuuuy��7  0w  `��lْ�'O��ŋ�+�ccc�����[����غ1    ,��������\����7��+������ύ�   ̇�  X��������ܽ{7��b��xr��͛�ޝ�����<���    �4>�7n��T�ŋ�+݆�y��   ̗�  X�b���λ�;���_������h&&&½��l�\����    po�ȉ��2���̭��t���y�W  �w  `ъ�ݻw�/��l��չ|�rX�;y.-�yxUg    X����9tޙU%[�jU����o�97�  �w  ��<��s9w�\�_jjjJ{{{FFF½���Ϳ>�7�ޚ�]� ��ٻ�/9�3��w眣��X�!
!$�P ���?p�Ú��0��$�s@����\������P���:��>�խ�9����} ��|:4��,_I������ʅ�   ߖ�  �iO?�t���G����%�8�����f��������������Z_    |3�����";7,_�������-���   �.�  �M�����<>��do��c6��_~r&����h��    ����d�{�|d���嬡�!jjj"������ݻ  ��  �b�ڵ�~���p�B�����cbb"�����1�J�[G?���*   ��665�;�L&X��A�d�|��#�De��:  ��  �&�������Bn�Qkkk���Ɯ��f|z6���I�U��   ����T�u�lnX �[�'����ƍ�[n	  ����  �7���{��K/��l6�����hll����`��LN�[��ƞ;7GyYi    �T:~�ə����������b>�����z(   n��  �W---q�������555�&ܧ�&fͧ�c�5ۻ���%%   P�R�Lnr���L�����Dggg�d�ɓO>   �A�  ̻��;.^���%�Q�*����`~����{��ǎ;6��  ����f���chb*X�������2�Ur����?  `>� ��o߾�����F*�
����:���c||<�_WG�w�/�C��   �b���ůN\��1gO����"�53�%����   �/w  `A$/�J�W_}5���/K.����"����\�`T���}�   @�����:<�$/��m��9�]�  `>	� ��bŊؼys�:u*�����hkk����`���:5��mMw    �?��������Ԕ���v�����  `~y�  ,�G}4z{{cl�Ԩ�WSSuuu111̿#��&�o^�    ��K�q��0�B�D㭭��϶l���L   �O�  ,�����?�t:���jjj*��l0�~�J.r_בߗ�    7�T����J_P8:;;s[ �UKKK�w�}  ��  ��K&�?�����o���\�W�%U�_�~=����oO]��X��    ��l�`��ܕ�p444��T�U2]��'�  ��"p  �ڵk��n��'O_VWW����/�_&������wl�   �|�`�^�^P��ʢ��=�ٮ]����2   ��  X4�<�H������p�e������f����"r|��X��    ��������LGGGn�c����;���+   ��  XT���G�J���J&3577���P�0��������m����!    ����G�7�.FV�^P���s��U�o߾=   ��  XT���ݻw�k��f���ihh�����$wF:������]�6EW��   X~z����(���������"v��   �A�  ,�U�V�V�~��������EOO���3I�~.vo�5��w"   ��K���N���$nO�<棒��x�'r�K   ��  X��\�z5��*//����N*��_=���m"w    ���܈�N\�LV�^hjjjr��Q��{ߋ���   X,w  `�8p ~�����l�W���199333�M�s��w�m��   ����s��3�lPX��<��񮮮�6N  ��$p  �LEEE�ݻ7~���Ŝ��_���}}}~.l&��_~r&����h��   �|sml"�9v>�q{!jkk˝�棪��x�'  `�	� �%�����sO��O
����2���bdd$XXI���G��ɻ7GSmM    䋡��x���He2Aᩮ�Ν�d���={���4   ��  Xr۷o�+W�D�W�����T���k:7��l�{s4TW   �R��_=�iq{!J򮮮�W��{o���  �R�  ya�������s�������鉹��`aM����NǓw��Օ   �T�'��-q{A������L6V�^[�l	  �����  �����ݷo_��'?s���+��444,�\���\�^W%r   ���L�}�\̈�Vmmm444D>�����{,   ���  �ɴ�x ���௒ˮ����o|z6���L��֨�   �hlj:���lLͦ�����|TRRO=�T�5  ,%�;  �W�n��.]��W����===��f���\&������E�   �������(++�|t�����dy  ��� ���L	�я~db��H.�ZZZbpp0X3�q��S�����P]    eh|2�:v.fR�p�����Ѻu�b���  ��  @�IV�:t(^x��d2��˯$�������l��t.ro��   �ohb*�:z6f���
Y2����=�Q2���G  �|!p  �Rr��k׮x��7cnn.�\kkk����Q2���OƓw�M��   0_���<z6f�����3�����ػwo   ��;  ��֮][�n��G��K.����ڵk��N�㍏NŞ�6Gs]M    ܬ���x���H��^ccc���F�)))�'�x"��u   ��  �k<�@.����>�\�������D�xr��ǧ�m����.    �����x���Hg�AaK&����E>���r��  ��  �{����^��7�)���ӑɘ�fR�x��ĝ��]�   |=�c�މ�ɊۋA����F�I�g�~��  ���  @�K.�8/������$?���v���l:���L��vkt4��  �o���|d�sA�knn�����7�cǎ   �Ww  `YH.]v��o��f�͹ LTWW�~.7n��l:o~r:ߺ)��   �_�:�yܞu�U***r[�Myyy�ݻ7   ��  X6���[�n��G��kii����H����Jg���ѳ��6�;   ��.]�ߞ�(n/"]]]QRR�$y=O<�Dnp  @>�  ��<�/>��joo����`񥳟G�m�+[   ��]�6$n/"�������7��{otvv  @��  �΁�?��?brr2��eYsss����/���9v.ݲ>ִ5   �.��g.ǜ��h$�ѓ���&َ�e˖   X�  ��SZZ�^x!2�L�����ӹ/_&������wl�   9�{���_���ܲ��+�MCCC�ر#   ��;  �,%�2;w�z�%�ioo�����f���K֌�{�|�ۭ�ĭ��   �c���_.�ť��#���+�H^�޽{  `9ɯwV   �����c�֭q��� ���,����ڵk��H>l�ӗ"�����oZ   ���\�ǯť��1���#����Į]����:   ��;  ��=��100��"���6w�6>>,�?��4�S����U   ���?w%��ť��"�]1�|�{ߋ�.C  ��G�  ,{���G155D������L�R�`�����LܿiMnZ   P��ss����HP\�s����;�Y�fM�y�  �	� �e���4:/��Bd2�(v�eZ21���/79��s��Z�>��|h��~O��   ��L6~u�B��ŧ��-*++#�444�Ν;  `��  !��y�����u&�Tknn����`i]�Mr�qǆ(/-   �p$���9~.��Mŧ��6���"�����޽{  `9�  cÆ144~����3���1==SSS�Һ:4�?:��m��
o�  �Lͦ��c�bx��K1*++�����'�f�={�Duuu   ,gn� ��r�����`\�|9�|Eroood2�`i]�1o|t*��ks�VV   �|�O��[G�ƍ陠8uuu�"�|���F{{{   ,ww  ��<����/榹��-����729�x2vߵ9��   X~F?{��퓳��8577GMMM�-[��ƍ  �� ��t����������t�䲭��!nܸ,�d������w��u�u
   |�������1��-�XUUUEkkk�U�V�}��   �B�  ����x�g�^�LƅcKKK������l���fS��ǧ�񭛢��.   ���7r#�=q>ҙlP�JJJ���+�g������;w  @!�  +�Z�{��x�7bnn.�Yr����===E���3�t����x쎍���1   ��u��p��Rd��U�Yr�VQQ�"�q���(--  �B"p  
ښ5kr�y���?D�+//ϭO�C2���g����Ǻ��    ��ɞk��W(rɤ�d�F�H����z*w�  Ph��  
��wߝ��ϝ;�.��������� ?d���W'���䊸{��    ��Ǘ{?���[2�=�ޞO}��hnn  �B$p  ���?���q���(vmmm1;;�T*�]��t&�ݰ:JJJ   X:���?}).^�[rN��Օ���/����rK   *�;  P48�?�|LMME1K.咉S���Vk�Wbbz6ٲ>����   �I��wO������������|�v��\�  P��  @�(//�C��/��L&�Y�V9��n�}��<8o|t:vm�U޶  �b����w����������룱�1�ESSS�ر#   
��r  ��444ľ}��W^)���uuu1==�㦑��7&���'��5�3!   
���T�}�\LΦ*++���3�E2E~�޽  P�  @���z(~���}��������/�ˍ��x��S���M��P   �����:y!f�Ž��ϕ��DWWW��|PVVO?�t.�  (w  �(mٲ%�������Q̒K�������l6䗩�T���xtˆX��   ��;�?���lqB௒�|�ɓ�;wF}}}   �;  P��)����Ŭ��<����ڵkA�Ig��αsq��5�yeG    ��dϵ���O�����/���X�re   �;  P�����?�|LLLD1����]�ݸq#�?sss����1>3�_�*   ��������O�t���/$S����#_lڴ)��  ��� ��VZZ?����?�q���D1kii���٢�9䳣W�bj6ܺ���ݒ    ��d[گO]��Cc_H�	�����$?�\�����  �b$p  �^uuu<x0^z��d2Q��˻������l6�s��193�ݱ1*��   ��fҙx����6V����G���QQQ����>v��   �J�  ����طo_���Ew�����0��w�F��t�ܺ)j+���   ����t�}�|�O�^Ǘ%g�uuu����r�8���   �J�  �_��;v�w�}7���X���Dccc��Yӝ�oL�/����[7F[C~\�  @�J>,��c6��[IP���� >���(/�r   �ͻ"  ���iӦ�q�F��O�b���333�/���l*^��T<�y]��̏�X   �7g�����l�4�%Sғ�%%%K�Rr�婧�ʛI�   KI�  �w�oߞ�^~���(f����l6�_��\���ܚ��׮   �sɆ�/�ƱO��JWWW^LKO�Gy$���   �;  �WڱcG.r���b��D������܅0��K�165n^e��   �,���oN]��Cc_���5jkk��e���{�7֮]   |N�  �O<�����/���H����hii���� �]���عuSTWx�  @qJ��s�|�NN|�$lOμ���͛c˖-  �_��  �'JKK�СC���8����X544���l�������D�z�D�ܺ1Z�~
   ,��}�{'��t*�U***���+���5k����   �L�  �5*++�?�A.rO�RQ����I�|��&ff���N�#���5m�   �����ݙK���|���������Xj��ͱs��   �	�  ��de�����_�l6�(����쌞����,7�L6�=~>��[��t   ��/�~���u����@��VSS���   ���  �H&��ٳ'�x㍘�+�)`eee�Ƚ���h�M��t��ո1=�o�%JKK   
I��ߞ�WG�NKKK���-�ˈ���8p�@^L�  �Ww  �oh͚5������_��wUUUn}���p�|��c�������Q    �ar6�?C�S_'�И�XjIԾw�ި��   �9��   ��w�7n܈�?�8�Uccc�R�������Ň'�񭛢��%*   ����d�{�|.r���LL���Z�%%%��O�G   ���   �����###q���(V�ī�����Ǎ��x��S�����!   `9�pm8>8s92�l��I���������~<�@�   �	�  ��'�|2^z��b�\�uttDoood]&/+3�t��3�}��ضƥ*   ����\|x�7�}��MtvvFee�R�����cӦM  �7#p  ���y�x�bll,�Qyyy��?w����}�p5�����뢼li��  ��2���oN^�ޑ�DKKK���/��ȅ�w�uW   ��	�  ��d���>���'''�UUU�.������������[7F}uU   @>J>����b|z6��������֥~�f͚x��  �oG�  p���=�\.r����b������1>>,?�S��_N�#����-�   �$�p�g.G:��&***���k�_Ftww�Ν;  �oO�  p�����?�A.rO�RQ����r����L��̤���O�Ķ5�����   �Zvn.>���>���JJJray�yq)%���   |7w  �yPWW���_~92�L��򰣣#z{{���/G�����t<|ۺ�(/   X
��}�b���6�����ť���O?�t   ��	�  �I2�i߾}�ꫯF��f���Gggg������\�<]�_|x2�cc4�V   ,����x�ą����6Z[[sC(�R��1�ۗz�<  �r'p  �G�
�ݻw��Ç�2򮪪�����~�z�|%Sܓ�����ǚ��   ��p��p����H�� nN}}}n��RJ&�'�z�<  @!�  ̳[n�%v����^QF�Ʌb*�����`�J�3�α��mMwl_�2JJJ   Bvn.>���>�������V��TVV����   ��	�  ����333��e�L�J��111,oG���&�?tۺ�,/   �O3�t�������m����6*.���駟�}   `~�  ȶm�r���#G�����"��g��vep$^��d�ܺ)jL"  `~�O�{����l*��J��+V��RZZ�w����   `��  �=�����q���(6�%c����7����LN�+GN���ƺ��   ��q~`(~�Jd�ـ�+*++��5<��c��/   ��  `�=��C111�.]�b�L�J.����"��z�Ke2��o�#�۸:�JK   ��t&���|W������%}?�p�^�:   �w  �E�gϞx�Wr�̋M2I+�t
���k�5�;�l��꥝�  ��165����UCCC455-�󓭅۷o�6   C�  �H���/��rE��������6��Pޘ�W���o_�Z��R  �����P��ܕ�w��������cI_�w�۶m   ��  `����Ƴ�>/��B���E�I&k�R�
�L:o=[Vu�=�W�;^   �2ٹ��ūq��Z�ͨ���+V�&�/�M�6�=��   ,,�;  �"J"������8&''�ش���"�����p��:C�S�Ȗ�Q[Y   ����_���S7#9SK���ϥ�v��x��  ��'p  Xdɴ��{.7�}zz:�I2a���+z{{s�;���F��������ʖ�   ��]��\��t:�fuww��ԖʪU�bǎ  ���  ,����������ܓI[�����=���c&��_~r&�����V.��p   �Fvn.�\�'{�̇������Y��'q��]�  ��#p  X"I���$����(&�ĭ�rr`` ����r�J_ޘ�G����
G   �bb&�>y!�ߘ�����ظt�����cϞ=  ��r�  ��jkk��������Yt�{2y���%������;2�9���;�  �����h��R̦3󡮮.��ږ��ɳ���   ,>�;  �K.�I�/��b�E���L&���Aᙘ�����;o鎻nY%%%  @a����6y}r�ߖ6�MUUUtvv.�󛚚b�޽  ���  ����8t�P���ˑN���$Sܓ�}||<(<I��ѥ���o_5�  @aH>���S�b`�{z�Oyyy�X�"JKK���I�~���%{>   w  ������<�L���?�T*�$Y��D�SSSAa��?���x�u���)   X�._��^��t&`�$Q�ʕ+���lI��l�  ,=�;  @I��<x0~���bQRR������Aa�N�㭣gc˪����UQ�  `�Ie2q�BO��0���dr{E��l���˝ˉ�  ���   ϴ���.�~���U�\vuuEooo���p��:�[_���룱�:   X��'�7�.���L�|K΅���� �۟}�Yq;  @��  ����ؿ���?�l6�"Y?�E�^L�w1�1?���$�d�;   ��dϵ8r�jd���[r�D�K!��:$n  �#w  �<���{���^{��b�du����ǜK�������D��x�ֵQU�   �L�����K�3<�ZZZ���iI�����<�L��;�   �'ޥ  䱕+W�SO=���zQE���b2��ڵkA�|}$������GWS}   ����g.�L:���룵�uI�]UU���+++  ��"p  �s�V��'�|2��D�d-u:�������O���O���]�+���$   X��\����8���,��������D��  �)�;  �2�z��صkW���[E�'�3�L��Y�^���W��o�F<�e}�WW   �ktr:~s�bOL,�$,������{���6  ���   �����2rO�T'��'''��p��D��ȉ��-��si֔  ��C�W"��,����X�bE���.��+**rq{mmm   ���   �H�?���_���"������닙���8�ҙ����?z#�۰&����  �X̤��3��ӡр��D�+W�����O��   ˇ�  `�ټys����.��=YW�������J���q��z���÷����   `~���g.����,��|���;*++���3��   ˇ�  `ڰaC�R0�ܳE�6<����ٙ���d��113o||:���{6����~�  �9��#{�L���Ő�����,�s��   ˏ�  `�Z�~}�ٳ'>\4�{�J:��D���=�W'��&>|��h�w)  �]����N_��3����-�����I���3�Duuu   �|�  ��5k��޽{��^+��;��L"���������x�/'��]�+���4w  �o*����/���177�Z[[���yџ�D�Iܞ�%  ���  ���+W�����W^)�໪�*����ڵk.�P����W��o�F<�y]4՚�  �ޘ�ߞ�cS���x������eџ[SS��  ,Sw  ��L4?p�@.r�d2Qjkk�;r�8]��W����׮�������4w  ���|H��Ձ��rod�>$��ihhȝ�,�$n��g��\  �\yG  P :;;s��_}��H��Q���rS�������ȅ����h<tۺh��
   >7:9���>4>���3��j���������   ˜wu   $�8|�g�'?�I�D��4�dj���HP�F�s���Y�*6��  �bw��z����Hg��)���l\lIܞ�����   ˛�  �������0����E�777�&�����+���g.Ǖ��x`�ڨ��  �b313�������*������dQ�����  �;  @J��db�O��H�RQZ[[s�����bwuh4~������k���   (����>�T&��***bŊ��'�`����  �;  @�J&�?��s��K/���l����\�>99��T:�=~.6t��}�DU�#  �p%S��J��l��(//��+WFYY٢>W�  P���  �������gff�tttDLOO$�����u+c�   (4g��Ǒ=���d��=�ۓ�}1%����   �;  @�����E�/��bQD�%%%��ٙ��g�$���%��?8s9��ƿ�zK�UU  �rwcj&>8{9�G��J29}ŊQQQ���M�ݻ7   (Lw  �"PWW?��s����d��r���+z{{#�J$�����|<��veܾ�#�a  ��&;7'��Ǘ{#��X*���$n���Z���  
��  �HTWW�&����gLMME��"r���t:�H�3��sW����x�ֵ�T[   ����T����/���ߒ����;w޴�V�^�?�x   P��   E$�tL&����Kq�ƍ(t�����g2��/���+GN��kW���]��  y-��~�Ӿ8z�?7��R����3jkk��6l��~8   (|w  �"SYY���_~���BWQQ������E�|I&��#���k�����V���   ����x|p�r�M��������_��%A�����w_   P�   E���4�}��x��Ws��]�1�=�������x�/'��]�u+��4w   �?{����8~u �Lm'OtttDcc�=/�۷o�۶m   ���  �H%�������q�ҥ(tI����-r�+e���蕾�28ݶ.��  `������^���T@�H&�/fܞ�������[  ��"p  (r{����{/Μ9S�ᾘ����/r�+�NN�k��[��������4   �l:��g��䓶��hjjZ��%��y�X�n]   P|�   Ď;���>��|�^UU%r�k%�N�^������n�խ�w�  ������=1�J����hnn^��%[�x��&>   ���  ��{�'����w����>3>=o=kښ�lZuU�  0�Ʀf��D�ȍ�|���---������x��'���=   (^w   ��֭[s����[�{GGG���͹28��c�uMWl[�e��  p�2�l��?�^鏬���dj�b�����hhh   ���  �/ٴiS.�>|�p�O7������N�;�R��]���G��n]�u  �]]�MmO6GA>jjj����E{^ru������   �  �֬Y�����_�"��t�$rO&�_�vM�ο4<1�}x26t��}VGU��  ����MŇ�z�|�`@�J�����E{^�<x0*++   na  �J]]]��3��O��H�RQȒ�T�;�F�\��nY��숒��   �g����<�{=�*������E���СCQZZ   ��;   �TKKK<��s���/���L�$rO.p�_�.r��I�������q��k���:   ����T|p��gN�$6O ,����ػw��  � p  �k%��?����_���¾�������I��T��x�r�xܶ�#��[�e.� ���t&>���z}���W__������+V��ݻ   ���  ����:����=7�}ll,
Yr����md�sq��Z\�{7����-  ��Cq��՘N��]r��յh�۸qc<��C   ���  �o����#����(d��n2]opp0�ۘ���_��kچ㾍k���"  ��1:9�?{%����Ŏ۷n���sO   ���  ������s�=o��v�;w.
YCCC��M&�[%Ϸuep$z��b˪θsMw���  P�f��8��@��:Y�!Y&3n/))���/n���   �E�  �����Guuu;v,
Y]]]�O�;�E&���W����Pl_�26t�  PX����ǑWc:�X.��wvv.ʳ��=�X�^�:   ���  �<������|�AA��"wn���l����8�?�mX-u5  ,��������T�r��������سgO���   |Sw   ���[���Y���[��f�P%�{�J�ڵk"w������_N���ָg����p,  �Q�!�/�������f1��d�߁���6   ��p�
  �MY�vm<��3���<R�T��26Y�=00 r�;K~w����hܱ�3�X��%%  �L6'{��'W�"�)�yS�������mQ����IܞLp  �o˻I   nZkkk<��s��$����P��Ԉܙ3�t��bO��Ms_��  @��:4<%Ƨg��Ōۓ��'�|2JKK   ��;   󢾾>����_��}tt4
U�wuu�"�l��>n���t�}�\�nm��6����   ����t�����X�3n߰aC<��#   7C�  ������Mr?|�p|��Q����s�{�ȝy���h.�ټ�=��neT��  �tfә��ro��n��Z�u���eQ��}���뮻   n��  �y���~ꩧ�wމ���lPUU%rg^e?��r��Z\�>�ׯ���  ,��������K�1�J,g��'gA?�p�_�>   `>�  X;w��8r�H�$r���>�;�fr6�=u1N^�{֯���   ^�ȍ��121�ܵ����eZ�?���bŊ   ��"p  `�|��ߏ������]�xeee.rO&�g2���28>�?9+��ލk���:  ��7�������t<�,V�^QQO?���<  ��"p  `A�z뭹����_�t�0׻�'��E�̷d��GN�Ʈ��{튨��  ��%ۓ>��g�cnn.`�+))�����9�B�������D   `�	�  XpI�}�С���~�T*
Q2�L��B���ř��q��Pܾ�3��銊��   ���t&�}�'{"��S3nokk�}��Eiii   �B�  �(ZZZ�?�a����199�(��W�X����ҙl����㮵+bSW[.b   ��䃣�>���zc&U��(N��®���T��~Κ5kb�Ν   I�  ����������w����M:/D���I�I�>;;�&gS����q�Ӂ������%  �����8r�'Ƨg
I2E=9�H�\ڝw�۷o   Xhw   Ur������݉w�՝&���}߽bv�I�b�	�@�!��Lz�O�+g:�L���B;�m�b�1��}�U�kL�ɮ*=�9�|�RUI:ǖ�[�{����q���(GUUU_���'�<S�q䃳�?8��]͍  ����8������������u�{9O<�D�ٳ'   �fp  ��x��'���#�y�X[[�rs�Amhh(���6���t�z�����mۣ��6  `+��_�?}v!7�C9J;�m۶-jjj6��������  ��E�  �[f߾}������Z���D����������Ym�l�φ����Dܻ�7����jo�  ���/-�{��K�Q(��Ԑ������@�o����x��7�!   ��UN   n��6���������oY6���{OOOnt����l���x������Hܳ�'��苚�  �r�����σO_��B!�\����p{U����҂��>��   7��;   �\KKK����9����QWWWnV��WW������H������*�  ���j!N_΋<�VV�YCCC���oz���{�G}4   �Vp  �(�������x�7�̙3Q����r����X�Ͳ��'>��b(��������  P�R���K�yQ���9/����������+l��{,��   �[I�  ����3�Dwww=z4��֢ܴ���0���hY�|��/��^�v�}]��  ����<�K��޹��_Z�
��w===�nO����?�C�:   p�	�  Pt���������B�妹�9�܇���ܹ�f���ˍ��v�Ǟ��Mo  �U(�ŧ#��޹�1���U��GR�f������?�G466   w   ���ݻ�����������Qn�E㴵���PY��)~�s��ӟ������bwOG  @�I��?��?}v!���onߥ��=���6�k����O~��  @�p  �h����/~�r����r������ҥK���p+�����F�C�]���5  �|16�����[MjmO�����o�'�|2   ���  P�jjj���������ܹs�������~r_YY	�UF�g��?������mۢ��9  �V�81'>�"�f��z***���7��7oN���������   (F�   ��M�s�=G����{��B�)�?00�C�KKK����L��އ���-��=�M  7Å�x��`^|	[Qz����/7�kTUUŏ~���>   +w   JFj���#G�D�P�r�.0���CCC1?���[�<zۚcߎ����  �����>���s[Uuuu�᭮�nӾFCCC�����d!3   �M�  ��r�wFwww��W�����('W�!�����b049oL~��ͱo��;  #��ua|:�=w!�f,�ek���͋�S�}�������   �N�  ��������J���188�$��S�?]Ԟ��(CS3���Ggsc����{:  �U
�>:��bL͗עe��U=5�of�����Gy$   �T�  P�҅ߗ^z)�~��x����ܤ
��6� �b163G>8���;�bOOG^�  ߥPX�OG����y���b ��͹Y}��T齓ÇǮ]�   J��;   %��������7ߌ���('�Bw�=<<,�Nљ���ߟ�4�����z:�R� �o(��e>��Z?o�l�������6Kj���O~��[   �R#�  @�۳gOtuuſ�˿���|������*� ?�arn!����B����%� @�ri4���`�--pYjkO�a���fI���?�|^4   �H�  �����/��r���188央�.�ҥK��,Bq�YX�?|t.����w�DU��; �V��Z��/�Ʃ���R�=��7�U}߾}���   �2w   �Fj&{饗��ߎ��?�Iuu�W!���ŀb5��<s>����;�����*  (o��+q����ɷ���Z������7��>;w�   (u�   ����ƿ��o�P(D�H��s���\@1Km�)��qGog�7��  �%�������xp4V�h����&/ZO�͐B�/���6�  ��$�  @YڳgOtuuſ�˿���|��+ۙ������T@�[^Y�.ǇG���ط�/�7�� ��glf.>X?��th,
kk�muuu9�^�I;[������(   ʅ�;   e���5^~��x��Wcpp0�IgggTWW�;��z:si4�����o{_l�l  J�ŉ�8}a8ΏM�����o���<�@<��C   �F�  ���."���K�?�!���X+�f��Op###e�sQ�R(*���Ƹw{o���Ȼ  P��b�O�����brn!�����-���7��{���;w   �#w   ���{,�������B�墩�)7����j@)���ߟ�4���bܻ�'���Mj6 ��-��1>�4��_���� ���x���+�7C}}}^ȟ�   �r%�  ���gϞ���_��W��P>��uuu�m۶�t�R,--���������_���==QW�m+ �[e~i9>�.����J W'�"��766n������s�=��   �3W
  �R����W^��^{-���X[[�r��'���ᘛ�(E��+������ξ��o{o4��  7���|���p|:<�By̕�f����������
�o߾x衇   �w   ���t��/ĉ'����erO�{{{cbb"(U+�����p��8�m�q������  l�4������_��&�v���9ܞ�o����x��gs3<   l�   lY>�`�ܹ3~��_���b���R�.�����Mx��)���81�GkC}�=�w�wGuUe  pc�WV㓡����P�,,p}Z[[���;/:�hy��f��  @1p  `KK���_ƫ�����Q.������CCC���P���g�ǻ�.����ս�^� �Z��/��ǗF��9��K����My�{�����   �"w   �����x饗����q�ĉ�i=��������t�R,//���4����8}q$�ۚs�}{gk  ���gpr&N��G���Ƥ�z{{���i�_���*�z�رcG   �V%�   _z衇r ���^+�@xuuu�����c~~>�\���ŉ�<Z����;��* �����O���C1����K�������|����Ə�㨯�   ���  �/�0��/�����s(��f���������r35�<s>�=w1���̭���� �U��/��ǗFce���H��nO-����<    w   �+����ӟ�4�z��������Aggg����{��L�RC����ő�ok�A�흭 ��s��ə8�~>t~l2��������QQQ�������]�v   p��;   |�Ԝ�.0���뱲�堥�%o����M����81�G[c}�=�{z:���[a @��_Z�O.��G��1����koo�����4G��O~���  ���   |�;v�����կ~���т���144����lrn!�~�y;s>vv��]��1��  ��J[�G�#���P�Cl����������m�����SO   ���  ��H�������~;���(5559�>22sss宰����Z�o���aw�� @)Im�g��r[���b �'͛������vC_7��ӎqw�qG    �+x   p�<�/n��曱���.]T���������[Eju?��x���Z�����n����<_���������)��   PN�  ��ٳ'oO��_�*fff�����f���^(�
�� @1���F{{{tuum���޽;:��   ���:   �F�i���E����q�ԩܨX�R����@���r�V�� (����I��}�����>��q��w   pu�  �:<x0v��o��FY��S�{
��&������蛭�w��f���  �,sK��ɥ��xp4f����|���?jkk7�uSX��^����    ���;   ܀�;w��/�����cxx8J]j���������R���O>�cg�Ƕ��t��վ���"  nTZXwq|:>���c��K;�������F����{�'7�   �N�   nPjx��OǏ�'N�ZS����ϕB��B!`+Ka��c�y�&���qWwt�4 �����3C�qvh,WV�u��ۣ��kC_3��?���y�4   ���  �y衇���o�W_}5����544��CCC���@���j|48�G[c}nu���;�k�� |��ť8;<�\���� n�+��555m�린�/����   p#̬  `���_����o�ٳgK��=5ϥ����HY��a#M�-ĉO/ğ>��m�q{_W��n����  X-��c�qfh,���r��	�A������]�6JEEE8p ���    n��;   l����3��'�|G�����(eW��&''c||<��Ka���y��:��o�����  ��t^0<=g������X.� ����������܍�Z����hii	   `c�  �&��;r��������h������p7<<�B!���������X��t�}]�T�q� @�]\�O�����ј^X���׺��6�5w��O=�T    K�   6Qj����~G����{/7:������O!���� ����B����x��`����ή����� ����872��ڇ�f(NWv%KM����*:�v�
   `㹚   7����s�[js_\,�Fǚ��r���� �[Z�ra|*�ʊ��������TU P:�n-�Ǧr����T
����]]]]����y�F���^x!�p   lw   �IRc�/��x������Q�***���),���B!�������&󨪬���)쾫�=��? ��������L|24�G'��s�����DOOO��n��:�����?�A    �K�   n��5zjz;u�T��(�`xsss����R W/�宄ݏ~R;����z��ܘ p}R����t|6:�F�ce����a+I��lO�ՍR__�>�l^�   l>w   ����;w�W_}5�����������ctt4fgg�vK+�q��h���v��Ѳa�� �w[[[����8;4�����@i�������|�(�v�Ç��<   ps�  �-��K���G����{/jJՕ�����t/�n���7��Ʈ��������@	 \v%�~nd">��� JS�cwwwoX���:~���m��   ��%�   �������;�����_�7��-�SS���P�����[\�.��R_�����jn�� ש��C�3qnt"ΏN���r �+�wuuE[[ۆ�fooo��G?��&x   ��	�  @����m����⣏>*�� ضm[nr/��>���x���<�j�c{g[���-Q)� �i����q~l2>���e���&���7,����}�Ѹ��   �u�  �H���{�'~�����B�������D]]]����t`����J��4�G
����Ďζ���5UU D�����L|6:��L���j 壩�)7����FHϟ��<�   n-w   (2}}}��+�ěo�gϞ-�pxkkk�ʊ�L�)����xU��1���])���5��`kI���s#qa�XX���MEEEtuuE[[ۆ�^
�?��ñw��    ��+\   P���g�y&>�����oKKKQ�R�}۶m9�>??��Y-���d�|�y��6Ů������u� �hvq)>��/�����v�v(_���yQx}}���^sssnmOG   �x�  @۹sgnsO!��>�,JU
����DLNN�t+=����lhr&�cg�����꾳�-Z6& ����\^Е���Q�V������y~y�R�<>�`    �G�   �\j�{��⣏>������������=r�{)�PjR�}xj6��g�����ho]-���-��n<$ �i�P��RK�����[Z`kHa����hkkې�KA������   @qp  �q�]w��ݻ��^�K�.�lz]]]l۶-FGGcvv6��ofa)>ɣ��2z[�r�}Ww{4�� ���Ÿ81_�MŅ�(������ڼX:ި������'�   ��	�  @	I�_z�8y�d���g
�(EiK������>66V�?�����)<��Ϝ�������;�ڣ��9*+* n���ZM����ߤ�G'cj~!��+5��yc������Ǐ~�����   ��	�  @	ڷo_n�����܄^����s�`xx8��R[��󨮪��������;Z�Q�; lay%�������ӱ����VUU�����ظ!��cǎx���Bk   �4�  @�J���������ĉ�������:bbb"�x��r�0�Ԝ��ܘ��;:��o7lH�& [K���ӳ���ߖ/ƧbrNK;���._)ܞ�7*���SO��&   PZ�  ��=��Cq��w�o~�nsooo�m�###���@qI�hF�g�x����������-1��]-Ӱ	@�I��\���cp},�hi�.-�Ls����y��۷km  �&�   e���9�����{q�رX]-��P
��v�ԟ���x�v�+a�q!jk���9�[b[Gk4�� [���rO����}n�c�oSSS�[��|�F��l���	   �t	�  @�������_���RTUU�����166�[������4���{-Q[�H�r���#�s�����T�����hii����iZ��;�����   e�U%   (3��^�ӧO��o�+++Q�R�!�,��ñ��@i�YX��������ln�����oo����\��ҴZ(���l�M������_,J��;�;R=�Ӽ�F566Ə~�����   �<�  @���{bϞ=��o�_|Q�M�i��������� JS��3:=�������2��Zrؽ��):���X
��L����l\����X-�޹%P��ꢯ�/��nD
��ݻ7~��    ʋ�;   �����x���O?�#G��dzn~���m�###Q((m+��8?6�G��͍����U轪�2 �5���ٹ�����}6��܈4�kooߐ���������i�   ���;   l��v[�ڵ+�|��8{�lI���m�o����177@�HA��L#5��6����ii�z�h��� `s,,��]6��f���ͭ� %�������7"��?��Cq���   P��  `�HA�g�y&���_����(5UUU9133ccc�ܡL�Pe
Z�����|_s}]�v����[Mu����_Z���hj&��g��[�����]]]yNz��������   �O�   �����x�W�w��]|��Q��v�)�022R�A}���,,�G�i��[��r�=�����(�𷤝{&��
�M����R l�������ɻq݈������;�3   ��A�   ��Ԝw�СػwonsO��&�%RXzz:�����uL/,��ɥ��qMUUt47DgSC��6G_{K��x��zR;���|��\nfO��+p3�E����9�~#�^�=�\��   [�w   `K��_��q���x��J2$����U����b [�����v������|_cmMt67FWKc��6�������r��Z��ٹd��_�83�ف['�Sk{SS��N
�?���gϞ    �w    ���w�uW��7�����(5555100��������$sK�176��.�^����ֆ��ji�M�)������P�
��7��1:���=5�;��Ecccn\����ݻw��*-L  �-K�   �����������s���;�������-r��Ғ�R��Rtrn!�3_�WSU����Ҕ�񽥾. n���jza1�G�fcd�r�}�P�b���]]]���zC���O=�Tn�   �6w   �k����~�ȑ8{�lɵ�����6���>55ZM�ﲼ��&g�"��[뢭�᫦�|��"
l�o6��������Uav���Pz
�WW_�e����������    p   �J
'<��3188o��F���E)��������Hm����p�R�}tz.�+M��W�j���>޻��r�{CmM \��啘�_ȿ_R�=ڧ�-�JN�suvv��nDj~��g���>    �p   �U���+q�ĉ�ӟ����QJ���b۶m1>>����WjX�YX�����W�7��D[c}]-M����u9�l])�>���s��}�򢙙��_��(})����55׿�/�՞x�رcG    |��;   �w=���q�}��믿�[�Kɕf�������� �(sK�y\��^�h8�W]Um���P�U�=}�\_������L�/���|nb���|�\?����e#Z��k�~�����Geee    �-�   �UI-}/��R|��gq�ȑX\\�R��۷o��������Ͳ�Z����<�ReeE4��F{c}�75\�7����������A������[�;:��ف�`#Z�[[[��g�����    �.�   �5ٽ{w�򗿌w�y'N�:kk��Jm����###��� 7K����i���B��ښ��ޯ��;֏5UU�<K++1=��C�s1�����t��QR�z�C�Hk{uuu8p ��    ��   �5K!��ƾ}����_����(%uuu�m۶�䞆�p��--�qqb�k���TGs}�������߷/�k���3Ky��t^tr���# ����===9�~�v��O?�t�C   \-w   ລ�����ş����農��"�����H��E�6��� n��s�����c�u�_��S����1��������斖�
�� ����'L�-���j ��R���+Z[[��5�<멧��y   �k%�   ܰ��/o7�ȑ8{�lI5�������@nr���m�@�(�����2������ʊh������M��9��T[�o7��)U�)����w=�M����ا�����\�������������~<�@    \/w   `C� �3�<�������6fgg�����}�澰� �,5X��oߦ��:��Gcm�W�)������6��fJ7ҮWB�)����q
�ϯ�N��P� ;�ƪ���m�)�~�����駟΋�   n��;   ��R���_���?�=+++Q*jjj��?==���Q(�\�q�siQ��_}���"R �.�kr���.ꫫr8>�S@�^<W!��/,_����������]LA���ʞ���jii����r�i���Ç���7    6��;   �)�����{�ȑ#q��ْjZM������>?? [Q���ڳ�����������h���������>௄��ǵ�I�Uė�Z�_Z��F�W
�ǥ���K���_������ (*i�ojmOs��������   ��$�   l����x�gr#�o����Q*��������9���ۭR��pU!����Z�k�*s�&�禀|uUU>��k�/�_[U���iԬm����K+��c%ԗV�o�p�j�?���r`==���Ws��PB�� �������^YYy��M�v������   �=�   ��K��?��O�̙3��[o���B������������v�ƤP�\j����W�O����c��J𽺲2��t_���]ݗ��5_�_��c��</=��2��ؤ0���JnL_Y-��k��j��K���5O�IǕ��Ǥ�.�ϥ�/����W�})��b���SWW�[���Z���in�1���   �fp   n��o�=�'Nğ���X]]�RPUU�C )̑�ܗ��~C1 �#��WV�n��K�o�������7�V��W]��-���_o:_K��o�˯�`3���J����A�kU[[��n�-    6��;   p�=���q�}�śo��ϟ�R��ܷm����y��" �mq��C� �#�J������~i8���8p�@�   p3�   �D
����122���Q
R�a{{{�������|   ����loll���yO���駟�s7   ��I�   ��R�����ԩSq���X^^�R��"}}}177���  p��pzkkktvv^W�z
�>|8z{{   �Vp   ��޽{��{����w��G���Z���H�����155   �JCCC^D\[[{�ϭ���Gy$��    ���  ����:>�`���1<<� }ߩ���9FFFbii)   n����<'I���*5��ڵ+�Ů��   `�	�   E���%~�ӟ�g�}����cnn.JAjIܶm[LOO���Xɴ�  �+͟���r��Z�����Ç���)    ���;   P�v�ޝ�ɓ'�رc���� Ls�}vv6   6Z]]]twwG}}�5?7�>��OD___    w   ���۷/��ݛC���_��B!�]jOLm�)�>::Z2�|  ��UVVF[[[tttDEE�5=7�:�����w�    �J�   (	)ı�����������Ν����(v�Mq۶m199�G)|�  @qJ��]]]Q]}m�y��{�7y�    (v�   @II���=�\LOO���K��>4�Z���se||<fgg  �j���Ewww^@{�v���ʋ�   J��;   P�ZZZ⥗^��/Ƒ#Gr�إ�Ş����������R   |�Լ���mmm������8|�p466   @)p   J���@���?��?�8���?���B�Ժ�m۶����A�B�   W�]�������r���=��S9   P��  ��p�w�q������+++Q욛�s����d   ����������������k׮    (e�   @Yٷo_�{���[o�G}kkkQ�*++s�b
��6����   ������؞دEMMM<��Cy   P�  ����!�����Ĺs�>�B)}}}177����@  ܸ�赭�-/|�������ٳ'��|   �\�   e���>�{��#G���x�kll������������  �/����Օ�^��ߵkW����   @�p   �^www��?�c�����b�+�����ԔC����  �����<OI�r�Eoooޭ*�    ʕ�;   �e�0��~������㭷��-�Ŭ��*zzzr�=�򗖖  (]�?5����\���\��'�̍�    �N�   �rv��?�����O?�w�y����q۶m��}||<VVV  (���y�jGGG�}5��N���9؞�   �U�   [�m�ݖ��ӧ��ѣ���Ŭ��)s bb"
�B   �-��wvvFu��_�M��'�x"?   `�p   ��{�'��'O����cii)�UjqL͏���199SSS���  @qI�S�����������Ӣ��<   `�p   �Ҿ}��HA�cǎ���r������� ���cvv6  �[���.7�����J�ݿ�a
   `�p   ��r߻wo������j�������ɭ�)辰�  �͗�������ժ���Ğ={   ���   ��Ԑ�~�����������������n� �r��)����W�����x����{�    �N�   �;\	����[o��q
�(V�}����������� @�kii���Ψ���������~���c    ��;   �U����C�Ł�w��]�;w����)h���SSS9辶�  ��hjj���X��q<�@    |7w   �kP__�>�l,//��o�]ԍ���֖�����133  ��K󁮮���������������   ��p   ���15�?��cq�ر8}�t���F1�������vOm�  \�T������W����_�   �:�   ܀\9x�`�߿?�=~�a���D1J��������sss  |�t���y�������#�ĝw�    \w   �P]]���>�hnt?u�T��S(���7s�}~~>  �������ۣ�������?�p�q�   ��p   �@�����=�[�}��8y�d,--E1�������t����  ��,�ӎG)�^QQ�M�ohhȍ��~{    �1�   6A
�?���y����'�:���ߟ��SнX�O  �,��=5��p��ۛ�����;v    K�   `��۷/�ӧOǱc�r�����4���bbbB� �����)ԞF����f�G}4�o�    lw   ���{��#�S����l����<����WVV  �IjaO���������---q���    6��;   �M��A��Ǐ���b����U�=5�� P�RX=���`{UU��}lWWW<������    ��    �ȕ����~��crr2�M
�477����t�WWW  Jɵ�SS{jlO��    �\�    ��m�ݖ���x���;q�X[[�br%�>� (W�c��ڢ���/�VVVƮ]�������    ��p   (��/���\��f�B���/�� (V���^SSw�qG8p ��   ���   �Lccc<��ӱ��ǎ�?���B�W��i\	�///  �J)�~%�����������   ��!�   P�jkk�����裏ƩS���ɓ9L^lR�{�y>�S0  n�fokk�㻂�i�fKKK�߿?v��    w   �"�:������ٳ��}rr2�Mj�LC� �����*7�_M����3~���#    �K�   ���ٳ'�������������(&W�����9辸�  ��R��Jc{
�������lO�   P��   JP����?cjj*�y�8�|
�(&y,,,�{: �����Ρ����]����;�3y�|   ����   ���=�=�\����ٳgcuu5�I}}}�� p�jjj���=����3؞X����o߾    �4	�   ��"?|�p<��q�ԩ<�����\	�/--���d���  |����������;���?�p�ر#    (m�    e���2�U�q���8~�x\�t)��֢X���FOOO!�~�B!  �����hkkˍ��&��n߾=8�w�    �w   �2500/��b���űc��̙3���Ţ��:��Spiff&�����  [SEEE455E{{{^�m�����x衇r�   ��"�   P�R��O>?���ԩSq��ɘ���b�BI����u3}_)込�  l�|0����i�I�#S�}�Ν   @�p   �"Rph߾}y\�x1�?�.]����(�����9��:��� @y����S��ۚ���۷o��<    �O�   `�_|1ɏ;gΜ����(�u>�p���*��y  nLmmm����i��=���΍��~   �<	�   la)D��O���8u�T�<y����uuu���9�>==]4��  \����hoo���&���P�Ν;   ��I�   �܊�o߾<.^�Ǐ�K�.M����::;;s�畠{�P  �[jhojj��������s��۷ǁ���%    ���   �����x��cnn.�;gϞ����(UUU��3�R�|
�/--  �%����zkkk^����F�;�37���;    $� �����X]]��}��t��jjj�   nLccc<��y�9s&�}���b��@����H�tO�w  n����lO#��}S
�www�������'    ����TW�&i����Z Ә����15B.,,��z�/��7"rR>]TI�ߦ�{���O����k��I�Bi�0��,  [��ߞG1���s��������<�(
 �͑�������jz��o��   �Ւ�ຬ�����dno�����������P����-�>S�&I!��q�L
���LGGGy;�� `�(�V������=���r�{1�I  �Y:�J�P�VY��v    ���; �*5������p}uL#��WVV��]i���Ǥ�tq&����<��N�  (W���D�B�4��*��  l���N
���ν�I[;    7B��dO��.�ŋ�1���b�Q�����Mi;ށ��ضm[>^�  �E1����UZ������N)��@  \���ޝ@g]������$d���"��	�E�E�}��V��ڱ�e��z�̙qڞZ���.ETv
HQED�N�	KH H��^�FDH����ޯs�yB�&3��w���ύ��wm��y.��     �-� �TVV���ڵk����ݰ`�W_}%x߉'\��FU�d��֭[�ѪU+5mڔ6#   �@mu���t7,%%%�6w�3  �8{���v�ׯ�ݭE��  ��a�V�gE���io[�r	gΜ9��<�_�=�۳{UVb���_��3tt�  �7� �lc-�(��u^^�kg����l��}�v7<l�زeK�i����  �`U��ݞ{7l���JHHp��ɓ.�na��@   ���Â���n�PUY8�
<z�꥔�   �O	Gii��=�n��[���x^-�^Wl}��U_=�JDl�`���� �[�@�ӹ۶ms�O��އ�`�sC�6�ݭ)33�I!   �N�v�ܰ֠��׻g^���7;dڸqcw�>�<��  �3�[���%���h�;u��m�   ��ٍ�TQQ�>|vX����׆'`_\\\�����d`mX����4�k!x  ���; 1�[;{nn������$5c'�?��37�m*edd���m"�kTT�   �``ϳ�{�v�6w֭[��{��kt���Y��!;xj�I6hu  ���y������۶�تU+��?Pll�    ȕf�����ڰP��9r$,���ކeW������.��ym֬��6m�� ���; ;�kA�/��҅����#���$=-�,P���]��ݳ���Fӹ�   ��Q�F>|�{�n�ڸq���{�c�.�,D�;  ejk�߳�^�z�I�&   �WZp�����s�v������q׮]n�+99مݛ7o�^[�hᆭ� �w p�w�>h�p����0o޼ٍY�f�)�gee�K�..�   ��mۺa����tZ�ܟhu  ��Bm����;�5F{   ��[��ؖ��f÷��ކec<lNbn�{V�g���  �>� `<-�6lp��C�	�.�Y��c'��u��6�lc�M)   ���(���ۍ��b7/�$���  ��kk�P�=�dff���/Wll�   �pa�j���矽I�u��a<������ۼ�}����֭[��L���  �� ��#,���矻ӨL��-��ނ\�R׮]]����-<   ���4:Խm!w��M��  ��kk��Gzz�z��ƍ   u���w�^mٲE[�n�Ν;]����ѣ���O�0�}�vw�_v�e�5..N ��F� ��B�_|�{����J�d��V�X�M�սW�^43   �y�����6�({������ǏwAw�*  ����			.�~nɅ=�dee��  �Pf�vkf��D۶ms�x=v���������e˖.�ޡC�j7Z �w �Cv�w͚5.�n��i�����0m�&Wvv�ٰ��t   �@�ZFm��jݺuڳg�_o����٨��PYY����   u���4h��~��Ђ�ڵs�:��   �������{vhOv�a׮]n,^��͗����Z���`0  �� |�&L"�P�ƍ݃4H,�~�z7<�����S��ݙ�   `%''k�С�m۸������'O����d��IIInX���ݭٝ��  �W�fF�a;;xW������֭��   ������Kw룽8���Z��kx��?�[`׮]���. @�!� >`M}j_�z���܇`Q��ݚ�z�쩾}��}���T3   �5jt6�~���<�o�>���,Tf#55�|�Vw�  \*+��@{bb�ق
[���7o���vc�   �Pd!v������@M����ؘ>}�[_���6hw���wc �"P�Z�J+V�p� �Y������HIIQ�>}4x�`���	   TM�4�����ۻw�v�M���Wee�_>���Q��f��6_d�  Ԅ��[������ξ�B�-Z�p�1�   �v�ڥu����>s�����%K��a�Ν;�2�.]�(::Z  � � �Ȯ���v��ٳG@(:|����kѢE�ԩ�����/����   hn�[��5�ە��`��֦j�Z�,�ns�ӧO  �|,�nm�6<7,�3Ezz����>    Y���O?�'�|���`�qڿ9v����z�r󯪇� �G* j)??�5[[c��S���X�;�l�aÆ�Y�f   �'�nϴ[�n��͛]3����111nXӪ�m�8qB   �hM�j���t��ڻv��Z   BV^^�>��cl?r� �,���ذ9Yvv�~���2@[� �w ����rwJ�>��a�N.�!�?�PYYY4h���y6�   �@T�^=u���O���/�t��#�nM��VV�|�9��;  �ǚ=�����;סC��   ����b�Y�F}�M�Xg��f�~���fw� ��� P���ג%K�z�jr���溑���������L   ��j�����r��URR◰�}>�`[ee�������ɓ  ��B���n��ƺ�YyD�F�\��]�v   Bѱc�\S�e0�������6��V�+��Bmڴ �{��l۶M,���k�`b�Ľ�3g���>\-[�   袣��3�O���͛UTT������Шk�4�v  ���x;�V5�nA���t�o�^m۶   �l�mӦM����׻5/ �ٚ�e��hڴ�������6 ��p�sXkߪU�\c{AA� Ԝ-F�ב���,6L]�vUDD�   �@W�������e�wE�?6�,�f"6��ۦ�5�[S  |�lѠAl�W[#���7V�ΝբE   ����>��C��~��Q�j����9s�f͚�.]�h���֭�� j��; �����裏\c;�*�{��k�2d����JEEE	   ��`M��6�ݻw��[ۘ�G���ᒒ�ܰ���naw�  ,UC�qqq.�n7�4o�\ݻwWJJ�   �Pe�7ntł�����6lp��q�����+--M ��#� 암����/^�'N�oj���?��_}��ns   &n{���/��_��OZH�Frr��[�����J ��g�v[���n��Z�r����   eV&h�|��:t萀pg_V��p�BeeeiРA�ѣ�� P��-k۳���L�P��P��ٳ�t�R:TW]u�{   JvK�cϹv���w��u�J�Fjj��fw��:uJ  �w<M�e����H%&&�P�]I+    �mݺյ���g�����zqnn�M�4q9�+��­� Ώ�;��STT��}�+��,lcA�E�i�����԰aC   �ȞemC�Fii�>��s�޽[ǎ��ϥj�����ݭ�  \����0{�P{JJ�ڵk��h�  @8�u��������v��! �c��S�L�;Ｃ����ꫯVZZ�  �F�@� �&��i~��$�  �P���p6�n�Ok�ڶm�����Q�x�|m�6O�8���
  ��~�Z�݆��GEE�q��j߾�233	�   lX��|�e˖�[�Nyy��J����_��vp �5� B^aa���}}��'u~E<��t�븮��w�3   �,�ֱcG7����]�}�޽�U�.Y0/11��[��vg� �wY���Y�ݮ��ז-[�K�.��   @89t萻���s�)�[�]�v�p���kյkWEDD �w !ˮ�����ŋ]K��`�!����?��O:TÇw�X   @(hڴ�櫯�Җ-[�ζAXYYYg���-�g���r����r�  ��:Tզ���T0���hi  @X�R��K���[��om߾]/���Z�h�J{����H@8"� �؆��\t]_��{�ky����j;�6�5N   �"::�5��0�����w=m]��[�ݞd�>�}lO�;�� �Pg����8�s�B�v��y�����v�v    \���kΜ9ڰa��u�n ����{������O^@����aavkk�?�ۄ�6��3gj���=z�z���U\   IU��-dna���<>|�N���a,�naw�9 
,`av�/��m�ֵ��4    ��ٳGs���ڵk	�~V\\�I�&��I+���+% �=�P����EEE�<�q��)33S��r�ڷo/    T��ƺÝ6N�>�;vh۶m����������6t���v�܆�+++ @0�\����Ҟ����eee�q��   @�dV�2}�t-Z���;��A�@P۹s��~�mm߾] 5X���U�n�t�m��Q�F   BY�z��O�!OkR���]m>v�Y]�p���6--��=�w�� ��iٍ$�s�j�Ϯ֭[��   �Â����6l�  ��j�}Ĉ�߿�[?�PD�@P��3f��� -����jذa����#    Xm�.]�0��a�wی<r�k|��a-��1������  @UU[����բEu����   ��Y�b޼y�裏X����	���[�օ뮻Nt% J�*Z�l�;=|��Io�T9�|�Z�J7�t����ˤ   a'%%E�{�v��߿_[�nUAA�JKK��Jik	��`BB���5�{��� ��ii��Av�_��͕��ō   �;v̵?/^��e0 /;�2q�D-Y��5����K *���<m�4	 ���ʜ�}�ᇺ���ղeK   �iӦnk��������u��A<����5�ڰ�}r���}|� �ڲUh�a7��P�6mԶm[   �0[����\㳭� ����+���}�|����� ;� ^aa��N��/��B p!�R���k���5j���   -��	����m۔����}���ׁ��aDSYY���w��  ��n�S�3$99�m�[����.s?_    \����^�Z3g��ѣG tmڴ�e&z��1c�(--M ��X��m���}�]�� T��C.]�T�~�������O    �f!�.]��a�6$;(ZPP��>u��?���H��ǻa,��	�۰gz @����9hoѢ�Z�j�v��)::Z    j&77W3f�О={ <ء�K|���:t����z�. ���;��dmr�&MrW� @m���(''G�|���NN&   �a��޽{������6=:��V�~}%&&�a쐻���^}�0 �/�9РA%%%�u��n�iӆ@;   p	
5m�4mܸQ ��W_}��F��>}����  XpP�������]+V�`�Wآ���iĈ��꫹�   ��sޭM=//O���:x�JKK}>_��^t��o!wϰM�  �EEE��������왙���    ^�	�ڨ��� >����^Ӓ%Kt�w�98 � �]�3q�D�` �d�vx�N&�;�m�   �8�m��c��{�����\ི�ҧ�Z}m����݆}N ��e�v�>n�v�D�ܹ��4i"    ޵a�M�:U����sٚ���g���W7�|��5 Pp�wǏ�̙3�|�r�/�ٳ�Mج��G?���   @�Y�<##��4ݱc�{�>v�***|���
]k��a�ƚ�,�~��	x�e� pa�}:::�m�7j�ȵ�ggg�aÆ   ������ɓ�y�f��X�ȪU�\	�1cԿ7��@D��_}�駚2e�� ��`a���&l����[   ��IKKs�w���ׇ�Ν;����f�s_� �'Li,`�iw��u� �;v�)..�؛5k�:�P�D   �[�����C���O ����2���Z�b���_�E͛7 � ���&N���k�
 �a߾}��_��믿^7�p�ې   p�RSSݨ���z?x�JJJ\뺯�MM			n���w���c@�������n��ܹ��6m*    uk�֭�4i�


 ��m�6������o�Q111�@A�@��k�rrrt��a�?�>}Z�g��ƍ����L���   �}~������]������� �������<�B�6,�n��w �.+�&���$�fҩS'7(	    ���P�O��իW�̙3�Ke�A,Y���&��=++K ��3�@4w�\͙3���������\7�|�$    �e��mۺ�QZZ��{��ё#Gt��q��x�6<l��v�໵�[ �EDD�����a���4]v�e�޽����    0lذ���ۺ	 x[aa��~�i���W��v�4h  �'� �]E>a��� ��,'Nԗ_~����]�   ��X��s��n��z���<�cǎ� �/DFF����6�(o�O��^9� TDEE����n�Zݺuso   <�&2c��Z�J �K��i�krss]��~ !�����g���>ۄ oZ�v�v�ܩ�����С�    ��5�7o�܍�����{�n8p�5�Y�ؽ�Z�-to��控��z?u�  �U�gdd(;;[͚5   ���駟jʔ).� u��ѣz��իW/t� �?p�36�z뭷�~�z@09|���|�I:Tcƌq�    �������j�޽ڷo�:��Ǐ{=|���X7<�e�>�O�݆� �}����vs5j���Lw+FJJ�    [ۘ4i�֬Y# �;d�}�v�s�=��� �%�Z |®�y���]� #kg\�d�����g?S�&M    0Y��cǎnxTTT���@{�����]�B����-�2ㆧ���-��	�۫/Z��/��cn���\{۶mթS'p   �v�ء	&���H �o��z��)P��n��l������zs� �%??_�?��n��v���_    ��m�ddd��a��v߽{�{���N�8���}l4����4�[�݆�[�����(w��^a���0O�-\c;   ��aks���ܹs�@@�nڴI��{�[�  _#��klSx���ڼy�  �X��7�p����.��    �X���t�Mָn�h���w�G�uW����u��Ӷl��6�-�n�w{�: �k_�� ���q��.�ޡC�o�   �l=�Zۭ� վ}���?�I7�t����*��)� �b۶mz�W�0 ��U�V�	�����Z�    �k[oڴ��*..v����B��QZZ���`����7��P�'�n!{O �^�1n��k�ݰ7�[�V�v��   a�� 'O��J�  ��:������_h�ر�> �w �l���:u��p�P�k�.������v�S�N   ��p��Ν;��t߻w��>|�l��W�[ ֚�m��j��3��qx�� ���SRRԼys�m�V�Z��f8    ��%���Z�~�  �X������]Ƚk׮ o#���l�N�X�B Nl���g�Ս7ިk���k�   �0�����;�Q��,�n�����Ǐ�u�_j����8�߫��W}���O�=>>޵��a���teff�fv�}    8�M�6)''GG� �cǎ�^���u뭷��� j��;�Z���q��iϞ=�pd���3gj����{'    ��kj>�5�:tȅ���ą����]�R������&6����s#pa���ns֚���m�7m��5�[3��>    T���g͚��r @H��e˗/�Ν;����� o ���6nܨ	&�X wve����'����q    �>��`��s����UTT����~d��'O����e���>��B��f;B�}}DEE��!��n�u��l����ccc    �`��W_}U����Pc%��?��~򓟨G��KE�@�ن��"~�w�܄۔oԨ���PPP  �8p@��_4v�X���S    PS��P�����n��eeeg��{���ǵ9��]�	�WVV������ EDD��u;�a�boذ�[�JMMu-��j    |i׮]z��ݼ B��T9n�8]s�5�����# �w �b����nM�-��g-U6�m��ܳ�mo{ެ�*>>�]�nv%�m�m޼YS�L�l���+��nЈ#�   �Uj��E���O��B!x��m6���]Y˺�m��q��JKKs�����   ���Z�J'Nt��@��u�(//O��w��@mppQ�!����+??_��gmT�a|���m���_l��:��k6Q�={���ۧ{��+_c    P]�	�;v̅�m?~܍'N� �'o�tS�P�5d۸�oYӻ��=�j;����~|�Oh݊<ֺ�Y�JIIQzz������	�   d6ǝ:u��/_. 7V��������Wff� ���� iZ��k����/��2eeei���:x�ڴi�m���&�m,�ƣM�|m�ڵ:|��~�_�w    ֘d�u�����F��G�����-o���	�_,ok�	�{T�����@`��ok��a�vd��ຕ/Xh݆�-Y�zrr�{��j    ���
Ǎ��;w
 }/|�'t�wh���� ��{mڴ�M�l���6 -�n�m۶n��t���/��m:������P �a�Uv��P�V�    ��:�����._ZZ�֒��6,_�ޮc�\7���$_��{� �������'$�ayO(�^=o��<A���m�ʚ��՚���ڍ���+    [�l����URR" w���o�����Z�j���Z�b�&N�ȕ��6-�ޭ[7l���/5jԈ�;pG�����7����:w�,    U���n4iҤ��[�����`��Z(�jS���m#�jx�s���V�Wf_���ws����x�/��<�s�����ϳn����������{�����������R���Ն5�[P    pq6�[�d�f̘!n?�y���z�ܹs�T �-_�\�v������. �b���p͞=���m@�o�^]�vUǎ]V���;�����^w�y�$    ��Y�ښ�mx���[���������m��y���sٟ;7�na�s� �6�{�/�n!����?�	�WekD>��������~�8�W�D�߳p:    ��ٜ��W�^-��ۺ��=��ږӰ���ڼ�s���y{�� ���IOO'�����|����/~�eff
 .��;���p���4j�ѣ��7v}�>g ���&Mr��#G�    ��<��6     �b�_z�%mٲE<�g�ԩ�Z�h�iӦ��zFF�Z�n��V藒����Di ���G��'�Џ�c���G �}�p�p��M����ճgO�j�J��q��pa�2:�������         EEEz���~!p4i�ą�m����k��^5k�̧a��!�|۩S���k����1b�yoD � \��g�a�����.�ޫW��^Y�l2f��^��V�X���2�w�}罢         @�۹s�^x�;vL𿤤$h�޽����2-[��?X�<�o�Z�}�ر�' |w ���'�t��Q7l�ԦMj��U(�8[}bb�JJJ��֯_�g�}V<��bcc          x�[�ε��W��X�`�Νխ[7eddl��)��O>q��_�򗊏� xp5�?��S:r��{vҰG��ׯ�kn5��N���-[����>� �4          H,^�Xo��6ae?����٭�݂����l��6�ѣG�v�ء����.?��* �C�S�w��3�<�UYu����{�V�>}ԠA�*��'�������O?�_��WJHH         ��t��iM�6M|��P��Vy����3(��� �|������ֿ�ۿ�C, @�C�|��gUVV&�NJJ��&X�pb�R�d@��ڵKO<�z�!%''         @`9y�^}�UmذA�[�Z�R߾}թS'իWO��2۷o��g�@,?���\�����af�֭z���U^^.����=z�䪦��g'���~��%          �Xy�3�<���|�nԯ__�;wV���դI����4�8˴������{]�
@�"����7��_֩S���`��\���o������         �����p��={�kذ�kk�ի�bccJ�T �WQQ�W^yEw�}�;� <p������~{ �w%''k�С�ڵkX�=�fP;�rM�=��Z�h!          �a{wO=��
߲v�>}��`����"�@͜>}Zo����!Y.@�	�' ����+''�����4h����ׯ_�N�j"""�M����+ �g-O<�|�A�i�F          �ݾl�v{��n�ZT���]� �Q�ܙ3g4m�4W�:|�p/$2��z�jn����pX���+�Ptt���w?~�]u����E          uc���.�~���7Z�j��:tP�� �5��۷O ��2o3f�бc�4z�h܁��g����_'��%6��֭�;��� |�M� xǉ'��s��7����5k&          ��{�nWDeAJx�ۇ��m�*Yi w�v,X�2pr� |��;�rss5~�x�>}Z�t������kմiS���d������O?����w|}         >����g�}Veee�wY�}ذaa{5{���Y�p����u�wr� w m߾]/���***�K����k��F�:u.�q���]v�����7�����         ��nݪ��'�=�!�����l¨���^�����t߫��իWO Bw ��ܹӝ(>y�P{����ݻ����*EGGՓ����9 �C��mroذ�          x�ƍ���/�ԩS�w$%%��+�T�=�VA�;����&���?u/ ���;B��٣�{�ŗ(33S7�pm�`��z_\\, �UXX�B���o/          �fӦM�۽�
��﯁�~}bi�wJ�X�f��Z���8H�(�$�q��=��3*++j'11Q�^{�:w�,Ԟ�8&���޽{��SO�׿��4h           ��c���⋄۽ ""Bݺu���Õ�� ����������p�֮]�7�|Scǎu߇ ��@8x�|�I����c�vkm'0z�,�y�f��ݻw���ׯ~�+���         @�؞�s�=��'O
��u�֮L�Y�f��Y���;�=+W�Tll�n��v-܁ g�O?���9"�\rr�F��v��	�a�1 ��}�v���Kz��%          ճo�>wk���ǅڳ�aÆ�gϞ4'�@ZZ��n�* ޳t�REFF�[n��A�b����DqQQ�P36��ӧ��lEGG�C���������}��ǂ         P����D���L�ۛ�֭�~����;j�L����?����뮻N Bw HUVV��_�޽{��IJJҍ7ި6m��׸qc��~�������4          �����.�~��Q�vZ�h�n�A͛7j��;�;�f�rM��\s� ?�@:s��z�-�ދ��ܹ�F����8�7bcc݉���R�y��)99YC�         ��*))�SO=���b�梢�4x�`���_���j��;�[3g�t٥+��R �w ͞=[+W���\���zwM|�&d܁�3m�4����=         8��]?��:p��Ps�Z�ҏ~�#��^b���a)// ���ɓ'���>}�@�"��O>�Ds���/33S�G�VÆ��aۼ�<��O�ք	����N-[�          ����z��UPP �LLL���^�z)""B��T�ٳG |�B�999��X��� 8p��֭[��믻¸8�ˮ���Yu+--M ꖝ�����#�(%%E         @8����+���ݻw5�����n���"�Lw���(p���z��ծ];>܁ a��_|�EUTTgW:�d���j2�?�9�g�}V�������8         �Ȋ�z�-���
��A�Q$�cd*��q��)��������t.܁ PZZ�~���Y�����k���jР���7 �طo�^}�U=��,:         ,͞=[+W���V$جY3���u�rwVh!���D܁ g'�^x�
�誫�"��gIII���r�~Խ�7jҤI���         ��O>�Ds���ǲ}����W_�������@�:x�ƍ��z��s@�`veք	�c���bbbt�7�S�N���8--M��� ����]��-D         �`�֭z���]���#G�s��B�IMMuō�O���a?rrrt���\��G�`���Ӻu�kڴ�n��V7@�����1c��٥K         ����@/���***��kѢ�n��f���u+22R���:t� ԝ5k�(==]�F���G�P�6m���/\X�4f�����Z��yny��G�$         E���.�~��q�¬�x���:t�k�X���;P��Ν��\y������X�Ǐ�*��	׀4l�0��	P܁�`�x����#��+        �Pr��)���*,,.����8;;[�/�TlٲE ��ԩSոqcu��I w ���kܸq�t1ί~��9r��w�..�@��srrt���s(         !�s��;��=��n�ͅ:�d* ������/�����wjٲ� &�@��<y�����KHH�wܡ-Z�---�imA��}��g�?����:         ���w�Ѻu��ڵ�+����e* �Oyy�^|�E=��JLL��C� ˖-ӊ+��KMM�]w��^��������Ç@`x��w����5[         zV�p�B��Y)����5d�!����_qq�^z�%��׿V��Di�@�W% 캬�ӧ痑���4h ��p���?��� 
         �8���n� kk=z�������20Ǐ �پ}�f̘��o�] w  ����W^QEE��]��ٺ馛\#8��ܷn�* ��رc7n�~���*22R         @09y�k�-//�/))Ʌ5�5k&���4�@ X�t�Z�l��
@� ����ӧ5~�xZ��G߾}u�׺k�|�RLvkȻ��         �`a����


��kժ��[;8�e*v��- �7y�d5m�T�۷��@��Y�fi˖-�w٩����Z^v�@`Z�p���u��M         @0X�`�֮]+�_vv�n��&EEE	��L8*++]I���G%&&
��p�h�֭Z�h��m��~�5��+���@�v���=��cJMM         �6m��n)�����O?��]���LX�9�B�=���ի' �E���Ǐ��^��ӧ�o���ȑ#գG!�%$$�k���;��c_�r�ᇙ�         `:tH���*��}�k��V}���w �l޼Ys��q�5 �E��I�&�	���o�Y�:uB�]�E�\[�l����u���         4�N�Ҹq�t��1���ׯ�1cƐ�R))).+SYY) ���mڴQ�.]��~��Gi͚5�7���[nQVV�Z����ݻ p�����ر�ڵk'          �L�2Eyyy·EGG��nc�/�YV�B�EEE8Μ9��^{M��\�' � �Ա��BM�6M��=��z�.\��ÕZ@೫'L���{Lqqq         ��U�\� ������Nedd��2܁�SVV�r���oU�^=�{܁:d��<yR��]�e��:���;��������'         ��B��ގoKHH��w߭&M���L��o߮��_�F���G��C�oǎ��<���C�1 x�\�R]�t�~�         �b�������˅o$''k�رJIIB�
 �͛7O;vTVV� �-�@�]����fW��=�p{���5�WTT@���.�LIII         �aΜ9.g�onMiii�Μ9�	&��SÆ��p���'�:;a����7�t�:w�,�>��NMMUaa� ���R����z��!         �.����\|�p{��|%%%z�7��_��P��u`�ԩ*..�~ȏ1B]�vM�����/�ԇ~�A�	         �+���?~�*++��Y÷��iMqqq���WYY� ��7jٲe2d� �mذA�V��v�uשgϞBx��1|f̘�nڰ         ��0e�	_������'JLLB�e*���r:tP������>t��	M�<Y�����էO!�؉r ���1슭�z�+�         �sk׮�@����$���?&�,����/ ��ԩS����#�<���H�-�M�6M��^�zi�СBx��N�6m�ʕ+տ         �bي�'
_KHH��w߭��d!�Q�]�vi�ܹ9r� �w�Grss9Y��u��Q7�p��,�n�gΜ��2}�tu��I)))         ��������L����5v�X����@p��{�.]ԦM������7� ��Z�j�[n�E����WLL��6���D �ˉ'4e����         �m�-��͛)66�5�7n�X܁�r��iw0��STT� �w�f͚��
w��{�m��~}����	w 8�_�^�֭S�=         xˁ��{�	Rdd�+lڴ�^���]����B ����z���5z�h�R������kٲe
wqqq�뮻��Y�����; 8Y�{VV���         \�3g���7�ԩS���ի�1cƨ]�vB������T
@�X�p��w���n�G�^d׏L�8ѽ�3;U|뭷*--M�Wj���ѣ�=�n�          .��ŋ�m�6A�����l!|YƆ�;\��[o��?����� �"�x�M�v�ڥp�Q�F�M�6�"���K��w��j۶�         ��***r�J����}�
�L�


4o�<��G? �"�xɡC�����+�0@ݺup.&c@��Ǔ&M�����:         ���=�7�xC'O�T��ҥ�,�L��ϟ��={�e˖�=�/�>}z�O�ڷo����J��$&&*&&F,R �mϞ=��?���C�
         ��+Vh˖-
w�[�֍7ި��܁�UYY���zK����U�^=�����jݺu
g��}��7�C��&���d�޽�f͚�^�z�aÆ         ����L���]jj�n��VկOt_#����<W8d�����Kd'��N��p�;�C���.��;���]���?��         ��>}��;�p֠A�u�]�������İ�� �����˕��, ���;p�/^����+\Y+��Q����&�b�w��:rРAjӦ�         ��ٲe�V�^�pV�^=�r�-��8�e*�����~�m�w�}p������Ds��U8�pcVV����J- t�9sFS�Lѣ�>�;         ߧ��B'Nt{L���k��@
��2yyy�֬Y�+��B]�t�KC�����u��	�+�t2D@upBK~~�V�\����         �>.ԁ�.��r���G��!S���S��?��?% �G���ݻw���Y			3f��>�.�N��͜>}Z B�;Ｃ�={*66V         ��>����+�eddhĈ.��;<�E������#��Ҍ3���,(�z�.��Ddd�RRRT\\, �����M�F�)         �\o���N�<�peي�n�M���pB�ܹsշo_W
�vxrj��>ӦM����V�Z	���pB˂4p�@w�         �غu�֮]�pe��G��@Ւ�����(�:uJ ��}Ϝ9S��w� �w��N�>�Y�f)\effj��j��7o��a���{Ocǎ         `,_1e��9sF�jذaj۶��ꈈ�Pjj�8  �o͚5.g���- 5G���e˖���@�A�3f�;a�Wj�i�ʕ�ꪫ���!         ��{��U��С����/�&,SA�o���{�1�v@-pj��ɓ�;w��5j�\
�@h��w�yG>��         ގ?�ٳg+\���h���.k��
 ��۷O}��$ 5C���E����D�w���ر��K�d]_|�6o���        �0g健��
G��k����X5���& ���w�u�;~. 5C��&�xY�=����ꫯ�qqq���WYY� ���3g�G��         Li�ҥ
WC�UFF��ڠ4=ǎӂ4j�(�>�@5͛7O���
7��������&d܁Д����?�\ݺu         "UTT(eff���w��Y�w��_W� 	�@���D�S9��֎�t���m����{g���1{k���tvg����*�(g-�H�� B!�����QAr�|>���gƙ�`5\��}]������~7��J=E&���@q����?�|6hx8wxW�^�w�y'�(��>��Ciƌq��� ��W^�e˖��     P2ǎ�ݻwGM�0!~��_e���J(�ڵkǝ;w�w��]��?�c G���C�&S6�gώ���C͕ZPlgϞ���?֬Y      ��o���N����~����RS!p��ٹsg���K1gΜ ������˗c���Q6�Dq�|UWW���� ���W_�U�V�P     P���q���(����X�hQ�PH�{�(�t ����}�˿�K �L�����_����(��>����w(�.Į]�b���     @��h/Mo/�����я~0T��ڻwo=z4�~�� ����ƕ+WJ9�=��)p��2eʔ����;w�P\���Z6ŽR�      ŕ�:u*�&}����,�������Pl���J���k _O�_����6_55^>��,�8��O(�s��ef��     �b���W_}5�h͚51����$p�b;|�ptvv�ҥK�j
V�
iz��mۢl֮]O>�d�pK2�;����x��gMq     (��۷���ts��/�0�cܸqq��� ��w��],Y�DK_C�_�7�(������x�F��Pi��|+W�      �%Mo�ӟ�e��ğ���Y�C-�|555eߵ�t���طo_,[�,���|��g������8Ə0�P�И�     �xv��.\��Y�bE<����%5w(�W_}5���Lq�� p�ظqc���D�̟??/^0R�P'N��ĢE�     �b(�������������&�Ŗ��wvvf�;�ew�O
�7m�eR[[?��OFRڌ�����_�pS�     P;w����G����?������dh �����X�t�)�� w���͛��>�2����S�NI�`Ŕ)S�ʕ+����>�;wn      �oiz�믿e�`��X�xq�p�C9��b���Y�|���{�nlذ!ʤ��1�{ѐ��ܡ<�|������       ����?ǅ�L��4�FB�)�D���� �����@���X�bۗ^z)ۄ�h�1cF9r$�rؽ{wtuu�6      �si�Q�|��ߏ�S�����L�<9�^�@�>|8�=O?�t ��� o��V���ٳcٲe�%�8�#]U��;�į~��       �����O��2I�m�;�	Iip����7ވ���sw��)�'ND�����mv��S��|�}����O~�Ǐ      �'Exe��ߪ��Y1�RSq�ȑ �o�޽q���hii	�+/�6n�e�dɒ�;wn�h�C�tww�����?�a      �/ip�C��L/^���#-� �C�������#p��_��gϞ=Q�����/��I�&E}}}ܺu+��x뭷�^p�     @���O�2I}�K/�0�ry����?�yL�:5 �;dRhw���(��k�:�ɘ�6d�O��<.\�}�Q���      �p�ҥ����L�{�9}�F���ŷ�~;~��_ p����m۶EY�i��?�|�X!p�rz�w�      9�q����닲H7��{�-QWW===���͛�'?�I�g�N�N��ڵ+�_�e��/d�;�NC9uvvFWW��      ����.�����_2������_(��7o���۳��N�N�	�e1mڴX�jU�X"n�r���-[��/~�      `lۺukܺu+ʢ��9�/_0ښ���P2�Ɣ��Q�T�L�N��9s&�=e���?�����;�W
�_~�娩�$     ���2L^z饨��
m�
(�.Dggg�������R{��w�,��������f�ԩY����@�\�~=����v     �1l߾}q���(��s��3�<0ܡ��z�-�;�'p��zzzb�ΝQiz��ŌE��2E�/^�|Ҵ�;     �صiӦ(�4��
�;������I����e%p��v�����Q)6���,m��PN����Ϙ1#      [._��Eve�hѢ�3gN�X1mڴlp`___ ����[�l�_��e%p���m�eaz;c]
[?��� �'mʶo�?���     ��%��[���R��/�0������ɓ�ʕ+��֭[�?�i�������R���#G�DL�2��vƼ��� �+:{���     Cz{{K5<pɒ%1k֬��f���w(�7n�|k֬	(#�;��N7���e���WWW�ei3�W�0�����x��      `lHQݵkע����W�X���ÇP>�������S:)l߱cG�A��h���c]ڌ��r���t�L�     0v���,���b�̙c���P^�p˹s�b���e#p�t8�/_�20����������Ҝ��lϞ=q��͘0aB      0����J31���*~���Uw(�m۶ů~�����S:;w�2H��;::�"m��P^w���"��{.      ]��ݲ���n3�555P^;v�_���R:wJe �+�u��yS#W�ǎ���{�=�;     �(Ka{������n�X6iҤ����[�nP>i`�}�b���e"p�T���[��޸q�bŊy�D<p����z�jL�2%      �;�˗/G̟??ZZZƺ4��̙3�Ӷm���RI�aˠ��#Ə�'w MٵkW���     ��غuk����?����Cy���i�{ccc@Y�)��7ofWu]�R�5k���H��}�;     �(���={�D<��1w�܀<�T@�����)(�;���Dooo]�>ˢ�<jhh�������	���?/^�3f      #k���q�Ν(��}�{y���@����{wJE�Ni�ڵ+�`ݺuy�nH��g�Pn����G     ��J�\L�<9�y晀�0�8q�D�?>fΜPwJ�֭[q���(�����Uڐ	��;     �Ȼ~�z)ڊd͚5QUU�ӦM����{�n �������/�PwJa�޽���E���|'��y��1��<y2.]��=     �������E����Ɗ+�$��S�LɾG�K�N��)�4	����룽�= ��@���{��_|1      )p/�e˖ń	�&5w(�O>�$N�:O>�d@�	�)�۷o������V�\�ƍ�3�;0 N�     �������2X�fM@�������۟��g�;� p����ۗE�E�����S�N�555EUUU)����ѣG�ڵk���      �4|(ݲ[tO=�T̚5+ �RS�k׮��/Ptw
��?�2x��c۶m����W��!#����c�ԩ���P?����w�      �>� ���v�,MpH���>}:�̙Pdw
-�q���Q===�	�����ĳ�>���Q[[�iC&p�;     ��z�j?~<�.��p�����+w�N�N�;v,�_�et����Y�~},]�4֮]���c]ڐ<x0 ���w��qP     `���i�`ѭ^�:�U�j	�s��� �-����Pdw
-M~-����/LuO�{[[�Mc����t3ɡC���Z      �4��*�J,^�8 �RSq�ԩ �����q�ܹ�={v@Q	�)��{��K�_y�l�{GGG<��1u�Ԁ�D���	�     �Ǎ7�ȑ#QtiB���ۿ��V���5 ����t���"�SX�/_����/����-[b�֭1o޼l�N*WUU�6�;0X
�����>      z��틾��(�������̞3f���˳^���> /��� I=ŏ�〢�SX����^:�|�ر�ihh�6o�W��ɓ'�����ĉ��>�����p�B477      Ck�޽QF/^�6��͛���-k%f͚0�8~�x\�v-�H�Na}����û~�z6�}۶m��SOźu�b��Q�TFZڐ	܁�=]�     0��޽[�����'v�ڕ=---�D�����������4�6����s����BJ/�]�zl`���i�b�ʕ�bŊl�6���!;y�d $����     ��9|�pܼy3���ٳٳ~��X�ti6pƌc�ԩS���:;���G	�),�;�t�ԩl"9�����ٕ\�6m��f'��͛g�;�Ήc`���h�5      ��{�_��ݝMt߽{w�H�VbѢE��bL����V^�x1 ������QS#�x�TSH酛���;;;�'������>`8܁�҇��V����      `h�۷/�j���q�ر�ihh��˗��իc����)5w I=ő#G��XP4w
����������T��k�ƓO>0������5�;     �иt�R�?>x8ׯ_�-[��֭[����֭�D�R	iMMM0��?�SHw
'M?z�h0�Ouoii�&�/[�,ƍ�L����q�Ν H</��r      ���p!���ӦM��+Wfτ	F����`�=������F�N�?~\;�Ξ=�=o��f���Ś5kb�̙�V:�N��'�����/      <�4��s���ذaClڴ).\�t#1#A�v���즑����"�S8�FGOOO�ڵ+{�������V҆L�Hq�ɓ'c���     �������s�����ٙ=3f̈�˗g�D}}}�p�������ի�D�N��ǆ����ׯ��K�ƺu벍<,2�~��     <�S�Nō7��w���l���͛���-�g͚0�Ə�&M����t3�����S(}}}q�ر`�����&��޽;�͛��R^�hQTWW|�;p?��      _��^===Y+�������hoo���ڀ����$p�j���E#p�PN�<�Ռ=�*�t� =�iGGG�Z�*�L�� w�~G���w�:$     �ҭ����g�f����c�ҥ�nݺ�1cF��HME� �+W�DWW�ފB�S()|c�K'H�l�[�n��T�ŋGUUU��tڸR�d�# �4��̙31w��      �����i+FIؘ&��޽���ĢE�w�[��Kؼ6P$w
%M'?Ouoll̮�Z�fM�א�f�<yr\�z5 ���;     ��s�ԩ,�f�n%b���z����qxX"V�~���{.�(���=��]��Mu߾}{vB9�TN'��o�+m���`Ǐ����     ��K�];�_���[�n��u��ł�|���� �{<E#p�0>��Ӹr�J�ow�ލ����I��+V�ʕ+c	A����ȑ#0 �      |;i�+c���ӦM�:��KL�81�A�N�555��� IWWW�O��(�;�az{�\�t)6l��6m��fS�[[[��p�p��/f�,�u�      <�Q06�]�|Y+�7JS��a�.��t�m͚5E p�0Lt-�t�t`�{
�;::�\}}}Plw�~�������      <�s���͛7�|�J�M�υ���ѣw
C�Na�8q"(�t���I�K�ƺu�b���A1	܁I��w     �Gcp`~��7o����X�zu̚5+(7Mp?�����BH�\O�>�G:���fOKKKvJyٲe1nܸ�8&M���>�u�V �     ��Do�����v�ʞ�V"����ʧ��) ;s�Lܾ}[CG!�)�K�.�F��Ξ=�=�ׯϦ��kVfΜC:q,f;u�T      �h�;���ĺu�bƌAy�����ݻYS1�����SB7���n'�H����իq�ڵhll      �Y�>�ܹsA���w�y��e�ĢE����:(��ST*������@���"�S�W�7pRyÆ�|��X�vmL�:5�Wj���Z�dI      ��N�<}}}Aq��9E��ihh�Z�U�VŔ)S�b����I�&����`�����@�N!���W�u�V�ر#v���rN�Bx�t�M�     �pR�Ny��y˖-�u�ֿ��/�����X�w�;0؉'�@�N!���7qR9��f�~��     �����ӦM��+WƊ+b�ĉA1��´f`�˗/Ǎ7� ����g�}�~�i��rR9_�N�555��� ��      �� R�aÆشiS,\�0k%Z[[�|kjj
���9s&-Z�gwr��ٳ����ʍ���I�իW;�<Ƥ�)r�x�b �p�B���9�     �zzz��V I��:;;�'M�����b���� �C���:uJ�N�	�ɽs��<�k׮e��7oޜ����[��^�T�ї6dw`���[� v֬Y     �WK��� 8�_WWW6�=�mmm�P@߿��x7�Pwr�w��ݻw�zR9]�bŊl���	��cC<HZ��     ����&i���]�����%
��������6y���ӝ;w`��~�@�N���p�t�RvR9Mv_�pa��kmmF��xk      �o&r�Q�!S�Y�~},]�4֭[3f�ƦJ��p��O`���糃/*�gwrO��p�����T��i[�jU6�}ܸq���b      ��R�����;��{��7o^6pѢEQ]]�-�������e�s��	�+�;�v�֭���OF�ŋ��c���[����W��Y�f�+m�ҩ����  p     �z�;V�+�#�;v,{b����`�)S�c������nw�L�N�]�p!`4���d'����Ғ�Tnoow��0����6�׮]���Q�@-�     �ˮ\����p���زeKlݺ��S�/^UUU��ijj
��H�	�ɵ��hK��ҳaÆ����6pN��t]N�s��<�A�a��!Zccc      �e�6����ӦM��+WƊ+b�ĉ��Ө ��"���	�%������cǎ��SOeWr-Z�(�����w�������ȑ#�f8� _%��      &pg�]�|9�iӦX�pa6���59i�{��:< `@�	��5��҆�����3iҤ�r��M�2%x����СC�k׮8z�hܽ{7 F
��ϟ      |�魌�������̞4Q���#k%����5nܸl(ا�~ ����Ν;Q[[�GwrM��Xw�ƍؼyslٲ%0�T�DUUUY���Ķm۲S� ��Z      ૝?>`���2MuO�D[[[�^�:f͚�t�@���ח5---y$p'�Dm�E�P~����<yr�\�2{�����7n�+W���e-      ���m�0Zzzz����3gΜl(�ҥK��F�6�nݺ�Mq�_Z��+�r+]m��!y�~n�~��x��wc�ٕ\���Q�T�Ҥ��^{-�= ��ҥK     ��������c��ӧ��7ވ���,v�6mZ��]�G��cǎe�N�S�WqЍ<��[W�^ͦbC^ݽ{7��ߟ=iӖ&��X�"&N�E��fq��۷`(�     ���M��
ƚ�7oƶm�b����0����UUU�WK��޽{㣏>�S�N��<������[i
4E�yްaClڴ)�,Y�Mu�;wnE�q��C�ٳ' �R�F�UWW      �3���,�����466fCӓ���ݸq#;�{������G!p'��䖉�Q
�Ӊ��477g'����c���W�������Z,����חE�/     �"Qyq�ڵl �ﾛMsO�D��^�T��zzzb˖-�s��lz;���y&p'�Lp������_�7�|3�����i�'ׯ_����������pIk�;     �	�ɛ4���?Ξ��_��bŊ�8qb�ɡC���^�}<�4D��ݻQ]]�7wr�w�"Mu���̞����r[[[�7.Ʋ������?����:     �e�g��wÆ�d��|Tw�܉�7Ǝ;`(��C���>}z@��ɭ�W���ٳg����}6ս��=�ݛ��c��y�f�����^k      �L�N
8s�̬�H�D]]]ɥK��׿�utuu�P��Wwr�ڵke�����^�����r����֎�?Z����o~�p�B ��tc      _dHEs���x�ײ��˖-�b�Y�fEޝ8q"����;nݺ Ć7�J�Nn	��4�==�ׯ��K��ڵkGu���o�G�	��bM      �E)�M�Ӡ�zzz���s�����������?��?q�Ν w�J�Nn��
_�>�صkW�<��Y�hѢ�����C���͛`$Y      |�����P��7FGGG�755E<x0���޽ �Ś����K)�}�v v�ԩ�ihh�+Vd�ɓ'���駟�+�����0�Lp     �"�Z)��7oƶm۲g��>�3g�������ہa'p'���I��pҟ�w�}7��>o޼,t_�xqTUU����?�1��`�Y      |QPe50���1V�\�=�Ǌ����Wܹs' ��իW�H�N.	��Ѥ��ǎ˞4�}���z��!��~�ȑ8p�@ ���.H�s�J%      p.$����M��w����+Ml��o~c� 0b�	�+�;�t�ƍ ���nٲ%��k��ٵ\i#�m�����lz;�hIuwwG}}}      `p 6x(�iӲ��+V���'��?��������0R$����͛7x<}}}q����ijj�U�Ve��'L��H��֭[�ҥK0���@�     p�i��`�/_�6d��.\�Mu�����СC�s�� Iih`j*F�P<�;��Z)P�7b�ƍ�������۷�h�6      ����^�����3{fΜ�loo����a��������o�)� #-Mq��7wr�w�7pӧO����,v������~tww�h�6      �\
ـ�s���x�ײ��mmm�z��5k֐�o����4�Q����7�;�dJ+�����^˵t��X�n]̞=���{���������A      ��ãK���ڵ+{ZZZ���i�{mm�c��.\�~M��b]@	��%��4���?̞�ܲe�b߾}���k     �����ٳg�g����P��k�Fss���^�������b]@	��%�at����x�k     �{��t#7��������w����X�jU,\�0���������ĉ0���:�\�}�v �'m� �k     �{Dl0������ѣ�3iҤ����b�)S�|�߷u�� m��GwrI� v�Ν      @���ƍ�e˖,^�7o^<�쳱x��/Mu?y�d�9s& F�g�}�7wrI� fm      p��FF��~�ر�6mZ�\�2V�X'N���m۶�X`�;y$p'�Dl �`�      ���`�]�|96l��6m�%K�Ă�СC08�F	�ɥ;w� � k     �{�������w���+��#�;�dJ+ 0��     �=�7 �6 ���R:� 0�w     �{Dl �`����\��� ��      ��� ����#�;�$b �6      ��ͷ �`w�H�N.�� ���      �� �Y�GwrI� fm      p�� ���7����R����\� �Y      �s���  ����UTWW���\J/�  �      ��� �������K��; 0�5Z      ����Y�7wrI� VUU      � �/�{�n@��ɥ�ِ �      ��) ��(L���% 0��     �=w �~&��7wrI� fm      p�	� ���#o�䒈 ��      ��J�  ��*��;�T]]  �      �� ��> o��RM�] �s���     �� �2��F%L.�7.  X      �S�T `0�;y#p'�Dl �`�      �TWW �`����\� �Y      �cB+ p?7��7wrI� V[[      ��
 |Q�ۭ��;�$p �6      ��`  `������;�TWW  �      �1 �ڀ<��K&L ��      ��� &p'��䒈 ��      � 0��y$p'���� `��     � 0��y$p'�� �`w     �{Dl �`���y#p'�&N�  ~     �g��� 0@SA	��%/� �`&�     ��{ `0k�H�N.544 @�����X�     $"6 `0��#%����  �u     ��� �`����\�4iRT*���� ���      �3� L�N	�ɥ���,r�~�z  ����      �SWW�u}}} ��y$p'�R�&p Lp     �\�R�&�޸q#  Lp'���V��Ξ= @���     �E���; �H	��-/� @bM      �E)p?w�\  H	�ɭ�S� ��i�     �� �. ��䖘 H�	      �H� $UUU1a����[&� �5     �544 @:�V�T�F�Nn��
 ���9i     p��ġ7�J�Nn��
 8�     �e�'O  k�J�NnM�81jkk�Ν; ���     �� ]y%p'�*�JL�>=Ν; @9��       _$f ���+�;�6c��; �XZ      �E&L�������	 ��z#���Zsss  �e-      �`ib�'�| @y	��+�;�fj+ ���      ��	� �;y%p'�Dm P^�J�Z      �+� ��RW1eʔ�<��k��� �Sڄ���      _6}��  �+u552a��O.���Ԕ� ��� P.��     |5C�ܬ�3�;�VUU���={6 �riii	      ̰  (7�;y&p'�R�&p��={v      �`3g� ��v#��䞸 ��w     ��6~��hhh��ׯ P>w�L�N�	����      �^
�� PNw�L�N��
 �3iҤl�      _m֬Yq�ر  ʥR�Dsss@^	�ɽ�"\SS��� ��n      �,� @�455E]]]@^	�ɽ���lCv�̙  �aΜ9     �כ={v  �c@�	�)�'�|R� %��O      _ϭ� PN� ���B0� �%n     ��555E]]]��� P&��ww
A� �QSS�f�
      �^�RɾW9y�d  �!p'��B���6e��� [�F+E�      |��	��<RK)p'�AB�Nkƌq�  �-l     ���Vv�� @9477gM%���;w�� J��'�      ��V �\��Ƽy����� ��Z[[     ����J���� ���"�Sb7 (�q���O<      <����GSSStuu P|w�@�Na�嚚���� ���ΝUUU     ��KS�� Pw�@�Na��=mȎ; @1��     �ѥ�b��� ��ɓ���1 ��ʼy�� P`�     �G�n� �逸�
(�;�"z�b�^     ���w,�J%��� (.]E!p�P�y�  ����9�L�      <�����5kV�;w. ��jmm(�;�2y��,~�p�B  Ų`��      ��I]� P\UUU��SO����I�� ��M-      �^
ܷm� @1���D]]]@�)��oݺ5 �b1�     ��kmm ����S$w
�tW (��S�FSSS      ����Ǐ����  �'��E!p�pR�6mڴ�|�r  ��      �㩪����~::;; (mE"p��-Z۶m �/^      <�����N�ӧO(
�;��d��; H:�     ��1� ��{<E#p��Ҕ�J���� �[KKKv�     ��3w��7n\ܾ}; ��H��@��)�I�&�O<�O�  ���,      <����hmm� P&�S4w
+Mq�@���t      �F��*p��hll����"�SXi��o� @~�)"��     :i�Ы�� @1���J�P$w
+�p�Ǐ����  �)�����      Cc޼yQ__�n�
  ��0`(�;��&���I|�A  ��lٲ      `�TUU�cϞ= �[�ܞ:I(�;���8�; ��     `�N� �����'O(�;���ޞ�P���  _fϞ���     ��Z�dI  �gz;E%p��b�ܹq�ĉ  ���v     �ᑆ555ťK� �/��(*�;���8�; ��     `���b6m� @>�7.�y晀"�Sx�ꫯ �'N����      ã��]� 9�x�⨭�("�;���O�̙3���� �C:�VUU      �����㣻�; ��I��@Q	�)�ɽ�� ��ʕ+     ��SSS�-�={� �/�JE�N�	�)��	� &L��}�
     ��Ja�� �gΜ91eʔ���S
s�΍����t�R  c[{{{61     ���4���? ��0���SQ
i3���7n `lK7�      0�&O���͋cǎ �+V�(2�;����
�`�?~|,Y�$      i��� �c���1gΜ�"�S����{WWW  cS� ���6      �����������;���?��a���c AD���QA0"���hS��[�&�$�MbV�ny$�dc��^+I���w<QO0FQ��>_�嚣g���z����-���3���TUU ��Ұ_h��䍂��2dH�q� 䦡C�      ��u�����_= �ܗ6�AC'p'�TTT� G�h�">�O�  n�IDAT��      �v�PN� ����,�t���	��+:t�N�:Ŋ+ �-餕���      �v80n��  r[ڔVPP��	��;C��@J�;      ��}��@=p衇��;y'�i��m� ��ڵ�8       �@nkݺ����!p'�EϞ=c��� ��Ç;B     �����o����  rOEE����!p'/��N� �!]|6,      �;i`��K�.  �2$ _��K�f͚���� �[�{��~`
     @�JS�� �{:u�;v�w�RqqqvQv�=� P���*      Խ�����Ɩ-[ ����o���	��n���f'�      P���n���O>�d  ���� ***����եK��ܹs,_�< ��1lذ(*�      W���w ��{������|�&"�~��q�u� P7F�      �C9$��g�x�� �{i���;y-�q�7Ć �]tPt��1      ����YO�hѢ  �Viii���? ���k%%%1lذ��{ �]GqD      �{�)�w �{C�����|#p'�5J� ��E�1`��       ��������J  ug����H�N��СCx���lٲ  jǈ#���GQ     �\UYY)p�:Թs������בG)p�ZRXX��@     ��5t�����~�ׯ ���5* _	��4(��w�x�w �Y�}�M�6     @�*..�aÆ�]w� @�jڴi2$ _	�!>�$�v;���� �f�3&      �}GqD�}��QUU @�I��JJJ���Oeee�v�m�q��  jF�.]�[�n     @�k߾}���#�,Y @�9������O�f͢��"���  j�رc     ��#Mq�@�I��:v�����	�G������Z P���bРA     @��~��~ϳf͚  j^�!�	��:t��rH<��� T���:*5j      ����1jԨ��� �Y�[���;�;��c�9F� լY�f1r��      ��9������o��7 Ps�<��ls�;�;��8 z��K�. �z��&M�      �OfTQQ��{o  5���$F���vh���w �&���ٱ�      �_GuT�w�}QUU @�>|x�������7:w�˗/ `�92Z�l      �_���ѻw�x�� �^1z�� >"p�Hocǎ�+��2 �=רQ�l�      �߸q�� P�ڵ�#w�C���n�-�z�  �̰aâM�6     @�׳g��֭[���� T�����ww����q�1��UW] ��K�G}t      �p�;6.��  �G�^��K�.�����СC���o7� �@����,     ��e���ѡC�x��7 �{���g	���ɳ&L����: �]gz;     @�TPP�Mq��/~ ���ܹs���3�O��NTTT�w�a�; �4����<      hxRKq�-�Ě5k �s�sL�y�4�;�D�@��D���  v�Q�F�{'      SQQQv����  �Lǎc���|��vA�y��?�!V�X �9rd�m�6      h��������w �C�&M2�>��vAz�<yr\r�% |����0aB      а�)��Ǐ����7 �:��_@�����ѽ{�x饗 رѣGGYYY      ��UVVƝw�i�; �c�=��v�w�S�N���� |VӦM�)      �S�`�u��1����n�ѣG���;/^ ���7.JKK     ��������U�V �s�'O6�vB����㏏^x!�m� �GZ�jGuT      �_���'�5�\ ��ҥK0 �/&p��ԩS�8��� �#S�N�ƍ      �gذa�hѢx��7 �|��0�vN�{�㎋�<6l� ��:w�     @~*,,�ɓ'�e�] �����#z����	�a�l�2Ǝ��rK @��>}���      yn���q��+�� �gM�6-�]#p�=4~������c͚5 �*���gϞ     @~K��L�?�� ���Wt��-�]#p�=T\\�w\\u�U ������b      >֫W��۷o<�� |�Q�F1u�� v���BEEE6�}�ҥ �f�رѮ]�      ��N8�X�xql۶- ��Q�FEyyy �N�{!�5s�̸袋\��W���b	      �Ծ}�9rd�{� ��Y�f1q�� v���R�Ν]��w�O�%%%      �h����裏Ƈ~ ��R�^ZZ���C58���'��>�  ��;��c���      ;ҢE�?~|�t�M ��m۶1jԨ v���A�a5eʔ��� �F���'�      �g�ر����ʕ+ ��	'�EE2]��s��TVV�C=/��R @Cu�QG�~��      �ER�7}����K �M�^������;T�4�v֬Y�����u�� ���u��1q��      �]�¾�}�Ƴ�> �/�&��N:)�='p�j�&ڎ3&-Z �Мx�QRR      ��fΜ/��Blٲ%  �����<�='p�j6iҤx�'bժU š����      ��ڵ�B�;�3 ��kٲes�1��;T�ƍgǋ\|�� AӦMcƌ      {b�ĉ��#�Ě5k ��W4i�$��#p�зoߨ����~8 ���>}z��>      {���$fϞmX  Z�>}bȐ!�=�;Ԑ�3g���?k׮ ��z��#F�      �iX`���㩧�
 hh���㤓N
�zܡ����f��/�� ��h�$����      ���¿_|16l� АL�81ڶm@��CJ;��?�x @}3u�T_      T�����4iR\�� EǎcܸqT�;԰�O>9�,Y��~ @}ѭ[�5jT      @u=zt<��#��k� �w1{��hԨQ �G�5�y��Y�~�e� �%%%1w���"      �Saaa�r�)���~7�l� P���[ݻw�z	ܡ4(F�<�@ @�;��]�v      5�S�Nq��Gǭ�� P_�n�:�L�@��C-�9sf,[�,�z� �\էO�9rd      @M�8qb<������ �71gΜ())	��	ܡ��7�y�������غuk @�i޼y�z��E      Ԥ���8�S������z���2z��@��C-�ҥK{�q��7 �Y�fE˖-      jC�Νcܸqq�w �eee1mڴ j��j��G�/��K� �#FĠA�      jӤI���矏W_}5  ���ٳ�iӦ��;Բt�ּy��_��_b��� u�]�v1cƌ      ��֨Q�8��S㢋.�M�6 �ѣGG߾}�Yw�鈒�����/ �KEEE1��hҤI      @]�СC����_�:  W����S�P��PG��� ԕ�ӧG�Ν      �ҨQ�b�����SO �����đ��� j����I'�˖-�իW ԶtdV�A!      �9s�ī����^ @.�4iRt��5��!p�:Դi�8����G?�Qlٲ% ����q�i�EAAA      @.hѢE6��?�iTUU �=z��G@��C�֭[�p�	��_�: �64j�(�`UZZ      �Kz��Gyd�u�] u�Y�f1w��(,,���!�5*^{�x�� jZ�Xս{�      �\t���ǒ%KbŊ u�K_�R�n�:��%p�q��'�o���� PS=��l�      䪢���7o^\t�E�y�� ����0 ��'p�Q\\g�yfvq�� T����3gN      @��رcL�:5~��� Զ�>4}�� ��rH:���N��/�8��� �K�&Mb���-      ��G��%K�ēO> P[JJJb�����Z�n�!����'&O�7�|s @u(((�SN9%�]      �E�=�ܹs�{��^��� ���O�:Pw&L����z��/	 �['N���      �7���:+.��ذaC @M:��#cذa�-�;䠴��SO����ov �W����{l      @}U^^�Mr���UUU 5�k׮1}�� ��rTځ�`����w�k2 {$����N�6N     @}6`��;vl,Z�( ��5k�,�8�(*��B.�9�}���$��.��d vKiii�}��Ѵi�      ��`�ԩ�bŊX�xq @uI��͛mڴ	 7�!�80�L�7�tS ��hԨQ̟??��      Eaaa�~�������z�� ��0mڴ�۷o �C����	����/ `gN<���ٳg      @C�N2NÞ~��Ė-[ ��СCcܸq��;�'�tR�\�2^|�� ��3~��8���      ��]�fC����� �=թS��3gN �G��D�F���3ό�}�{Y� �h���1u��      �����2^y�x�� vW�-b�Ѹq� r���t��W������k׮ �.M��;wn      �Y�f��o�K�,	 �Ui��g��[� 7	ܡ�iӦM�s�9��(6n� жm�콡��$       _�@q����}/V�\ �3ip�)��|p �K��P�.]�d�\rIl۶- �_�Ȭ/���-      ����8������~�_�> ��L�0!�@n�C=u�!�dGm�� �S�ƍc�Ѯ]�      �|վ}�8묳�'?�Ilٲ% `G�'O �	ܡ9rd�Y�&n���  �řg�ݺu      �wtP̜93��� �t��i���>�;�s�&M�M�6ŢE���PXX��zj���7      ��~����;��w� �]۶mc�Q\\@� p�`ڴi�aÆ���{��-�$�5kV2$      �O�2eJ���{��� 4o�<�=��hٲe ����;�|�ɱq��x����k���1r��       >+5�g��"��{. �_ib��g�����/wh �ک��[�n��{, hx�N�GuT       ��Q�F1����˗/ �Oaaa�~��ѭ[� ��;4 �My�ܹ�$�g�y& h8�=��8��      ع&M�Ĺ瞛E�+W� ����<@�$p����(�<����OK�,	 �ѣGǤI�      �u��O|��_����z��  ?��1bĈ �/�;4@���q�9�d���e���k���1cƌ       v_YYY�w�y�$���{/ h؎;�;vl �������,r�����믿 �?��9s�dGg      {�]�vG��֭ ���:*&L�@�'p��iӦ��/9~��śo� �)n?�3���0      ��ӱc�8���A��ׯ �#�<2N8� �;4p-Z��o|���$^}��  �2$N;�4q;      T�Ν;ǹ�?��c�ƍ@�p�a��̙3h8��5k��u���K/� ���ʘ5kV      P��u�.����g�y�� �~4hP�r�):h`��}۶mU4hM�6��|�+q饗���? �Q�Fŉ'��      jPϞ=�3Έ�.�,�n� �O}��y��Eaaa ���}[ ^III�s�9q�WēO> ����Ǵi�      �y�����O?=k(�S �Oڬt�YgEQQQ O��]����=�B���+��� �V�֞��q��      P{_�җ�k���#|p,\�0���h���>�AI�{څ�&�?���@�Hq��3b���      ԾaÆEӦM���/�-[� ��o߾�`�q;4pY�m�6�!��)���]���O
 jWz�3gN><      ��ӿ�8묳��?�yl޼9 �M��z���ـW�a����yh���&M��m�� Ԏt�5o޼��C      ��_�������cÆ@n:th̝;7(4|Y�y�f��@�<yr���č7�UUt �IiSQ�MܧO�       r�A�~���?�u�� ������O>9�
�,pߴi�������m۶q�W:n���l�2�9��ҥK       ��k׮Y�����$��� �n��m�ԩ�v�3Y�q�F5+��V�Z�%�\�"���k�.�=���      �]�;w�����o��o��� u#��ӦM �l��.p2ݺu�/�0.������� ��ںp��hѢE       ��}��q�d���U��ړ����1v�� �S�oذaK ��6m��7��l���e��=7x���;wn      P�~�k_�Z��\�2 �y)n�5kVTVV����}�ƍ&��RZZ�~�����~8 �}�G��3fd_      @����ƅ^�^zi,]�4 �9EEE��C=4�������� ��?0�m�6n��� `פ��ٳg�a�      @����w�yq��Wǣ�> T�f͚��G��=p� ;��O�4)Z�n�^{mlݺ5 �|�[,��:(      ��!��7o^���P�R�v��F� ��w�}wc |��ÇGYYY\q��nݺ �:v��&N'_       ��!����կ~eH @5�o����=��l�}����Q�F�yz����ַ��K/�7�x# ��~���i��M�6      ��9rd�j�*.���ظ�\Q�=շo�8�3�I�&�IE��|��Ѽy� �"i*�7��͸���'��|��4�7.�N���      �e�~��/�5k� ����2N>��(,,��q�~�z�;�KJJJb����hѢ������* �Q�A<w��0`@       �e����/�0~���������KA��3��#����q�nݺ �UiJ���㳋�+���k�w:v�,����       �S�V��.�+��"�y� ��A���~zr�!�E>�׮] �+����|'.���x�� TTTĬY��-      ���~o�p�¸���㮻�
 >+<묳�C��3w`�����׾����\�ZQQQL�6-ƌ       ��̙3��_���y�� �#i��y�Y�f�+>���� �S)��~�v���ƍ�!�w�}c�����      ��:4�N|饗��ի �ĸq�b�ԩ�}�]e�;P�҅Z�.]�+���˗@C0p��8�S�$      v�s���o}+.���X�dI 䣒��8��ScРA���@�+//�/�0n�ᆸ���* ����l�1c      `W�h�"�?���馛bѢE�	 ��~��3ό���/ ��ǁ�{� ե��(fΜ�rH\u�U6� �N:6��3�p�      ���6mZt��-���X�~} 4t�/}�KѴi� �S�k֬	��ֻw��������+��_�\WPP�F���?>��      �7�غ���cŊ��M=�w\�?> �ƺu�����m۶�E�:�j�*;v���������iӦ �E-[��9s�D�~�      ������7��͸��⡇
���u��1���ڵk �w�y���֭[c�ڵY�
P��D����8���i�z �A�ŬY��y��      P�7ns���n�򗿌?�0 껁f�KKK�:|*p�����I�ȭ/�0n���l��# �R�&Mb����&      ��6x��l������/� �QqqqL�:5ƌ �i͚5��� 5�Q�F1iҤ�ݻw\s�5��[o@]H�Ci���       ��u��q��m�ݖ���� �/Ґ��O?=:u� ��3�W�^ ��{����|'n�����`�;Pk�6m�|�92


      ��f8��l@�ڵk ����#���ӧg�j�g�U�V@mJt�M�C��.֖/_ 5�o߾1{��(++      ���~������q�u��_�� �E-[��9s�D�~��&���۟�W�\ u�s��q�f�n�y睱u�� �N͛7��3g�СC       ��h�",X�?�x\{�~�� ��ʆ	���@MK=���EEE1eʔ6lX��W��^x! �V:���";+�P       W<8�v�W_}u,Y�$ �R�&M�ޢ��2 júu벍~�
��y�زeK�ԕ���8�����믿>>��� ��ڵ��O>9z��       �A�֭�_�j�u�]q�M7ŦM������7��^VV �����n?U�WUUŪU��}��P����4ɽw��q�7d�{z���5���:*&O�l�      P�nb̘1ѿ���//��B Ԇf͚Ŵi�Lm��ʕ+�ۢ}A�䊖-[�ܹscĈ���&�x� �"iZ�̙3�C�      P��i�&�;Ｘ����w��]lذ! jJ�~�b֬YѪU� ������ً@.9蠃����v�}��q�-�ć~ �Զmۘ:uj<8       �4�=MR�ӧO\w�u���@uJCH�0�C=4 �R�ؓ����_ f�o6,n���,v���
 �5n�8ƍG}t      @C���ƹ�O?�t��W��5k���Hh***bƌQZZ um{Ǿ�	� �,}�J;��_}������Y�w\���      @>�ׯ_���#���+��ضm[ ����/f͚ݻw�\�>Ӭ\�2����=MDN�@.�֭[|���v&�������~;������O��"      �KM�6�x8�u�]+V��]Ѹq�8qb�;65j �⭷ފ-[�d�?�oڴ)V�^mڴ	�� �L�ӧO�+��[o�����0�k�.��>h� ��      �����}��ߎ�~8������������O�֭[@�ICڷ+����׿
܁z%�&3fLTTT�����{ol޼9���e˖q�1�Deee       I����rH60ܶm[ lW^^�������ԯo��B���_�v� �7͛7�3fdG��v�m���h�z���$F����M�4	       v���4X;���o~/��R �-u���0a���@�[�|����v������,fϞ�}@K��Q\UUU��*��eʔ)ѢE�       `����q��O<����cժU�t�CEEE��Ѳe� �Ҁ���@���י;wn�3&;��駟�C+..����?~|�j�*       �})n<xp���/��l8��h�z��ӧO�N�:@}�~��X�f���a�z������y������.�7�x#n��l���r�����{��      ���!ci�؈#�^�{�m۶��t��!��~�!�@}�����,��'�)�i'@C��~������}ѢE���ݡ	�      j^t:s��8�����o�'�|R/D�֭cҤIQQQ���P����>7pOO�U
��Ν��R���;��G��[�P;�4iÇϾ��       �#Mx^�`A����D���~:��)m\7n\�=:;��>K��?�s�W^y% ��;f���ɓ��c<���q�� jF˖-�� cƌ�f͚       ��k׮q��gǲe�⦛n��K�P?���ĨQ��c��4/����,p����IGqM�81����{�>�z�o�>ƎÆ����       ��x�����=���,tO�݁ܔb�#�8"�>�hC����ߏU�V}��-��}��X�fM���@�HG�L�4)&L��=�X,Z�(�x� �L��ݳi�����        ����+[)t���G�"l��ޞ|��� �&M�N���J�q�u�]��%�m��K�?�zh�7.��o�       �~��?��q�m��08jGiii�=:,شi� h�v������@�K�q���[o�����ğ���X�~} �ֶmۨ���#Fd�!       P?���7[i(��w��<�LTUUP�Z�l�~xu�Q�v /��w >R^^3f̈iӦ�SO=��w_v4䳂���ٳg�80
      ��a�P�+V����x�Gb۶mT�4X��#������� ��s�k����ǿ0pOaӦMѸq� �#EEE��i-_�<���裏Ɔ�ž��Mj9rd�j�*       h�:u�s�΍I�&e������ظqc {�G�ٴ����g���믿�����-[�dS��dV >�s��1{��9sf<����T�^x��\4HisG��6lXv�i�       ��M�6q�I'�ԩS��?��O�z�� v��#��ݺu�|�dɒ>���{�t�R�;�N�c��Ou_�jU�S9-q4]�v��Çǐ!C�Y�f      @~kҤI�3&F��<�L�u�]�����Ś6m�vX�7.��� ߥN}Gv�^������H��^{�x衇����k���[��C=4F����       ���� ��뗭7�|3���l��ƍ��.]�DeeeTTTD�ƍ�����x饗v����Jl޼9�N��IN�:���_�b�'�|26l��kZ�j��N"�޽{��       �:t��3gƔ)S��G�{�'V�X���IC��#�8":w� |�o��֭���v���=E�tP �g
�W�^�J���X��<�z�����J:�o߾�n�t���      ��JQo�T�ֲe�����'�x�Tw�F�n�b���1t��())	 v,�<;ܓb
��G:c��\۶m��_~9��{�X�vm@Mkݺu���ߤv       jԁ��Y�f��O?��w_���QUUА���ƠA�bԨQѩS� `�}�����.�/Ύ��z�i��/�N8�X�|yvA��3��k��Pҿ�t��!��m����E�       Ԛ40aK뭷ފ?�������;�P_e-�a��ݦ>�]�y��X�t��~}���_=֭[��2�f��]�t�֤I�����B���#��:���ݻw���o߾��      �	���q�q�e+�{衇��G���? ץ��ݺu�6kTTTD�������/~a�K���m۲�aҋ2 ��m۶1z��l���?�����q�x�.>i����={F�^�⠃�F�       �� �O��/�Gy$�aÆ�\����]�Ɛ!C��C�}��' �;�>��~}��$E�w�����J�rZ�ڵk?��S��r�� �l�{��E�)h/))	       �o� �tByZi`j"R���O��N�HQ������L��۵k T��{���ˁ{*�Ӵ���@�jٲe��9�$�K�.�b��^zɄ�h{�޽{�8����͚5       hH��~��e��O�_|1�x�,xO}Ԕ��"8p`�Lj�i��Ά��r�f͚X�bE��[R�N��~�F:��W^ɂ����}ݺuA��.��1li7p
�S�޸q�       �|QTT}���V�׿�5�y�xꩧ��_6���VZZ={��xS�a� 5/]ߙ]ܓ��@����4i�M�N+It��߲�=�˗/�6-����6(��״R�~�DYYY        ױc�l�?>�}�ݬgK�\�����LAAA6l�w��YО�� �����sv+pOǼs�1@��>�w��![Ç�K���o����)zO���Z�z��5$�,o׮]v�ݩS���vGZ      ��iժUTVVfk۶mY���/���?K�.�-[�$i�`�=�A�)j�i ԝ͛7ǒ%Kv���
�_}��X�vm��@����[�5x���ߴiS����J�{���B��қ;���j۶m��v�Ƃ��?       P}���Ӊ�i����D�ϥ��˖-������6?t�AY�~��Gyyy ���sjwf��4�7�}�/ O�ƍ?��������J��ʕ+���;�|��{ｼ�,..�����w�}��6m�|����͛       P7�4i�M�N+I��K/��MvOa]
��k8R�ѽ{�����n ���{�]z�n��O<!p�Ci�{���J�(��)rO���5k�����V:�#���׭[~�a��ߗ&��h��㕎�J�z:�$�O;|SԞ�       �)x�ӧO���8��S��&����kٟ��?r[IIIt��)�x��f����xꩧv�y��/^�8�KKK �K�}m�w&]��}����Ziwt:~d�ƍ�u���9�o?i��?)MUOk��7m�4������4�>�O�����o_�b       h�R�бc�lUVVf�}��Y�|��W:�^�^wRϱ���G�Ν���o�>kB ����U�v鹻�����'��#F ���޽YU����c} �����$jlJM|%F�ֶ��M��δ��&M�S'�tҙ���bZQ�5���@�"��G��օ]XvY��.��۞�BMb"�}�{��3�s��=砻�}��ږ�       �PK>���[��\.�x�hjj����ؾ}{zL>Ş��,,L�����~�A��z�@�X�r����������         �����'N��Λ%�ޓ�}ǎ���;w�L��'[i�O�筍;6N?��ÓD�g�}v�v�i�V} J[]]�������ק�B;餓         �E����.H��
�Bttt��{[[[�޽��$�'�8p JQ��|�����$dOfܸq�ׇ���Ç �)�4��MaG��|>�V�W]uU         @����8w�&]]]��ٙ.�ݳgOz<�8�������><�\.�BUUU�=���5*��IB�d���'3lذ ���r�ʣz�1��˗�        �UWW�3~��#z}��P���חｽ��$��e��^��%�9�~��d���M�#G�L��$^O��#F��O��m���t�G������]c��rJ          �+�
h�: ����hii9�s�9pO��UWW�\sM           ��-[���9��=����          �f�B�+V�y��oڴ)v���ƍ           H�_�>:::����
ܓ�>��~���           $�.]zL�W��X�xq|������           ���߿?V�\yL�w����7n�.�            (o���ӹ��'�-�w           �,Yr���K�����ԧ>���          @yjll�m۶��������k�?���           �i����u~��E�	�          �TOOO����u�~ܷo�1a           ��$q{.�;�k�[��H���          �Oғ�~ܓ���o�ѣG           ��7ވ����N��i�~��W           �?��'�5pO���+q�UWEEEE           P�zzz����_���{SSS�[�.���           �m�������/����=1o�<�;          @����`��~�ހ�?���c۶mq��           �iŊ�k׮~�ހ�_|1n���           �4͟?�_�7`�����S�L��c�           ����>^��~���}}}��K/�'?��           ��̛7�߯9`�{b��O|"F�           �����X�zu�_w@�\.K�,�뮻.           (s�΍B������=��/Ƶ�^Æ           ��޽{���v@�=��{{{{�X�">��           �m�����; ���=��/�����FEEE           P����.��J���Ԕnq����          ����/FWW׀]P��̙3��.����           ��twwǂ������Ĳe�b���          @q�;wn��A����/�<����           �}���K/�4���Ҽ��-�.]��G          ����s�E.����*�9s���ɓmq          ({��W^yeP�5���ݻc���q�5�           ٖlo?p����kH֨?��q�W�	'�           dS��|ѢE�v�!	������          �lJ��<xp��7$�{��矏�|�#1r��            [v��?��O��C��ݻ7�ܧL�           dˏ~������{Y���7o^\q�q�g           ٰaÆ�����i�~��������o�=           z�|>�z�!����_�n]L�4)           Z�-����!����������          ����3g��3�777��ŋ㪫�
           ���ٳc߾}Cv�L�g�y&>��Fuuu           0�v��/����2�wuuų�>7�|s           0����+�����ߐ��=�`�����?g�uV           08֬Y��P�T�����G?�Q����m           0�����,�T��H��������K          ��5w��رcGdA����?^xa�=:           ���1gΜȊL�QSS����          ��W(������ȊL�ŋ��_]tQ           п�f{����%��������c���          @���쌚��Ț����֘={v�t�M          @�x��ǣ��;�&Ӂ{b�ܹq�e����           �U�VE]]]dQ��|>������O�Æ           �M.���{,�*�{���)�ϟ�_}           pl�~����般*��=1k֬��K�3�           �N}}},^�8��h��������aÆ           G���'}��(
�eE�'�瞋o�1           82�=�X���F�U���3gNL�4)&N�           �v+V�����(E��������_��c�ȑ          �[koo�3fD�(��=�k׮x�'��[o           ~]�PH��wwwG�(��=�t��x�{��Ї          �_6gΜ����bR��{�����'Ʃ��           �-[��g��bSԁ����ӕ�������          P�zzzb������Ŧ��ĦM���矏?��?          �r��ODKKK����gώ/�0&N�           ���W_������bU�{�:ڴiq�=�Ę1c          ���ر#f̘Ŭ$�Dggg<����/|!��J�?          �m�r�tixr,f%U�o޼9jjj�[n	          �rP(�?�Al߾=�]I�����y��'O          �R��s�E]]]����3f̈��>;�=��           (U�֭�Y�fE�(�����7���o�=�����          Pj����{��^���(%�'��~����������          �R�,��w����RR��{bժU1gΜ���          �T<���e˖(5%�'fϞ�x�;��/          �b�p��X�dI�����B|��ߍ��+�=��           (V6l���z*JU��\.=�P��?�c�;6           �MsssL�6-<��,�DGGG<���q��wǨQ�          �X�ٳ'�N����Q��&pO$�X��w�w�ygTVV          @�����q��ݻ�ԕU��X�vm̘1#����<           �,������c۶mQ�.pO,Y�$�<�̸�           ��|�����~�,�ď��3fL����^           d�/�/��r�����B<��q�i��ĉ           +V�\�.�.7e�'z{{�[��V�}��q�g          �Pۼys|���O�z���������/��t�;          �Pijj��z(]�]��>pO������ߟF�cƌ	          �����<�@twwG�����;wƽ�ޛF�'�|r           �C=sggg�3���z��������          �������tttD��������:uj|�󟏑#G          �@ٻwo��{׮]���-���������>��1bD           �����4n߾}{���`���1mڴ��;����&          ���r�4n߶m[���ۿ�������������          p�8���7���1�e��QWWӧO������aÆ          �����I�������	܏�����_�������Ç          ����S�FCCC���Gh�������w�#G�          �#�w��x��b۶m�o&p?
�� �w�}�w�wQ]]           o���3퐛����N�~������}�sq�'          �o��֖�ǭ�������[��׿�����?cƌ	          �_��Ғnnooo����m߾=����������i��           �$�q�����#8r��k׮��7��F�g�qF           lٲ%x�����
����8�޽;��~�w���          @�Z�vm<��Ñ�傣'p�����&��n�->��          P~�,Y�=�X����F��Ozzzbڴiq�-�ĵ�^          @y(
1gΜ�5kVp|��(�����عsg�|��QQQ          @�:x�`���G,[�,8~�0��hkk��n�-N8�           JOWWW|��ߎ�7�C�>@^{���7�w�qG�|��          ��]�v�ԩScǎA��������W�w�yg�?>          �������ַb�޽A����_��W�����.          �x�X�"y�������}tww�}��S�L�n�!          ��R(b�ܹ���8}����|>555�������cĈ          d_WWWL�>=֮],�� [�lY477�����~z           ٵm۶�6mZ�ڵ+x�!�lq�������[�K.	           {jkkcƌq���`p܇H.�K��q����M7�          �|>�<�L�������B���ҿ��q�m���ѣ          :��|'��'pπ5k�Ŀ������g�}v           �o�ƍ���Gggg04����_��W��o�+��2          �������矏Y�f��:����3f�ڵk�3��LTWW          0pv���<�H���CO��Auuu�y����g?_|q           �o�ʕ�ꮮ� ����=�P|���O~�QU�G          �!����O?�-
�E5�a�B!�ϟ�֭��n�-�9�           �]cccL�>=Z[[��������򗿜nr���k���"          �#���c޼y��$����l�����x��'c͚5���~6N9�           �^[[[<��#�q�� ��Ef�ڵ����q�M7ŕW^          �[+
�x��x��#���'p/B]]]1cƌx�������bܸq          �����x��G���>(�"�f͚����������xTVV          �����x��c�̙q�����܋܁���&~����g>�?~|          @9jhhH��777�I�^"6o�_�җ�뮋?��?��*?Z          �C�4z���1o޼���A�RA����^x�X�zu��}	          �l͚5���G[[[P��%(�H��~��q��W��ܫ��          JI{{{<��ӱ|��t�KT�P��_~9�-[���Ǣ�ʏ         �����,�9s�DOOOPZ�%���;jjjbɒ%q�-���_          P�V�Z?�����-(M�2���S�N�I�&ŧ>��?~|          @1غuk<��S�q�Ơ�	��̺u��K_�R\s�5����1jԨ          �,ڷo_<����K/E>�J����������c�ҥq�7��{eee          @$���'?�I�r��|��XWWW<���ӟ�4�L�_|q          �P)
�lٲ�5kV�ܹ3(?wb۶m1u�Ԙ0aB|�������          �%	�W�^�nlojj
ʗ������fL�81��O�4.���          ���nݺ�����[���5�7o�{�7���wŔ)S���~w          @J��g�y&��mڴ)����ǤI�⦛n���??          �x$˘�����>�W	�y[ɻc֯_�^zi���Q�s�9          Gc�ƍ1k֬ذaC�o"p�
�X�re:�z׻�n����}QQQ          �V�u�����s�ECCC���s�6mڔN����k��ɓ'����          ===�lٲ�7o^���)�;Ǭ��)f̘3gΌ���:>�я��ѣ         ��w��X�pa,X� ������������f�J�a��8���7n\          PZ[[��_�W^y%z{{����~���b������/�<����x�;�          ��B��ׯO��5k֤_�����������6��������率�O<��          ���ٳ'�.]�nkߵkW@�3��o�5551s����>W^ye\t�EQQQ          �C��-Z���Z����Aq���X�bE:g�yf����+���N:)          Ȧ��������F[[[�@�3�ZZZlu         Ȩ|>6lH����ե_�`�3d޼�}�رq�e��?���0a��         `
�hhhH��W_}5:;;����Lhoo����3nܸ���K��}�ĉ         @���Ew2g��݇c�SO=5.���;         @?ٲeK��֦a{GGG@��ɴ���ñ�Yg����Ɍ?>          x{ɦ����X�|y����d������ܜάY�����y�{bҤI����7F�          �BWWW�_�>֭[�W�����!p�(%��-Z�NeeeL�0!�����E]�w^TTT         @�H��oݺ�pԾaÆ����F�N�K��nڴ)���'��nwO���8jԨ          (5���KC�$h_�jU�ٳ'��	�)9����t��t�����|g\p���w�;��>bĈ          (6]]]�q�ƨ��O�۶mK7�C)�S�<��O&1lذx�;ޑ��'NL���N:)          ����-bӦMiԾ}�vA;%O�NY���͛7�s�駟�nvOb�d�9�t�;         �`��r�u��4hO���_���΀r����ܹ3��������������8�����Ϗ��ǧ����         �xuww��طlْN���� p�_��磹�9��K�~~̘1i�~�Yg>&��G�          �*	ٓ%�I��t����v�
�	��utt��nݺ��UTT���g���駟�N����N��#G         P�:;;�`=	ٓimm=|ܷo_ GG��!�(����t6l��k�5jT�;6N=���8nܸ�x�'�)��'�tR:Æ          ;8�����ݻ7=&�r������w���� �ϡ�����_VQ���QOOO�ر#�ߦ��:�ޓc��}��ч'��G��F���UUUq�	'�����Ǉ$߷1        �r�,������璖/���������/r�\�'����$�O���+ړ��4;��笇.���{�ox�{��}����* (&�w�u��        8F_��ϫ���@Q�,�l�뮻FE�*            �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��       �v�X    `���4vG   � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �  Ԯ�6 �h ���T���,Sĕu�@�'pg���8        �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��~�y�_˲� �<ϗ       ��^��x <�i�~O��~Ǿ��[>         /c۶�[> ���           $��k����    IEND�B`�PK
     t$v[��n  n  /   images/6b551873-9f16-48c5-b1b9-2fc6ab10f815.png�PNG

   IHDR   d   �   +n/�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��io[U��Wl'q�fh�6miZ(P(C�2�|x��
�*\^!U�B|������ $�2�I@�g(3�<�i�$�<��ݿm/�4��Nb;��U�:�9�׸�^۷v�Z	����as�J|*0���o��Y�FNt
��[�1m_��?(}Q>P y�2�I�2��d��0��a�$�(H�Q��< Fy@2��d��0��a�$����SOɓO>)Ӧ�1���/((���By�g�D���!x������<�hKKK�u����TWWK �/�A�_��|�/F#�x�
JKK�D�U�V�=z���s���/���<���E�Ge}��O���.�����r�9�șg�)ӧO�_�F��2�O�W��ϟ�ɕ��Ef@���� '������o�m۶�P�%<���򴵵Y ���3g��2(�P]��G���zc�� ����<>묳���[��w�{�C���t�M�b�
��@;O�!� GU=����7�xþf��E]$w�u��D�y��C��}��7KGG�lذA|xW��8��8r�<��#5��z����_����eƌqՔ�� :88h?��,..��<����ò<`䫗
�U܈�***�ꫯ����� ���#�������r��!�wsB<1<�e˖Y`���O(�Q#�{�n��?d������ky?/^,K�,��<s#@����R,@ ��_��_]�9b_}e:�mٲE>��+v�^{�}�D�xs��ak�qaǒqi�o������n��.���%ڀ�u�A��5��������k�9��ڱc������}�Q�n�:9x�\��8�r����s�=g�ǢE��s���)���q�mmm%��}��ɽ�������NXTT$?������L��>Y�`���w#F�����+	ut��y��g���ώ�/�Ђ�:��h6���>��o=Z7�D����nG<����=�!?L�%}��6�d��ZL�qګ��j���[��K/����!��������vl�駟�7Q�~����|�r����~���	I���g>��SH���x��N;�4��#�@%�p�裏�w��~�Ao
�{@
���ᤵ��V7�L����%����#�i�&�=JJJ����'*͍0�dxq�4���@PI���f����I֯_oG<��t�RkS���c^4�sҪ���u�jµ�`��/�l@E�}��V:b����Μ93> �'F���h�y<b�J�g#�l��Ih
��~+555�����7�6�-k	����u��D�H4¦&��� �JB��ro�n3�%�C��`?�s�o"��ƛ��pR� ����ܹs�n�AG{�z�68�(()�� �� ��_|1a��#%�\�*� �u�1�\`A��W�w�6���'�������/�8���� F�HU�@�͛'W]u���/�]����\S'|�y�g�ډj���ґ�(#��P1�P)�}T���'Su�o�ݺ��[���<`y4��	�0��裏�+��"�y_7"2_�j�̚5+)ҡ �t�v��dp8t^�kU�G�hpL��<���L��c�=&/���͆�#�{T�Xj<f�#�?��CV��k�ڵ블	7���f`w��ɂSQ90~�޽6�RCc#��jj�#Xm���=��q4��xnj#⻤����P�H�XUI��95̡ǳ�q+u4�{�6e���q��o�H�����Ǎm޼�zy���n���M��&���ß�)�g϶G�~s���d2��kll��L��ʄ/'�tR��Od�&\J�?� 8/�c2�����n�߄Yc��t:�q�Pka�atõ��7��T�s�ZhH���x�sq�\+��)��r�{\�x4Ƹk{�m a8*f�ƍ�@j�NrdN�<���eV���5Sf�AQkF^yY��N�F���_::�䰑��C����Ez��#��B�0#Q�ؙ�J�+L�2���E#����Q�,np��`�a���e�YK�43�j���Q������2��2��a^
T�6��J�4̑�b����a���l���wȠyn%J�͇�3~��6͚�L�I�(3��O?ّ�TM#L#�/�@�_|�̬��ζViڹU6:(�248��Q���{
�WX$e�RS7S�<�t�	�ɮ��rd`� � �R���[���Λ�)��7Jf�:$5�j��������/)/.��[7��쐞��F�cm�S��Q� ��~T:����l_(�J�>���A9�;$�<��ະae
 *ݩ���`|��W֋rf����"�,�V"��e���d���� �����{b�|pN{d�%2��H�t�38q a���V���⊈�.J �����TQH��r�,�.�B�G�6J��	�`T'���3�,/�ș�e��{P{�1��T3�H��S}�F�/��b� c4�߂�2i�*������_Zp4@C�_J|���/((OXRv��i#~���	"�Ci��۳g�5�c��)5e2Ϩ��y5*-�J��k������V�l$L�QA�r@{�׿��kk #	?É��K�'a�f��k)���Ԑ�*	��Rm�S7�\<�AUU��܊i�V�`(q]uFR��h��5�H
e�����ȓ�kQ0 �ʸ���L,5���I�p@Z��#���@�I��J H�C�y)��3#nQm�}�fn�/��{( ��p^��r$$u�A*(e�  �z���o��3��@����{^E����鳪�()q+M�����cS�"�>�̭,�h�P
��|s߰t�=AJ�:<��#�}�)%� �='f��C�7#/��@�Po�I�P([���$e���$%�0��t� =�bVyqVH��y��'e&��ZՅ=dS�P�MI�Y��Ө-��ߨ�l"X�nTW����s�X�46�0�V[)��w��|��7����H��_u�O��Bb�O�d������P�2��}�4��h�I�%��*1*�g$h]`@���E2)%6�Y��+/�I��@�K����t��H�V�$���ǩ��d�9<fl$;�VJ<�{�'����${�$��p�\$ӡ�쇉?
�Y
E�Bj�+#��v��{c�j��2ɤ�K�h-ģ��l&��A5B���2��:�P,����<����hVˈ���pd��{LE�$��۲�l�e��6��7�#���&��$���H�>���[2�QH*԰�������@ h�

}٫�
B�;��үS��kcG�gP�;lt��X��
̠
�0ނ!  #�Z�.!�w8���%������did��S�:l���= F��TBXA�n�5����������30hT�h�����(���2�c��r���=��/���2�B� �%T�3�2>�9׏P}���/��[����0e���c۱:d�ɤ�KEJ�]Qe]Ds}C#���'��*�M�.Hl��!i�鋬[�5�1+�� BA˸��eDy�>���!��+%��&�utK�qL�U��V�H�SQ4���2�|;�������]�i���,��=-!�HS������J$�h��ֶV9`�dѬ�22��6H����FB���*��XYU� =
�c*4Q:+v78,3��O��փGl�)��d؏TUç�r�~��!�k���=��"�����9u6��d"_u��K��f �,{H��[��dPJ�(�� &aޠ���o{�dn�4)-.��
�Y��Ws�d|���6�r�HJ��ѷt1`1����
i;�.w7ʕ�J���Ǿ&i��^``?h�Ò��p�x$g�q�]9 ���<�*3*�dɼY��|��E���;o�� ׍!�+C�WR�|}��H	�-R�4m��(�b�o�|���d�v��w���VK(�`���A)Dq,��=9��Lp���|�u�\m���)0:���-�lv��o�����0J�C��nA,��(~`xX>۴S�0�d���)5�j�/��ξ�H��8�A�tu�N�*\n7�!Z�
�����7�e'ϓ�s�lf%]ޗ��3�^�o�97�/'���Ő��y@Zpc,1V#���������+�Ε2��.M%,0~hĸ�����f;l!����%�\bU�xvJ��1mt��� �
3o��P�4wt��sda]�-
��J���1��O�V��0�ל.J{��A�#Q[�π�=0h��n���"g̝)sk�I����:�x���oj�-�Hc[�Mr��$H-�ߍ7�hw����@S�Hk��O�%�۠kK�FCk��������D̨��T��m�����F����#�����t��fm[���Æ["��_$��Q�>�[lLi�,n���l��Ma�.��X�f0�����(] �+ʤ��T*K�RRTh��Z'��a�g$�hO���xN8����x"�PQl9���=���N���ʋ�ԛ�h#)���lS��vx`�g[�zCK���C�CxG�0@�ZC"F�Փ�v�M�z}�c-c��'���������Pg�Ήxg	���H}�Z(4�pɄN�ŝ~�u�u�YF
�x�W�Ą��Q58 �1��nq���g+8H�o�ħ��I��������9���DS.q�޹tc���/m_D�Fps������W^iG��<�E��k��L#}�9YhI�E�m�H[h0f�Z��m�)=�^��d	o��}j��U�!�(���&��`L@`8K��>�7C� �Z0�xK�n�ak�׉�2
�#�d#F+��1H+��Vm�1p`�Y
���&� ��-a����=2o����ZF��O�g�F��Uu�7Dʈ����J���6c��p� I���РF��n2�;+��E�u���
��DM(s��%��*����o�۳U�4J��1jv얂��޲�wi5�!ZL@�L0�w�y�e
���F{��=�$������.���s�F�����B���-�!�n�Arcm)F@ ��5����21ʈ(I9Fs*����v�`����R��ڦ�-qZܺ
E�T�Am���]�=����v�A5 &�-�@訊M��@�F�RC���嶥`�]�Hc`� l���q�}N�H��%�梨 y����d��5G����s�v�7��q�]�
ށn���xQ��-���X'�8!���d&ݤˡu�F\\T���`g�`�"���m�Ǩ*�7��0��܉�Ts�TB�d�(6�$��r�U	IB�%�m�G��������%�7�R��%7U�.�x���7ri�6�|9l?ՐO��3n��� D��b 0Q"e��sIm�ц7ZH>b�>a@���B6Q@k���b̝I�k≐��O2���S;�m���?�1��⫉n)HP�vn�k�/�X�º�L%J�i���p�	�'��۫1I"D��ʕ+cnH�3��f�5u��#��X�tH,�o I6ܹ\2�c�{�~W�^-�֭�Y�x�d i'7�<�8ad�1[{���(� �(��G�D�p$�	$#��P�_�B�ސ!Fs���e�5�{2F#���c3.MiG#��a���q��y��)��6#iJ��	��0��&��0��i�h�g.}�z��bef�=�R��^�6�D&����Lx��0���A�|$ ��z������]ɗM4�I0-a��^���K/ى�B.{H�D�ԟ�4�}�v�iY�p��b+��P^�KZ����y���T�x46�L�9�ׯ��)�ݱ[�:~�Ɉ�_���m���d;��}�����=�*��۶m�h^f!��[���r���������:��ۺ�/��w�o��<���:;;�� �f�V�}�RM��K�����gÆ?c�!�K�e�He�s3y72�an@wL>�)\��͹!&������ O?���/d͚5r��ڵk��q�NJ����[�韔$�(H�Q��< Fy@2��d��0��a�$�(H�Q�#' �M��S��iR|q�g���c<*I�s'1I��;��w\e���7㳑Y��    IEND�B`�PK
     t$v[�9�L� L� /   images/b9037746-96b4-41bf-a651-5749520ed4a9.png�PNG

   IHDR  �  �   :�/   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx��ڡ�0 ��
t�]�0�?DT�    ��9� y{����3     ~bp           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��; ���� �uև>ﹻ+k-a��L���:�&Mj�iJ�`���)�G�ȅݳ�P��;i���t:Ljj�v�MpL�@���j��!7�L�&t�v��6�I��6[�c��s��q�HF�w����<3�y�9��8C�=�o�        @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;   �Ut��w�<��`�� CaϞ=��~)3oo{�����   ��B�   pUU�7��] �p�����5|   �U#p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�          �w           A�          @#�          h�;           � p          ��           4��          �F�    pUUUu~ʲ�xV�{>x��7��6_o�c�'�~?!<����y�?I����I��Ǧ?f���u��n�����_�>�?o�Y�����r�~     `��    x�:�N��}�7?�|��Qw9�����`0�o�Zg�o>/�,���o�     	�    FH���������Ϡ6��~;�I!��)���}��׃���>    `�	�    fsx^G���|6�3z��v{��s�sԑ|�����    �Y�     ۨ�gs�~�����{.����霘�8�a>�i     �>w    ��p�8}���ph����i.5�O����ٮ�     �G�    �e��t���?�>���:0�*å��F�t_����ϸ    ww    `d�!j
�c�E�6�ۥ���y�٤������:��    uw    `(� ���7��A{�ׁa��yUG��Ν���B�����F�t�N    �a$p    g0R���o~&\�U�>i.§~p|:7��k<    �Dw    �K��Ӗ�:���m� \���?����[�7��u �>    ���    ���7�����ә�~@3�F�-����z�{
�c�:�O��    ���    �,)`�P�^od�Zۂ���?�Ϟ=�U��������    �\w    �l��^��i���6>�����4�6�o����    6�   ��J�z����vH��ϝ;�1�]l������	    �'�:    #,m��7oc���l��S��"�z�{�����    �O�    # E�i�z
��)bO! ��o�:{��W}�"�͓��ŧ8    ^w    )XO�_�ne�qR�{p�<�/���   �p�   @���1{z \\Y�ٹs�6f�z�����Ƥ�t�(    h�;    �:\�ʞΪ�2 `k���={��3��[��轞��	[�   `�   `�X�B���  ;�b[������i<    �}�    �R����ld�q��{��   `k�   �2���gle�G� ��b������F�v��B    p��    p)`K!{
��=ݧ�  ��OrIs�����Rܞ6���}p�{
��    paw    ��j+{
�����5 ��J?ݥ��y���[�S�n�;    ��;    c%�f�V�t��)p ��O�I_�9u��Ƴ�����{�   �8�   0�R�����c+; �T�7�9}����V��{=    0��    ���	u0d� � }�^��gϞVo{O�{��3=   �a'p   `��+����� ����~�ԩ�g�w    F��   �F�����e  |Ņ��drrR�   �P�   �u�^O���3  �̅6�F�iҽ�   ���   �#ʲ�����iR| ��I�����zꩍg)n���Ȯ���;    ;N�   �UQ��g
�  �Y�k�z�{��y~~�{
�ӴZ�    ���   �-���7"��g�n�� `����S���'�|r�Y��>55���3E�)�   ��$p   �9���== `��z��9}���}�[�S����s    �Rw    .K��^of��v  �O�	=�'��yꩧ6����)t߽{�-�    \�;    �����h���S�  �~�O�uc���OLL���N[�   x6w    γ� ����ar}}}cN�:��lp�{��   �	�   �T��=M��� �v�Ж���[�ӴZ�   ��$p   ���4). ��4�u�O>��lbbb#xO[��999i�;   ���   ������e�O�>��  �A��ۘ/���i�{��>   Mw   �����ofO1{���6L  v�k��i���}jjj#t���ވ�mx   w   �!������g�i�%  ����p�8͗����g�����y�   0|�    Cb0hO#h ����NN�{��>11���޽{c�    �A�   �P�A��3g�~��  _[���<��S�w   �!"p   hA;  l�;   ���   �A;  ��;   @s	�   �����o�����7�Z���]�  �p��}jjj#t�Ͼ�رc���{�d    l;�;   �6i����������W�n���  ͖��s��mL�瞅��?���������WVV�3    ���   `�����]�v�\��������N�<}�  `hM�oX�������������?~��H�dyy��g��   �w   �+433�ڷo�+�<O1{�ڿ�,�]�3A;  ��=�Z�y0�dEQ�e�����Z��?~�s    WD�   p���nj�ZA{���8�O�C  0�n�3�fz�^
�?�I�{��O޿�   pI�    Ϣ(�B�~:h��q^l;;  �5����y���0^?�9w��o����g    \��   `���Lk߾}���������P  �+Պ��y�,�;'''�(��Si�{�������?�   p�ߜ   ��������}!�[㙢����>  �b7ę��j��륟��x�H
�˲����ҩ   `�	�  ��s�رݽ^,�>�M  `'���K���������O��,//�A���    ƈ�   �����,��ׯ][[{U<w��J+  4���M��<��y����x���ޒ����_�    F��   I�v{z׮]7�ey[���x�8  .�=��!�4����?��'���ö�   �J�   ������Z�����R���eY��   FC+����<��*�b5^"��p�O,..>�   � �;   0�fgg�ٻw�ʲ<o��oV��  �X��P|J�+��?������#��ˏe    CJ�   ��G�޸����­���eY>/  o��}oI��yV�g��#UU�<}��o<���g3   �!!p   mff��o߾W�Z����^��C�  p17�i�W����^{f~~��<�O����?~�s   @�	�  ��y׻�����������WU�  p�v��w���^�}EQ�Q|�p��KKK�%^{�   E�   4BQ/!�������׿/>��   �jߖ&��T|�����˲����ҩ   `�	�  �S�+B3��֪��=N�   �Z^�P|;������?����������3   � p   �����k������,o���(��WU�  ��v��w�����.,,��x����///?�   \%w   `[���}�!�o_W���  �&˫�:�y��U���׿��ܿ�':��Z   �M�   ��+����q�?�w��3   ��7�i���n���cUU}tzz�cw�}��3   �-$p   �DQ�!���[���  ��>����3gΜ�����<�O�Z�_>~��_f    ϑ�   �"�N'_]]�9����7�G/�g  �ظ&���{��{����x�P�/..�Y   p�   �%;|��x|wY��=���3!��K��  0�Zqn��*������ӱ��,..~&   �Dw   �Y���鉉�ׄfʲ|c|t]zn[;   �����4EQ|6ޟ��---=��P   %p   �ʱcǮ?w�ܭ!�[����\�  ���)Α��y�(����UUu���}|eee=    p   6=z��^���x�浵��Bhe   ��^��9ۓ��ݢ(>���C7�p�ou:�^   �=�;   ���(n���!��^���̯   p��0N�,�v���B|G����!��  `��Mk   3�v{�����S�o_O�>   �N�>Ρ��zhrr�EQ�L�����?��t�2   `l�l   ���̯	   �\/Ȟ�ݻݮ�   ƌ��  �%j  `��  `���m   !�|�;�~bb��UU�9��'�   `4l���,�_���C�   �C�   C�رcן;w��zS{UU��  u)v���|������(~z���:�N/   ����  �!�n������������6��   ���g_���DQ����/,..~2>�2   `��  `H���^3==��OojS�k3   `�q�ey�(���돤��KKK��   CA�   633�zы^�=eY�H���8{3   �R�8Α�(�O���UU}`ii�g   @c	�  �a:�N���z�ӛ�o/��   �\|C�;���EQ|&��������'   �(w   h����ps<���vgB7f   �vxyUUw�w�^����_^__hee��f   ���  �ZXX��x����;�|S   \-!��K399yOQ�B��ӧO�x*   v��   ��cǎ]����檪~$N��2   `'�qn����޽�xQ���}mm�+++�   p��  �*8v������[SԾ�����h2   ��8������/E�������ϫ   �Vw   �&�N'_]]�9�phmm���ho   ����}�(�?�׿�j�����q   l�;   l��(^�C�n�GC/�   �Q��8w���;�׿���>t����f   ���  ����q��o��j6޾2   FV|�?��V�����qzz��w�}��3   �9�  �z�[ߺwzz��OG��ϐ   �B8σgΜ��(�������w��Ϫ   �lw   ��N'_]]�9�p(��pUU{2   �,�.�۫�z{Q���*�reyy��   p��   p	�=��^�w{��m�n�    .�%q����'�����/�e�����S   ��   p�~^����xy���&�!   �ty�[���%��(N�y���������   ��"p  ��N'_]]�9�p�,�;�ym   ���3S��LQ�����[ZZ��   8O�   ���ܷ�Z�ۻ��!   �>=Ν!�;��+�O���<�T   cN�  ��j���MMM�^U�l���xf    WSUU��3�wﾧ(����_ZZ���Q   cH�  �ؙ��;��y;^�QUյ   �Λ�s(�p�(�����Y>q�ğf   0F�   ������y����۫��[   @s�8Νq~b~~�Sy�����}teee=  �'p  `du:���'�xuY�i[�TU5�   �<�p�������_,�⡲,O,//:  �%p  `�9r�eeY���v,޾$   ~/���󼽰��X�^)��KKK�2   !w   F����5{��-mk������B   0���:��	!��(��y��,..~2}�  ���  0Ԋ�xE<�y{UU7��k   ���83eY�E�?����~������   ���  ��s����eyG�|G�o�    ��8�i�Z��(����'N|*��  �!#p  `h�����]����=    �M���4EQ�I<�Vw   ���  �F{�[ߺwzz����Ҷ�o�    �Tߔ}e����y�������Vw   L�  @#����e���f    \���}�,˙���?!�?���   4��  �Ƙ���fϞ=��e�!�    �R!����=eY��  @#	�  �q�~yY�?/�UU� ��   ��lu  ���   �w���מ={�-UU��,���    �[��EQ��?s�ĉ��   `�  ���9�~���3g��x��>   �)v���4EQ��x>P������3   �J�   l�N��?���.��h��C|2    ���'��VŇʲ<�����   ���  �ms���{��l�۝��/�    6{��<o/,,<V�彽^�C+++�   l�;   [nnn�@�M�^�w(���    zUU!|`rr򧋢x0>Z>q�ğf   ���   l����k���(�p,޾2   `T���8?1??��x޻��t2�U   ϑ�  ���ȑ#/���o��?��   �q�����������OMM��=���   ���  ����t&VWW�B�������B   ��
!�,�Y[[���(~�,˥���Og   p��   \�v�}����l��=Bxi    ϴ'�;�<����ceY޻��v:�^   �@�  ��477�-y���˷WU5�   ��PUՁ����,,,����ݷ���x   �B�  �u:�|uu���H�5�    \����.wMNN�Ӣ(~�,˻���?�  ��  x�v�}����l��}W�2    ������PQ����۷�#�N��  ���   l(����mUU]�   ������[���/,,�l�^<q��   cO�  0�:�N��O��,ˣ��qB    W�_���x�Y�C!�s�}���  ��%p  C�~^UUo�v����f    ����s���CEQ<B8�o߾�t:�^  �X�  �����o
!��,��x{m    �sKUU�t������p�,˟_ZZ:�  0�   c`~~�U!�#��MqZ    4�ߨ���¿*�������?~�s   #M�  0�fffZ/|�_/2��]    ���9�������x��O�8�{   #I�  0b>����~,�?��/�    `4�qnM����XY���߿���N��  02�   #bnn�<��eY�3�^�   �����@��n���(V����_YY�R  ���  ����y����g��    /7�y����OE�����{�?��  ��%|   B�N'_]����y�\�}��V�� �� A \DI�����[d'�g�q<�D�����u�)іDі�6%K�%��zی���'9���9�I�dNF�iS�.X�������ߍ�܉��~�s~��nU�����n����w&Iroq��    ����555��c������   �;  �<��ۻ2˲_�M�dk     �V-�]q�4�/I��Vgg�7����   �� �  0|���8==ݓe�]��     �����GFFF�m4��Zm�<0   hi�   -쮻�uzz�155�U�    ൺ9��'&&~��h��j_y��N   Z��;  @���oO�����w�I     ިy�zbb��4}xɒ%���C
   �w  ����W~g�$��?    ���������z�4��I������#  �� �  0�z{{�NOO����ȽI��9     ��V��y�ߞ��-�/��   ��p  �#���+�<�@�eO�ds     ��_K��ߥi�h��lذ����M   f��;  �,����^�V�β����     ����$��GFF���C����/}�R   `��  ̒���U��O۟>�   @+ۑ����������_)�;w�<   �q   3�����dYvw���b*    �/:�$�����i�����o�ڵ�H   `��  ̐z���$I�ɲ�]    ��VsW�Z�N��_���   \s�   �P___exx��I��jq��    XHڊy_1?���Ȳ�o�Ν�#   p��  \]]]�%K������{�$yk     �J1�T*�L������   x��  ހ��ޥ���?�$ɧ��[    ��$ż+N���5��/}�8�   ���;  ��p�w^�lٲ;�,�x�$�    ����$I�]������GFF~oϞ=�  ��D�  �5����P�V?Rl�y��
  �{Y�����}|jj�E�����r�T*�x�����Z-$I�� 0o}O�^��6l��^��xO�{�w�   �*�   ������,  ���x�(�k�ǰx��y&&&ʿ�����c͐y�o�4�Ϳ�:������7�v��:�dɒ2T�`}s��\���}���v���|����5N|,>���iN� �k����?*އ�z����ŋ����}m,   ��  ^F�^ߚ$�G�퇊�  �H�7��q�z���TP�ٌ�답��ʚa���϶f���||,��i7�����|�� > �"pc����˗ߛ���{��ݻw_   �(W�  ^D��ۊ%6�w�  ���A���7���f@��m�ǶsfN3\�B��xo������}�y �yhc1��e~��h%I������  �p  �J��ؑ��'����� ZB���f||�%������+^�� uؽ���ⴷ�k� Z������I��`�����   @ɕ\  �Boo�[�,�D��� �� ̰<������+k��
��������J%,]���x�A���x3��� fPg�ONNޝ���,˾�s��3  `��   ����U�ՏgY���  ^�f�6��GGG�5�֯�7��5�\������8�Fl|o�_l:::�0|��sE  x�VsO�RI�->?44t<   ,R�  ������=Y��j�}w1I  x	1�/_.C�q�������r�&�܁�cjj��K�.����6�f�=�ߗ-[��|\�� �`E1w%I��4M�X�000p4   ,2�  ������'�,�� X��ns��l\�zbx]px%�/qΟ?����mmm/�7[��� ����U|��4Mw'I�EAw  `1p  �����T*���] X������gh��X�̦x���rA�j�Z6�7�q�<n���`QXV�G�<��i���3�}�v�:   8w  `A�����,�b����$ X0���.]*'Fc`�y��ׁ�(�@�弔Z��/_~��=ߛ�q�q�� D[1]�j��t/^�]�;  ��	�  ROO�wW*�OfY&� �T�7��WO|����XMNN��gϾ��W����{�f~Ŋa�_�<T��<��i�~�x?з{��c  `�q�  XP��w�y���� Z^lW�A��/� ����6v ^�Wj�okk�|o��c���� -mi1]�Z���4����燆��  �B�  X����V�V-�s�v h1�i����W��q���SSS��711QΙ3g��s1��l{���]�; �����U�v0݋���=��C'  �<�
$  0��i����b~��J  f]lb���f{����gY �?�y�y>1K�.-��/6���e 0ʠ��Ԕ�;  � �  �Roo�[�,�D�}O1�  ̨f�=ׯ��}|<>��0>>^ΩS�^�x���v��뮴������ߙ��`�e_عs�   0��  �J�^K�$�fY&� 3 ������A����_Yc�}jj* �K����ĉ���f����2��r��2���V�*��kjE1�����;  0	�  �BOO�M�J�/hl�kbbb��7ٛ!vm� ̄��f�����/x����J�=���5N{{{  ސfн��h�V�z������   ��� �����{C�e+��X�Z? x�&''��z��=N3` � ���ԩS�\mɒ%W�� |\c�; �����I�|$M�/���}�   -J�  hIi��+��eYvW�v �e����s�ΕA��٧�� �G�5��ٳ�\-ߛ-�W�;:|t�W�Y����$����?   Z��;  �R����:::����bV �b���{sb�- ,������\-�c�}ժUW��q��� �7�y�`1w7�ϝ8q�w���3   Z��;  �>�я.m�{�Y `�˲,����̙3�ڜ<� �B1�_3�\�V��A�իW_	��Y�&T*�  �ܶ���W7l��F��遁�U<�'  0�� �9����v���;������M ��u�J{��=٧���599N�:UNS��X���ǉ��8K�. ��%�����cI�|f```O   �C�  �����[2<<�����O�7 Xb�z��=��Ϟ=[�̎�� `��;�4\v����c������E��<���$I>900�  �p  fU___��ɓ?;22��$I� `������C�q���Z��u�T�{��Y�jU|��%�f`���<���z�����W����{   �E��  �&Mӟ>y��g�<[ �djj���6��/�A���!w `~�����]m�ҥeؽ���v����� `�H��ǋ���4���J�����  �Y �  ̸����T*_(�?��y ��,6�6�͆�.�q �������Ǐ��$����3Y��t����$�=�  �p  fL�^K�$�^lo 0MLL�A�b?}�t��a6 ��b��+V�����V� �g*�ܞ�y�mzz�S�v�   3@�  ������$I>Yl?XL5 �<055U6��{s.]�  ވ�/�s���+�-_��J�=���u�_�0/�[�tU����i:8::�?���   p�R  \3i��+����b� ��,�ʠY3��� �i�Gtq�9R'I���2�jժ�f͚r*�J ����{:::�L����׬�����  �&� �7���kY�V�-���* @�+C�N�*'� @+��<�?�������1����=6�@�Y_��Y��4��uvv�N__�_�  o��;  �uuu����>Pl��<� ��0{lc�z&'' �|255u��yMeн����1 -`[��_=y�do�Ѹo```O   x�\�  ^���h�;˲�����  s$��^�p!�;w�J ���S ��dtt49r��(I�p�uוA������Y��q �����˿���X�T�x$   �F�  �k�����y��_�_��9 �-6�^f?}�t���  �Q��_�q��?����1�nݺrb�]�; �-I�x���4�W�j�W��<   ^%W�  �W����{�,�b13 �,�f���1� ���?l�w��-���{�e˖ ��!����鿛���b�o׮]�  ��  /���{K�Z��,�>XV ̐\���'O���q  �~W���߿�|l�ҥe��ڵk�56��K 3�VLZ�V�H�t`tt�7~��  �%�  /�^���T*�����aG �k,��7��q={��vv �YDx�ȑr�Z�V�ݛ�k֬	ժ߸p�-/枎���6��N�8�{��   �A�  x����Z[[��<���� �����022r%�~Ⴒ6 �V099N�8QN��W�^}%�'���5�%��nذ�ÍF�o```O   ���;  pEoo�gY�`��) ��O�:U���z���  @�w�9s�L9�<�L�����Æʰ{ggg��p�7 ް��9��^��a�Z�x��  � �  �2��}Y�}��	 �:]�t�lg�a���y���  �����߿��H��k%I�X��H���?==��]�v  ��&�  �X��ۊ�3Y���X�  �Rl��p�Bf�����>::  X^,���k׮7n˖- �T���Z��+MӯLNN~~����  �(	� �"t��w�����x��H1K ��h?w�\8y��@{�Z   ���8�*��x��-A��j����+�ʃ����  XT� `��;ڗ/_�቉�{��U ^F�� ���p��>55  �������+Bgggz߰aChoo �2�s�ew�i�����  �EC�  �z��SI�<Xlo
 �"b )���0��c����X  �k��ŋ�8p�<��1�~��r��� ��7��4��b�{pp�[  X�� `�k4ߛeٗ�$��  W'O�����  0�{������$IX�jՕ�{lz�T* ������4M�Ւ%K>��C
  ��%�  Tww��j��ky��B�$� LMM���@�ٳg  ̵<����q�����jX�n]v���~�!x ��bp����;�4�/^?>;44t1   ��;  ,0]]]�j�Zo���b� ,Z���eH�ԩSe�=N @+��c�2��ݻ7,Y�$�]��J�}����EmY1�$I��F�q_gg�����e  X0� `�H�ƻ�<�b�� Xt�͗�0Plk�2�� 0��;]x_�lYt���8K�. ,J[�<����ȇz{{�����	  �� �  @���_,_���� ����X8q�ĕ����D  ����������D�V�
7n,'6�W*� ���Y���4M��$�]�  0�	� �<V�׷&I�����$�/6��9s&?~����v  X�Ν;Wξ}�B�Z�֭+��7m���� ���<�"M�]�J�S����  0/	� �<�я~t������<��8l ,h�.]*��###�:99  ��hzz��ݍ����/_6l�P�c���%�X�ڊ�+˲�4�Ϟ8qb`Ϟ=�  �W\� �y���o�nܸ񃣣��� ���T8}�t��~�رp���   �v�Ǣ���/�R�����2�C�W� ,X�y�?X�����444��  0o� �<����}Y�}%��� ,(Ź=�;w�JK�ɓ'Cq�  ���c_�����^ݯ���r��j��/'I��4�f��500�?   -O�  Z\ww��j���,��[&�a||<�8q������  ���*'I��nݺ�q��rV�Z XPޕ����iKd>;44t1   -K�  ZT___�ɓ'{�<�Lqx] `�;�|8~�x9�O�.�� ��ߛ�;)ŉ��K�.-���=�K��Z`�(�$I�[��ehh��.�  @r%  ZP�^�������� ��5==N�:Uڏ=FGG  �������J%tvv�A�-[����� ���%I�����������  ��� @i4o����b�� 楱��022�;N�8���  0eY����y���ʕ+�f�8k׮I� ��+���J������?�k׮�   �w  h===k*�J_����}:��R��ùs��@{lj?{�l   ���ϗ�o߾���v%�aÆP�� �J���U�՟J������?���7  �9%8  s����2<<��$I�Xn �����ɓe���ѣa||<   ����D8t�P9�J%�Y���o޼9�X�" 0o�.�����4���c   挀;  ̑����>22�P�$� hy/^,�qb�=6�  4eYN�:U�޽{�ʕ+æM���{�'I hy��y��4�fq^��Ν;�  ��p �Y���Ʃ������ -+�Ϝ9�;V��ǀ;  ��u���r�zꩰt��2���ׯ__�����U��<M�/MNN~~��ݗ  0k� `�tuu�����SSS�-ݣ��P��ӧÑ#G�   o���x8p�@9�j���p�e�}�_����b>Y��>P��ehh�  ���  �,h4?��y1o �����022R�c[���d   �)�3����ˉM�k֬)��cཽ�= �r�$I��4M�(�ۍ����  0�� `uwwo�V�����}��111N�8Q��:55   f[�e�ԩS�|����V�
�_}v��� -��y��4Mw���~���  �!�  3�������V���3šo#Z��˗�ѣG�@�ɓ'� 	  @���<�={��'�|2�\����Y�n] �%Ԋ�����g����}#   ל�;  \c�z�I��y�� ��:�|8~�x9�  `���g��۷/,[�,lܸ���5I� ���R������žwpppo   �w  �F����T����� �Dl<�A�cǎ�m�  `���m���_�ҥKæM�-[Bggg�T*�9�b�$Mӝ����|��/  �p �7�������V���3��u�YC�O�G�	����  `���y8PN�V�v߰a��;�ܨsWGGǻ����CCC�  �"�  o@�^G�$y��5 0k��  B����*G�`�mN���i��Q�{�  �up �ס��{K�Z�|�}_ `V�  �4aw���b�$Mӝ����|��/  �5p �נ���V��b��b� f�P;  �k'�0�j������3�z�#CCC�:   ���;  �J�z��Jeg��o ̘�C�q���   ���;��ښ$��7�?(���  ��� ������T*}Ŷ��o� f@��<y�li?v옦v  ��a�͛7��q�Ɛ$I `f�y��b��F���������.~ ��p �������%I�b�> pM	�  ̝v?x�`9mmme�}�֭aݺu�� 3�#��OgY�����z�  �E	� ��H��MŲ�� \S�ϟ�?�|�j  �{���崷��-[���� \[I�ܚe��������Ʈ]��  ��  p����emmm�����- pM�P��#Gʶ��/   Z���Xx��g�Y�lY��¶m�+ ����j�o6���������,   %w  �s�z���$�J��� o���hj?z�h8u�T   `~�|�rطo_9+W��7o7�xcX�|y ��X����'O�|_���x$   �  ��ݽ�Z�>Plo �!��'N��
���  �P�;s�yꩧ�ڵk˰�֭[�ҥK oL���X��������'~��  1w  ����%'O�L�<�Lqx] �u���Ǐ/C�1�^�W   S��������vX�~}��iӦ�d���ހx�������z�ޡ��o  X�\a  `Qj4mdddg��� �k�eYf����p{�  ��İ{�{W�n�!���aÆ�$I �u�\�C���黋}�����   ���;  �JWWתZ�v_��� x�bp�����ȑ#����a||<   @455U�:N[[[زeKv_�n] �u��b~,M�������g�  ,�  ,�z���$,�[ ���������P���X   ��311���_�ʕ+ˠ��7���� �ɲb�߰a�߯��]CCC�=  �" � ����յ�V�}�ؾ; ��0Blj��{�N�
   �z�M�ݻ7<���a�ڵe�=Β%��x�r�$�o��Cy�������   ��  ,dI���P��_,�+ /+˲0<<:�=��g   �k!~ƌ?����c��믿�lu߸qcH�$ ��b����w��z�����  `�p `Aj4ߕe��<�  �Ξ=[��>���   ̤����aq���Ö-[¶m�ªU� �h{�$�1M�o���]�v	  ��� ���q��+V��D���&I� xQccce�������Ew4  `n�ϧ�>�l9+W�[�n-��K�. ��wU��o7���������,  �!� ������W�<s �/�yǏ/��'N�(o   �����a�޽����ׯ7�xcؼys�V���:������^������   w  潞��5�J��b��b� �1�>22���p���055   ���ϲ���崵����۷o/����$��b��4M�\�T>���?  `p `^k4��y>Pl7 ��p�Bj�m��   棉����ϖ�f͚�m۶p�7�Z� x�xb�gzz���6��  `�p `^���޾dɒ��y��R�e�رc���e�   ,$gΜ)�����¦M��V��^ \-I�[���Ʈbo��   �;  �M�h4>������. Ξ=[��cc���T   ��,���ȑ#�ttt��[��;v�e˖ J�<����3�F�>00�o  �#�  ��z��$I~;�� ����p�����p�ܹ    ����hطo_x������Í7�6o���j X��<�T,�&M�=����ݻw�  0� ����������r�� �<�Cq>,��cK���t    ��g����rj�Z���V�U�V ��Ź�����}#  @�p �����|������� ����X8t�P8p�@�t�R    ^Z��Y��Y�իW��[����mmm`ې$�����˲�ghh��   -J� ��t�w��X��y��[��	Xt�,ǎ+C�=6�   ��ٳg�y�����͛����Cggg X��<g�$�5�O������,  @�p �����J��w�<K Xd.\�P��<x0���   ������?�|9+V�۶m+��Z݁EjU���l���088�/  @p �etuu-��j�Vl?VL% ,SSS��1�~�̙    ̜�/��{��'�|2lٲ%�ر#�]�6 ,6I��p�<���iϞ=�  Z��;  -��h��<ϿZl��E"���߿��ǐ;   0{b�{��Z�뮻.�x�Z݁Ũ���ׯ_�s��������   sL� �9���|d�����<�Pq��.˲p�رp���0<<   ���[ݟx≰iӦ2�aÆ �X$I�W�,��4M�\�T>���?  `�� 0g�4����ɝ�vc X����cS{�OLL   ����9r��f���;B�V �@<��S��v��w�q  �9 � ��k��ۮ ��ik  ���;[�o���nݺ �|W1������ 0� �U===��]l7�jll,:t(<��satt4    ��խ�W�۷o[�nK���X��I.�����h�100�H  �Y�7  �Bk;���y�?^���8q�<   ��gφG}�lv���M7�V�\ �������� 0�� �qi���?om� �f[������˗   ��MNN����V�[n���'I ���=��w6�hs `�	� 0c�����p��~��Qm�   ���V�Gy$<��ca۶m��o���`����mŢ� �'� ����,DSSSe�=��]�x1    4����}���g�y�ls�馛5k��� �'� �5��X�b����,C�    /%˲p�СrV�^�o�n���P�V�B�� ��$� �5��XH�<###��g�Ǐ    ��ٳgã�>���[��o�喰lٲ �@hs `F� ��im���~������ҥK   �����,D�7�_�>�|����� �6w  �5w  ސ���wNMM�v�� 汋/�_2<x��   \k�q����X�"l۶-�ر#�j� 0ϕm�Y��doo������4  ��$� ����յ�V�}����y��y(˲p���A��ɓ   `����ݻ7<��Sa�֭�[n)C� ��wgY���4�����v��=  �5p �5���?�$�׋�-`���M�1�~���    0W�����_Ά��7����� 0���R�S���FOO�?ܹs�S  ^w  ^�;}���}����T�<s���p���p�С0==    Z���p9��}ǎ�T�.����W*�?I���ׯ_�ž��,  �� � ������ݕJ��� �H���ȑ#e[��ӧ   @��x�bx��¾}������V��K��y��������^��944�|  �W � �����[222�����b��<199<X�/_�    ������SO���~:lڴ)�r�-a�ڵ`�I��ǋ�ۍF�c�  �w  ^Roo�[GFF�^l�7 ��.]
���/C�    �]�e���^���oٲ%T*� 0�������z���_8  �E� �b�F��,�(���<p��ٲ�����嗾    Q���#��'�x"l߾=�ر#�j� 0_$I�y�?Z�׻����u  �� � �twwo�V��(�� Z\q�
'N�(o�}���    �XĻ��ݻ��.�u�ֲ�}Ŋ`�X�$��i�������p� �+� ��^��?I��b{] haSSSa������/_    �U�:Ɂ¦M���7�:;;�<q���������Ν;�   @p  ������xK� ��b�=~agrr2    ��;�=z��իW���[�l	�J% ���sտO�thrr��w��j ��	� ,r�F�'�<��^ Z�ٳgó�>>�,    ��x-�G	O<�D�馛;B�Z -,)&��j?����ޝ;w��  ��%� �H�}����y~W hA�u�ĉa߾}�ԩS   ���ҥK��O=�Tؾ}{��t�� ���\�T�[����'N|fϞ=� �EG� `���������$ɭ��LMM���g�y&\��N�    o���DY"�w�7�[o�5,_�< ��%y�z����^��ohh�  ��"� �����-��,�>�$I- �������sϕ�t   �ښ�����7n��v[X�vm hEI��@���F�񱁁�� �EC� `�h4;FFF�Ql� ZH�Uvl�_��/Y   �Yy���Ǐ��nݺp��7�͛7�0i h1+�s�W�4��b������  ��; �"P��ߟ��`�] ZĹs��3�<>�,    ̾S�N��|��p�M7�S�T@���bޞ�靃���!  ��	� ,`����,��b���E�/L���W6�   ��]�{����O��۷���mmm��l,�i������ݻw�  X�� �z��Y���b�9 ̱x��G�����g�    Z���Xx��'�;�Š�������@�H���jo���}o��  w �����������u�`�dY�9�z�p�    ��055U�ܟ{�p�7��n�-�X�" ���fY�G�F�s�������e �C� `�������ؾ9 ̡���[Z��/    �X`p�С���χ�7�7���a͚5���<����ȏ���844�|  `Ap X�F�qW��Y����a�����g�}6LNN    �<������ٰaCx�[�֮] Z�;�$y�^����  ��'� 0�uwwo�T*_���'��p�B����b�    ���p9�����n+� slU�$�4Mӟ��>44t1  0o	� �c�z�'�$�z��> ́���_	��/    ��'O��jժp뭷�n�!$I ��������i�����?  �K�  ��w�Ѿ|��/��b|[ ̺s�΅��z*9r$    ���kE�<�Hx�'ʠ��m�B�R	 s�b�[���\gg�}}}}n;
 0�� �3�z�-I���b�=`��:u*�۷/?~<    ��.]�}������7�v����j ��<�?=22��F������� �yC� `����O�dg�] f�`;    ���˗�c�=V^O�!�[n�%�j� 0~,��G�4�spp� �yA� `�����j�[l�N �E1���O�3g�    x-����kK�=�\�馛�V���� 0�����4����ɻw��}9  ��� Z\����<ϿQl��YP�s'�   �&&&&�kM�<�Lضm[xӛ�����,J���jo����;w���  @�p hQ}}}KN�<��<�?UV�����G��_6�?>    ��455�}��p��AAw`���R��Q�������W��<  �r� ZPww������+�? fX�>|��_�x1    �L�Π�m���.] fI{���i��b�����S ��"� �b�����$,�+�ʲ,9r$<���ҥK    f�Fw`��t1������;w���  -C� �E�}���ۻ�������O?�t    0��A���۷��iK�R�Oi�~qxx�W���3  �s�  -����������ؾ- ̐��۰�|�I�v    ZN,f�A�X�����7���R�=7n�����ߵkב  ��p �c�z��Y��,���h۟z�0::    ����Y1��iŠ�m��:::�L����W��G{zz�عs�  挀; ����]�e�W��� 3 ��p�����O�K�.    �O���p�e�������T*�>M��������o"  0�� �@����,��y��9 \c1��ll�|�r    ��,�:T�9�F�7��Ma�27EfLR�]###?���������  �*w �ٕ4���<��b� �!��    ,d�F���۷������`��ª?N���y  `�� ̒���ζ����y�� p�`�ѣG��?.^��'{w�y߇�7 �]�D�Dʢ�/E�%G�#[��-��8��8U�g�x�[��	zN{������$���M�Į�8v�4%Y�HQ����	q@��EX��Ne7q-[�>�s�������,x��;�    �Y����S�FwAw`M.����r���뻯��ͱ�  C@� `�Y�����$�� �B�   �~�����s�̉���ǘ1O�GkkkW���577�  ��; � jjj��������?ר ��   ����}��šC�JA�Dmmm \aK�$y*�������O  �F� `�����uuu�Yq�� �~l߳gO�?>    ���A�#G�������t���I�<���������mmm� �+N� `d��_�����ű. ���{zz    xi����w��R�=ms�={v�����+���K������� �%� peer�ܿ*^�Cq�
�����ӱ{�����
    ��|�rl߾=���_jsO[�݁+ha�$����o777:  �b� ����ƺ$I�kq�B �F��ݱk׮���    �ջt�R�ر#<Xjt�5k��;p��K���\.�r���k>��O]  ^3w �+ ���l�P���8# ^����Ǟ={�رc    \9/^�m۶���ϟ7�|sd2� �>z�ҥU��w���|�3; ��D� ������'I��sm �J.\��{�F{{{?S    �^\t?t�P,Y�$n�� ��5jS>�olnn��  �Up x�r�ܵI��yq�# ^�^x!8PZ�B!    �����O>�d\s�5Q__ӦM��h|�$������뻯���b  ��	� �
�lvU��L&ss �
}}}?����    0<�������ӧ�-��W_}u �F���]��fW���  ^w �W&���?�$���1�
�a����}���B�    @y�����Θ1cF)�>q�� xn�d2�����jnn�|  �	� �L�����&I�+�
?;�ȑ#�gϞx�    (?�>ޱc�����q��7ǢE�bܸq�*]U�\��\.wO]]]cSSSo  �S	� ��\nE�P�bq� �@�@,}�k׮�p�B     �/��;|�p���ǜ9sb�1z���5tuu�\�f�y�C �O�� ��f����S�56 ^�'N��ݻ���'    ���������������ٳ���& ^�$IV??6g��{[[[�  �$w ����f'e2�?.�
�W���;v��]]]    T�^x!�o����7��L& ^���ώ��r�u}}}�hkk�  ��  ?F.�[��d�*I�� x�.^�{�쉣G�    P}�=�m۶šC�bѢE1s�� x��_�||̘1˲��Z[[O  ���; ����r�-^�K�$S�e�������ڛ
�B     խ��'6m�S�N�[n�%�M� �D�$wg2�����Z[[�  ~H� �EMMM�;;;�}q�W� ~����R�=���9E    F�3g��c�=3f�(�'M� ���L&�1���?---�  �� 566�uvv�Eq�� �)�$��Ǐ�Ν;KG    #[�_x��ɘ5kV,Z�(ƍ /S���d>�_V����O}�S `�p F�l6��$I�Po������l?w�\     �@�P�ÇG{{{̛7/,X�F�
��#I�_�tiycc��׭[�;  F0w `D���I�4Wm ���ݥ`{WWW     �����ػwo|��ߏ���7��L& ^�E�B��|>�ϛ���  #��; 0"e��I�˟$I�� �	.^����#G���)    �r\�t)�m�V�[\�tiL�6- ^���$�|.�{c__�'���� `�p F�5k�,����R�$��z{{c���q������     ��ٳg����ӧ���'O��"=���G�^�������� 0�� #J>���$I>W\S��H��i��{��^�(a    �+���#6l��f͊E�Ÿq��'�d2o���ݖ��?��ܼ>  Fw `Dhhh�3f��%I�6 ^�ɓ'c���q�     ��҂�ÇG{{{̙3'.\�G�n ?��$I�����UKK�� 0�K �^CCô����'IrO ���;v숮��     l����틣G����o��洩9 ^Bmq=����?~�o~�S��� T5w ���r��˗�kV ��˗/�޽{�ȑ#�$I     �t�r۶mq�С����뮻. ~�]�tiɚ5k���#�
 �*%� T�\.���及k| �#����J��     �SOOO<��q����-���'O��pkMM��|>����� �*$� T����ѝ����8> ?�رc�s�θx�b     ���'OFGGG̚5+/^cǎ�cj�$���r�_WW�o���
 PE������gtvv~�8�L �#��ݱcǎ8}�t     ��B����{.,X��͋��� ���z���sICC�G���� @�p �F>�C����! ^t�ҥؽ{w=z4     *E___�ڵ+����ǭ���]w] �ﮭ�}*�;���uO  Tw �*����$I��1P400�������f    �J�����O<ӧO��K���ɓ�G,�d2O�r�����  �p� @Ekll[(��$�� xѱc�b�Νq���     ��~���3gN,^�8jkk�����*���~]]ݿijj* @�p *�}��7�P(�Uq�3 ������g�-]    �M�$q���hoo���ܹs#����������x��_{��� @p *Rcc�
������xiS��;����    P�z{{K{�G��[o�5�M� ?�$ɻ���r���ZZZv @�p *N>�o(
���ٛ0��ڊ����E     �$�Ν��{,����R�}�ĉ��d2�'���o���~)  *��; P1���q'NlK���x'O���۷ǅ    `$K�KO�:s�̉ŋGm�� �dR&��B>���ӦMk** @p *B>���$ɗ���h�ϟ/�;::    ��%I�҉�ǎ�%K��M7ݔ680�e���ogg�ʆ������� �2'� ��\.�"I��Ǜ����c����o߾(�     �8�/_�g�y&:˖-��S�@�;kkk�Z�f�{y�� @p �Z6��p���5>����=v��Yz0    �Ow���ظqc�ɽ��>Ǝ�����������[��[ P�����z��QӧO���� F����������    �+w���8q�D,Z�(�Ν�L&�mj�P�f.���---�  eH� (;������-��`D��퍽{����M�$     x����bǎ����e���k�`DU\���rKǌ�[=�Х  (#� @Y���?>``ோ� F�B�����c��ݥ�;     Wιs���G��3g�ҥKc����h����;�����mmm' �L� e#�Ͽc``�ǫq�����g�����     `�;v,N�:��͋�FMMM #�����>�����u��m
 �2 � ��|>�$P��s���صkW�h\     �F�ݻ7�{��[��`ĚQ(�f�����~.  ���; 0����q�&M��$I~=��P(����c߾}�)     ��>�x≸�����>Ə��46����\.�3uuu���&o �a#� ���o�Q���$ɪ F����x��g���'     ~i���'b����p�¨�q�.�P����֬Y��Gy�;  ���; 0,���]�L����y�0�\�|9v��G�     ����@�ݻ7���cٲeq�u�������'׬Y�Gy�{ 0���!���>T�|���q	#D�$q�ȑR����/     (_.\�'�x"f̘K�.�	&0�,�����b��� `	� C)���7I��`�8{�ll۶-���b	    PI�?�N���������&�������\�߶���^  w `H|���x�ҥ?O��}�iS��={�СC�w     *���@�ݻ7�{�ۢ��.�eTq}2������˷��9� t� �����f^�|���qe #±c�b���Q|�     ���矏�<n�馨����c�0�4�=zΚ5k>��#�8� T� ��Z�f��kjj��$��T��ǳ�>    @�9z�h�8q"-Zs�΍L&��P|��|qm����nnn�  �D� 4�|��I����8>���Q�o߾�*
    @����;v������n�ɓ'0b�K��\.������ 0�������$��s U��ɓ����/     #��ӧcÆ1{��X�dI�-�#�5���|>�577� �+̝ pE}���x���?K���j��zl߾=�;     �L驞,�/[�,f̘��0:I�?��r�}}}�����  �B��+&��ϸt��W���T��aŁb�޽100     ���<��S�������Ǐ`Dh������|��>  W��; pE466./
i��uT��g�ƶmۢ��;     �G?~<N�:��Ϗ�FMMM Uﭽ���֬Y��Gy�{ �	� �Y>�_](>W'P�Ҧ���}����$I     �K���rv_�|yL�:5���d�������� �� �E&���N�$���T��'OƳ�>/^     x�zzz��G�Y�fE}}}���Pզ&I��\.w_KK�g �Up ^����1���R?@U�|�r�ڵ+�=     �j���9r�T����_���P��_��i.�[VWW�����  ���; ���]�vjWWח���T����ؾ}{���     �Vi���O?]����b	T��wvv�lhh����6� ���; ��466�����zq\@չp�Blݺ5:;;     ��S�Nŷ���X�hQ̟??2�L U�����7�������?}*  ^&w �e�f�w
��Q��*�����={�D�}     0Xb׮]q�ĉX�|yL�<9��ug���l�ݭ��� �ep ^�|>��$I>W�PUN�>۶m����     ��r�̙X�~}��}���QSS@U�1��<���>���� �S� ?M&���n�$���T����ؽ{w:t���     C-ݟ޷o_;v���^W� a�RW�W�����E �� /���q�����$I�kT��'O�Z�/]�     0�.\��?�x�t�M�t��3fL Ugt&�i��r����655 ��p ~��k�N����J&��� �FhO��i�     ��ѣG�ԩSq�m�Ō3�J���|]CCï���] �!� ������޿)����]�vE___     @�z�⩧��믿�t?~| U�}����mll|��u� �D� �'����$��qZ U!=�u�֭���     P)��H���oǢE�b�ܹ��d�*�
�'_�o �	� ?����Y�$m�qL ��~��ƞ={���?     �Ҥ���ر#�?˗/����*��2�P(|'�������  ���r������T_@H[۟y����
     �t�O�.��ϟ??/^555T��I�|=_�����  F<w ᚚ�Fwvv�ǆ *^�P�C���ݻc``      �Z�'��۷/N�<+W�����:��1��$��-niiy���$ �K� F�l6;�����L�T����Rk{www     @�J��7n���������\���ljj� `Dp��������Lfy -mm?p�@�ٳ�4    @�K����bŊ��k���������> ��#� #P.���x���)�����lٲ%Ξ��    �ȓ�?���ܡ������������O��G Q�`�����$I���8%��U|������    0�is��u���������Z�n��  Fw A���'I���qL �̙3��3�����     �_�6��7��7����1z�XT�$In(�G������� ���/y !�7��o�*�� *���@�ݻ��ܞ6�     �T�~������(��O�6-��7�����|>�knnn ��	�@�[�z��������}T����Rk��     ������<�Ν�/���ot�$���洴���⿵A@��; T�l6;����/�7��
�"
�سg��v     x��}�ĉ'b���QWW@�{0��]����[mmm} T%w �R7���|-I��T����زeK�?>     �W�m�gώ��zm�P��Ymm��okk; @��; T����%�B�o�$�@�I[����[jmOg     �;|�p�:u*V�X��*�����n����lnn> @Up�*����,
S�PqzzzJ��gϞ     �ʺx�6w�˒$ٜ�����ܼ# ���t �"���o���8����M��={�hm    �A���wtt��ܧM�lF�$���{Z[[ �*�@�(ް�[�q��������ӧO     04�����}Μ9�6���� *�5�L�[�l��Z[[� @���*���,^>@�Ibv�����     �$I�������+W�����:��46���e�����3 T4w �`�W�UWW�\���\�x������     ����鉍7Ƽy�bɒ%��d�8��$y$�������� T,w �P���c���T��     P~
�B�۷�m�W]uU ��\.7��������9 �@� P�֬Ys����W3�̛�/��B<��3q���      �Swww�_�>/^�������7:;;�]�v�z�K Tw �0�|~F�$�(��P1�;۶m����      �[��k׮8q�D�~��1q�� *�{z{{7444�b[[[W  C� *Hcc�B����o
�"���[�n-m�     ��̙3�6��K���7�@Ź������������� P��B�Y����B�k�qZ �ԩS�e˖R�     �L����2��Ǐ����c���T��Of��w���n ��	�@��r�-^����A([z���      �CZl��o;n�喘={v �#I�2�̆��{KKˣ �5w (s�l�_/-�5*�����O?�t<���     T����ضm[tuu�m�����T������쯶��~9 ��%� e,��=X�|2���$I��=mn/
     T��{�r_�|y\��T�q�L��|>���� @Yp����r��x��({/^�-[��6�    ���������1w�ܨ������ *¨$I�(���iii��  ʎ�; �����ѝ���/�#��w�رغuk�HR     `�IOx����o�=�L�@�x0��M���{����� PF���444L����bq|g e-�?�����     ��������wb���1���d2T�Ǝ��k>��֦�
 ʄ�; ��x�꾾���7P���-[�ĥK�      U(b׮]��+W��q��P�2�̯���^�v��<��C @p�2��f�����fq\@�J7�������$I    `$�����'�رcKA�������+5jԨ����2�=�t�����˗K�^x���r��/ڇ�buttķ��������o�"�b�hC.�{WKK��  ���; �|>?;I��Y�P�ңE�~��8w�\     ��G��)S���W_]�^u�U�P���%-�p��W�G���gϞ-�ߡܥ?�ؼys?~<�/_��} e����x�}���3��̱  ���; ��q}�$WgP�8P:R4}�    P�jjjb�ԩ1mڴ���+��'O��LfX�_�0}�~T���Ϝ9]]]���Yj}�rt�ر��u�ʕ��P�n5j�c��������� � 0Lr���/]\S(K����=}@    Pm�y��1cF)�~�ז��]���ח��?>:::�ԩSq��	�w�Jz��w���X�`A,\������쁁�G���;Z[[� 0���� �P�F�����k| e)=2t�֭���     �b���1s��R�=��3&�����Ν[�w����+mxO�$`8����ݻ��#��o�=&M�@Y�>��lhll|Ϻu� `H	����r-^���j(;��Ν;����    P���4�>k֬R�=��D��:uji�����˗KA��G����>0����X�~},Y�$�͛@Y�������l�#���_ `������H����c��C���͛7��     �l��ѥ@��ٳ�����2nܸ�3gNi]�t)�9R*99{�l�p�;v��ӧc���Us�T�������r������y  CB� �H���$I>@Yjoo��[��6�    *Ք)SJ����痚���Ə�/.�3g������������0���F��o�=�M�@�J3v�%��Nkmm}( �A'� �/�����x} ���>�H���=�\     T�����馛J��k��6xy�N�w�yg�A�СC��}/Ο?0��S���	K�.ѧ-@�+�=3���kii��  ��; �իW��>}z[q�X e'm�y���    PiF����+�'N��:cƌ�E��K�ڻv튎�����$I<x���bժU��P���rZZZ�/�I  �B� ISSӘ����V%���n�ݻ��Ɠ�     �d�ر�dɒX�`A���WFڜ=s���J�۷o��'O����X�~}�T�o�1��՘������e���
 \q� 0&tvv~�8�-�������wuu    @%I�Ӗ�[n���:���>}z����|)����ƩS��Bl޼���[�lY�}�����9��������� ��� WX�vJmm���7PVңe�n����    P)Ҁ�E�b��ť�v�Nt�[�����a��ѣGK��U�VŔ)S(K3f�Uk׮]��C]
 ��p�+�x�:������ �F�P��;w���    ���x�q��ǤI���3cƌ�����å�{zZ(�����w��ҩ�����$I򮾾�o|�c{�g?��� \� p�d���{{{�gq\@����)�^    *�ԩSK���A���dbΜ9���*{��-��`J_c;v숮��X�bE�3&��$���Ǐ_�������r: ��L� ������L&���Qu�����R����@     T�ѣGG}}}��9TS~Ҁq4�?~<��q�ԩ��v�ĉX�~}�/ӦM���^\�����677 �5p��(��.~1�>3�����[�l)m�    T�3f�w��&M
��UW]o}�[c�����3ϔ��a0]�t)��X�pai���PV�$I���5k~��G9 ��&� �A��te&��Fq��,�={66m�.\    �J�6����s��	*O���8ᩧ���Ǖ�2��$��{��NX�jUL�81��2���fC.�{kKK˾  ^w x��T(��8N�,8p v����f     T�����뮻Jm�T�4d|�=�����F���Swwwlذ!V�XQ��PVn*�ǲ���Z[[� ��	�������V(�\'0��c_�n�ǎ    �JPSS����t���d2AuH�ܧO����w�̙3�)}>��0{����[K�+@٘^�~_��������T  ���; �Bk֬yW�$_*��vgϞ�M�6Ņ    ��m�ozӛb�ԩA��2eJ��mo+��ݻ7`�>|���~�w�N ��5���|>������ �l� �
o<W'I�ߊcm �.ݰݾ}{
�     �3f̈7��1v�ؠz�5*n������kK�����)-ڰaC,_�<fΜ@٘�$��r��/����}  /��; �L�l����?ߟ0��#7�m��=�\     T�[n�%n���d2��0{������G�������Iz�m�����[���&��0��Ґ�[ZZ� �O%� /C6���L&��h�Y�@�n�^�p!     *��ѣK��{�낑�k���������ǉ'[zn�<eժU1q�� �Bzt����G����* ��H� ~���}I���p;����غuk    @%?~|���o�k��6�Ǝoy�[�駟�}������ذaC,_�<fΜ@Y�$�����Z[[�, ��$� ?A.������`X�������=�\     T�)S��=�ܣA�������;b��ɱe˖H�$`0����Nŝ;wn��ח^�����d>���F���|6 �K� ^B��������͛7���?     ��뮋��;ƌ��-Z�������Q(����̙3�j�*?���0���$��Mjii��  �� �co$�]��;����Rs���@     T��3gƛ���=�#y~�ٳg�B�>�h�Sl��ݱ~��X�re̘1#�a�)��_lr��  �	w� �Oe���J�dm �&��O���=�\     T�o��n5jT�O�����Ć����쩧���s�F}}}���0�Ґ��f�W�����  ~H� ��4���I��6===����>     *ɜ9s�g~�g"����]w]����\�Y���/`(<x���jժ�0aB ë�wCS.������ ��@��իGM�>���$�� �M�؞6�k�    *��ٳ��yU���J!�o}�[��2gΜ�o�۱bŊ�9sf ���\.7�����8' #��; #^SS�����?/�
`X
�رcG:t(     *��^�:�v^�iӦ�=��Sjrrg����M�6łbɒ%>�`����|���9=u^��M��-mn�����n�as���xꩧJM!     ��n�7��QSS�ZL�>=~�g66n�Ce߾}��4�V��q��0|�$��-~'4455 F(w F�����1c��e��]]]�y��R�    �Ҥ���;F�p%̘1#��x���Ӑc�PI��lذ!��Θ:uj �'�������LSS�o	�0R	�0"o�ttt|>I�_
`X8p v��i�    �HW]uU�m{�h�ݹ�f͚.\�g�y&`(��D�=�X,^�8,X���XWW��իW�_��c= q�i0������/d2��0����K��ǎ    �J4v��x�[��ƍK�,��/�޽{�R�P�]�vEwww�\�ҏx`%I���ӧ�M�-�� ��_� �(/�ۿX���;�|<��S�+    @%JÞo~�c����)�M����C�������w�y��;^���HC�&��H"����b��K����t~۶m�w    �J��=���[&����+���oƹs�����?7n�+V�̙3��vvv�455}D���B�����q���_`H�GY�ܹ3<     �l���1{�쀡R[[w�}w|�߈������mڴ��ٷlٲ�/�a����3���𑶶6_ T=w ��ڵk����~�8�5�!u�ҥxꩧ���;     *Y�ھ|��6y��x�����w���Ç���'��7n\ ��WjkkӐ�����v� T��݄^x᫙L��R]]]�y��|�r     T�	&�Z�kjj�Í7�����Sa��>}:֯_�V�*���3f�W߿nݺ ���; U+����~�8���ڷo_�޽;�$	    �J��d⮻��X̰[�lYtvvƩS���/�O<�D,^�8,X��K��]���{������納P���J��0<���b˖-q�ĉ     �K�,�믿>`����_��ף��7`�
�صkW�={6�/_����wN�0!����; �H����O|b�K��p�[2�?�|<��q���     �S�N-�fC��8qb�y���c��cǎŹs�J��ɓ'0�2��;���c�ڵ�{衇. Tw ���>���.]����� �Lz��͛K�     �`����7�!jjj�ɬY����=�90����7Ɗ+b�̙�����~��{��%M� Tw �FCCÄ��ڿ�vR���ݻwG�$    P-���)S���;�#:::��ŋí��?6m�,�%K������M�4���{�{���� T���S���H7+�y���     ���k��E���1c��ʕ+��(i)ҹs�bժUQ[[��I��&N��6��O��j �@�{1������ �ą��'�����     �&555q�wj ��͚5+�9�����ԩS�aÆx��_�'O`H�}	_nll|ߺu�^ �`� T��k׎������xO C"ݘܼys���    @���[b�ԩ���;'Oڳ���EI7n�+V�̙3:�L��B!����; �L���U�!�������s��h�ݻw�G�    @��4iR���T����ǭ��[�l	('����iӦX�`A,Y�ĩ0�ޙ$�ohh�P[[�_@P���HMMMc�����8�3�A�nB���Ǐ    �j���5*��,\�08�Ν(7iyR��\�jU���04�$���{�/���>T\� F������;;;�p��t�1�O>�d���    @��>}z�t�M�������6��S�N�^����c�����wvv�!��Pi��(/�ۿX1�A�n8n޼9���\    T�L&��~{@��9sf̘1�I����Pi�ƍ�c��W`��Jggg����!w *��; ��p���{t�q�;w�L��    �j6{��:uj@%K��'N���O����M�6łbɒ%�Cb��!�_r�R�Pj;::>��d���*
��3�D{{{     T����X�ti@����c֬Yq�ȑ�r�o߾8w�\�Z�*jkk���HV�^��_�� ʜ�; e�x�5����ϊ�/0�.^�O>�diS    `$�7o^\u�U�`ٲeq���R���S�Nņ�������w/ )N4�%1�dq%YN��U��i��ؤM_��-K�XV��$M�Ǥ/M�:�S���&�;�e;���v�bk�$Q�$�"EQ�<�L�t�;�ʕ�H������ko���Z6�����b�q�W0�r������w/[�쟥�/
 F4w F�,�����I��\ C���ñf͚8}�t     T�����3gN�X�mָ馛⭷�
麺���g��{�7��� ��#ɲe����; #��; #Vn����b�$?��ڽ{w�[�NE    ���v�m1y�䀱䮻��۷{�Ϩ���/��b466ƝwޙU�`��ӎ���t^��$ `p`��544<.�C+=����_��[�    @%�B��g�k�L��_}�ر#`���U;v,�ϟ����Y,{Z[[ ���r�Tk�$�"�!�U�x饗���    Pi� �ԩSƢ9s��3�<x0�{������&�!��b������� Fw F���?�;���!����W���Ǐ    @%��;ƪ3fĕW^���N���{��^�w�}Q[[���W�B�h[[� A�Q��⯧����9t�P�Y�&zzz    ����N2��y��J����bŊ��{�n`h�r�_+
}mmm�) `�p`�(��>��m Cf����ꫯF�$    P�fϞ0�]}��1u��8q�D�hS*�bݺuq�ȑ�Ї>�|>�����~��!��
 ������WY����_��[�    @%�0aB\{����[n�W^y%`�ʊ7uuuł���:������K�P8����; ���; �]z�ԔN�`H���ŋ/����    P��oUUU@%���[��^+WÆ�*{���3���]	�!�K�555u-_�� .#w .�B��Hz������ŪU��    ��,��b�ĉ��v�
�N�<�>�l̟??2�$I>_,�[[[�8 �2p�ijjZ���n��0�jY����;     ���1mڴ�J�Uqpg,��ye�����hll`�d�n����tj���O \� \�b�$�R�sc��۷ǫ���q     ���o�4W]uU����ӧF���צM��]�������R�!R�oOeَ��ֿ f� �������?
��`ЕJ�ذaC����    �d!�k��6���r�����c�֭cŎ;�ĉ�`���`H�O�W���nkk�^ �0,`X577�T*�i������2�^�::;;    �����+� �X�E��g�y&.\ӧO`HL��r�hnn������ ���; �&��y�T*�Y���Yֆq�ʕq���     ��n�ᆀJ����&M���$�7�����������!QS*��nnn�і��� �@��a������p{M ��������===    ��������k*U.��뮻NwƤ����;�3�K���jnn�ᖖ�� ���; C�X,6�7:�N�3T��틵k����@     ��jkkc	��k�pg�J�$6m�T�z|�=��7u ��6�755=�|��� CH��!�裏^�����t���ڶm[lܸ���    �3���*]CCCTUU)�Ø�cǎ8u�T�w�}1n�X�k�$���ŋz��'� Wr �G}������4�R)֯_�v�
     �M��������e����������555�[Ə������hmm= 0��/������t������իWGggg     pn�&M��3g��fw*�����{��^,\�0f͚��J����/>�O|��~��N 2w ]ss��R��rN ����+V�Z'Nx>     p�x�UW]P)z{{�^�{�7��� ݂I�&}�ӟ�����g>� 0��T�=�ؤ������ ��Ç˕�{zz    ��W__�;�O��Ǐ/��J�X�vm�<y2�� ��O��zss�O���x���p`�,^������$I~8�A�w��x��c``      �0uuu�#��Emmm�۷/��lٲ%����{�|>��I��o�ӗ-Z���z�)/�� ��F�jܸq�޸�� Ͷm�b�ƍ�C�     ��TWW�+V?�u5p��ܹ�\�}��N��I��g��/�=]���? .��; �!����xz����]�u�b���    ���*Ug��Ȏ�T��g�y&x���2eJ ����c���� \"w .Y�P��$I�E ����/V�^���    �����5kVy��T����x��g����{�'������_ �� \����W������ʕ+��    �4ӧOཪ��˕�O�8P�z{{cŊ��8���� կ655�Z�|�g .��; �X,~*��} ��ȑ#�jժ���	     .��;|�3f�S�J�R�����c��;�,w6 G�$�Y(:���> p��(��ϧ�o0(</��b���     �nܸqq�W�~��]�v�u��r��y��E>�`P�R����tb���_ �@� \�b������t���A�s��x�W�U"     ӦMS��@wx��{���,/\�0���UI�|)˘���~' ��pA�.]�0��8��A�y��زeK     0�To�3s|��uvv�s�=�����0(Ƨ��b�GZ[[� �'�D �[SS�]I��E���%ɪ���꫱cǎ     `�M�2%����v���x�g��� O���[K�.}���# �<�p^��������%���_|1<     ^8�q���ĉ�����WOOO<���1�����+u�|�;�B������ � ��9577וJ�o&IrU �${ �r��8z�h     0t&O֐�&�"�,+X�f͚�����o`P\�����c�}������ ��pଚ����vz���%�Z�Z�*N�:     -���M ���|�R��ׯ�����;sz{{��P(|����d ��pF�=�ؤ����s�܇�$�.���c*     z555��c�ϖ-[�������r\����'���?���� ���@�-������t�� .�޽{c�ڵ�*     ��������ل	8?�v�ӧOǂʿc�K���>�$��/[���Ët �G������2���� .ɶm�b�ƍ�O    ��8qb g�8�����=�\<��1iҤ .M�$�����H�, �5� �O�P��t�D �$����    ��?~| g��;\��Ǐ�3�<S�O�6-�K�$I�X,lmm�� ��B���Ho~)�>�E+�J�v��ػwo     0�w��l��s���x���c�Q[[�%��b�x����s �'�������Y�$��E���U�V��Ç    �ˣ��:��p�����+V���s�Ƶ�^�%������˗/�r @��}�b�'�$y"]��(��ݱr��rkB     .���� ��q�&����K/���v�m\�|�$_(��[[[� T<w ���yAz�����\�'N���N�
     ./�]87�	��7�C�w�uW�r���%�Z�|����o���� *� #@���'?y����7��� .ʑ#GbժU���     \~��pn�|>����[o��ӧc޼y�-�4W$I�?�,Y��O<�# �X� ����ꁁ���S] ���#V�^���    �Ƞ�.��.��{�Fooo�w�}Q]]��I�䪪���,Y���'�x�= �H� �����R��?��\�ݻw��/���`     #��.���_VkŊq���Ǆ	�h�VUU}�P(�h[[�� ���T�e˖�ooo�Z.��'�����o�k��&�    0�J� ��qC�ȑ#���ƃ>�'O����r_^�l��M��� F��¤�����?Lo>�Eټyslٲ%     �'�sp������=�\<��1mڴ .�O����~:��t��� � &�����\nQ ,{!�ꫯ����    ��k`` ��p��u���x���c�Q[[����r��X,�hmm�w@�p� MMM��$ɣ\��!�K/����     F6w87�	����X�bE̛7/��� .گ�Ŏ���� Tw�
����$�\����X�fM�!     �T��sp���i����M7��E�l�P������ `�p� �b�'�$��t���d�W�ZG�     F�,D����O�$��+�ĩS�bΜ9\�|.��b�X<�������&�0�
�����p·���+W���'O     �GOOO g'��o�֭���w�}w�r���E���777����� `�vÊ�bc:�E:�pA�?+V�(Wp    `t܅s�.��۷������G>���]Q*��Q(hkk� �I� c��ŋk�$�F.����tvv��ի��     }/�ss���o߾r���Fuuu ��\.���K�~���? �9� c�c�=6�����ty[ d�����/F�T
     F���I��We\83���ʊn���q����ĉ�`wVUU�Iss��---ڒ �1� c̲e��_L��pA���k׮�$I    ���ԩS1eʔ >Xv� �WMMMTUUpq�$��t|>]���?�1C�`�����\:�t d����ꫯ
�    �'O�p��Ȏ���:�̙3'n��� .��
�����~% 3�Ɛ����$Is d�֭�iӦ     `����
��#pyd��,XӦM`p�r�_.��[S�� �0F455-J��7� ��     c��.�Ytww0�������{���:�A���bqOkk� ���;�����P�T�B��p�6l�۶m     ƞ�'O��l ����cΜ9q뭷0d���b������k�QM�`�+
��J���ˉ��$Ib����s��     `l:~�x �رc����X�`A̘1#�!W��?]�d��O<�Ď `�pŚ���J��7�e] �%=f⥗^�}��     c�ѣG�Or�\ ��л����{���� �͕UUU��c�}䳟��� `Tp���I===O�r9=��<Ě5k����    �����'N��+��"��p�����cΜ9q�^��erGOOϟ677����' u�F�E�U��_��r8/}}}�jժ8t�P     P�9"� ;6��QSS��Ϗ�3gp��r��J���-[��Q
 Fw�Q����sI��� �KOOO�X�"�;     T��J�7��d�N�<��ꪫb�ܹQ]]����;::���/ ���;�(S(~1I�� �Kn�����    @e���/;.�$	`������;���1��
�������!�0��şK���y���*Wn�f     *OGGG9ț��xGv\ ����&�ϟ3g�`dJ�?W,w���~# �F�B�0?��{:<���Ul���O�     *S___=z4f̘�;�a�\u�U1w�ܨ��`D�JǗ���hkk{) ��F������$�v��pNG���+WFooo     P�:;;��p�K���cΜ9q뭷0j��r�?-
���v #��;����|E�$O��� ��СC�jժrU     hoo��n�-�w�)�fҤI�`���9sf ������B��Ѷ�����%�0�-^��z``�k�\�8��
On���     �8p �w8��\y�1w��?~| �S.��p�$_Y�h��yꩧ�I�`���nI��pN��     |����r��3fT�}��p���|466��ߞ�c��������~+]~* ��F�b��o��_pNY��5k�D�T
     �����+�N�ˊuttpa&M���ϏY�f0v�r�G����Z�|yK 0���@�B��L���9	�    p.Y����
�d�	.ЕW^s�΍���0�$I�٦���˗/: Q�F���y^z�?�e>���*���K�Mg     ��tvvFoo��"m�����|>���q��gU����$�b�Px���� `�pA�,Yrcz���tY�Y�ٳ'^~�e�v     �)��{���[*Q�>e׮]�ۤI�b���1k֬ *\.�?����kii� �� #Dz�|E�T�Z5pV;v�W^yE�    ��{ܩT���q�ԩ ή��>�Ν'N��\=00�t�P�h[[�� �p/^\]*���.�
ଶo�����p;     d���q��i�E*�Ν;8�|>���q��G.��������ˋ-����zj  ���F�q����t�x g��۳��     p�J�R�ٳ'n��րJ�ڽ{w lҤI1���5kV �'�K:�� �p�̊��/�Ӓ ���7ߌ�7     \�����;�&�^��������ży�t� ޕ$�c�B�����e#�p��?�N�1��ںuklڴ)     �R<x0N�8S�N�o��V ���b���q��� Uz^�lSSӛ˗/�v pY�\&�B����2�m޼9�l�     0�m����*��ӧcϞ=�@V�}�ܹQ__ g0.I��,Y���'�xB�y��@��2(
W�r����� ����_�7�x#     `�����q��wG>�c_��}`` �w���ży��!w�s����������ZZZ:�a%�0�y��N�O�q] g�aÆr     L��ݱw�޸�:�j��k�w�r���;�����8O7|mٲeKGo 0l��Wn��ɿ��8�M�6y�
    ��ٲe��;c޾}������n	�����p�r��CO��O �F�`��_N�����p�֭[     �����СC1k֬��j�������6,XP�\�Z(6���}6 � �$����t�� �H�    �ᒅ?��EG�����T�\.��v[�y��5��J�%�)
�����< r� � ���'���B������    N�v튮���<yr�X�z;�,��>o޼����A���r_ljjzp����!%�0�
�������Q8�v     �[�T*���$�%�ƍ;vT����X�`A9�0�&I���%K�{�'��!#�0�y䑉��'�.�$�    ����oƝw�555cņ�8��466���\. �ЍUUU_knn�XKKKO 0$��Nn��ɿ���@��     \N�g����N�<o��v@%ɪ�ϝ;7`�|�T*�N:? 	w�!R,�]:�| H�    �� ��~�wĔ)SF��^{M�v*Jmmmy��ĉ`�������˗/�L 0���@�P��t��@��     �Yx�ƍ�p����nǎ�;vT���Ƹ��;#����$�njjں|���A%�0Ȋ�������>��     �4o��V̞=;f̘0Z�_�^�v*	b�ܹ��� �Y>I�?ljjzp����A#�0�}�ц���?M�5��믿.�    ���$I�]�6>���F���={��u���1���8qb �S�k�?onn����� 
w�A�x����������x�,���o     �D�ݻw�u�y���Um��ƺ�o�9>��E.������ח-[�7�� \2w�A2~���$I>��lذ!�m�     0��[�.���ꨪ�
-��G��n�ᆘ5kV���Ƅ	`�HGG�M� ��	��b���$I�E �q�F�v     F�'N�;��u�]�Awww���kcݡC�bƌq����|�W�T,
���~' �$� ��X,��t�� �'{	��o     �YW�뮻.�O�0ҭ]��\�ƺ�'O�����]6>===Q[[�\. F���Բt��-�?����Ep�K�,�1��8�O�}�l�o��F     �hR*�b������N2��ݻ7v��P)���cʔ)���]]]������1n�����R�����Դ`�������
�"
�)�\��tY�{���[�y��     �Ѩ���ܡ���1`$ʪ��Y�&��$I;v��o�=Ə_>���W��^SS #Hmz����?��|�3��
 .��;��ɥ~/��
�=�p�k��     0��[�.��ꪘ:uj�H���/ǩS�*���@l߾��)벑u��*�O�6-f̘ #�=����#��#	 .��;�Ehjj��$I�YL�v     Ƃ���x����|>0R�޽�\p*U��#��~�5׼�gǎ+Wt���s�F���X,�bkk�o D����?�$ɯ�������     ����7Ƈ>���� ��^�:��eU�'O�ӧO�Ϻ��������������-
����< 8o� �����R���2�����[n՚$�j    0�lذ���\N�{�+VDOOO �v�I�&ń	������������6jjj`��r�/���[[[7 �E��<���J������ ޕUAx饗��    ����+W������'\.Y7�������عsg�v�m����F]�T*Wx�6mZ̘1# F�����b�8����P pN� �a���Y����qs ��	�    0�uuu���?�������z��x����u����k��wǎ���ި���|> ��M���e˖�D:���p8�Ǐ�\�$?��:::bժU�
     0�e��_y����?0�� �+�3��[N�<���www�7�444Duuu \fO�Y�)�? ���;�9
��$I!�w>|8V�^-�    @EٴiS̚5+����������<�L���pf�w���0a���.;�����������u�P������ ���΢X,ޛNO�#G����d�     �Ҭ\���̂�0Բ�Cٻ��b�������|�}��joo�iӦ}`�w����_�t���� �	�����>�����g�rR eǎ+?�n    �Re�ȟ}�������<yr�Py��cǎ�����سg�Y�ld�;{{{������ �dbz���ŋ�=�䓝���|�e˖�����r��6���Ǐ�/�P~�     �,Q~��ߍ�~8Ə0ضm��7o��:t(�L�3g�<��d��}��ECCCTWW�erCz��E�=��SO �!��:::�k:�p e'O��+V�    ��eU��{����QU�TY�5k�pqv��5551q��3~M֍c���Q[[[�Z���o����z:�b �� M�P��tj����+���8}�t      ?p����3�zHȝA����:�&I��)�J�cǎhll<�9������6mZ̘1# .���Դ~���_ �%��W
�{r�ܓ�����ʕ+��    ��J�Yԏ|�#���.Vggg<��3��������]�vō7�xί�:rd�����lV.�\�$�}ɒ%��x≍@��;��=��c3ӛ֯�K�� ���W~ ���      �l�Ν1nܸ����.Ƒ#G����p;�츚:uj̚5�_��������Q]] �lrUU՟��y���� w�̢E��z{{��.o
 bժU�j     �����[QUU���Wɝr����˿��ri`pe]6jjjbҤI��ڬ Xr���-�0�1�hѢꩧ��	������s:=@�J�X�fM:dS0     \��[��C�<�@����s������I�$�o��g�.oB:��]iGGGL�>=�M� ����������@�p*^�P��t�W��]�6<     ��۱cG����C=t^aJ*ׁ�g�)�{�NOOO�ڵ+n����g�L�9R�x�Usוf�\(^mkk�j T0w��-]��C���ҥ;RH�_�>���     ��۳gO<���{uuu�_�{��x�b`` ��w������,��WWWWyJ}}�K�pʥ~�X,nnmm� J��XK�.���翞.'6l��;w     p���������G~�Gb�d����-[���/�\��l�QMMMy����{v>ohh�����0����/^�x��O>y, *��;P��-[������tyK ���Ƕm�     <Y��o}�[��̙3�ʖڳ`{p�_vn߾=�������}Y�����G]]���.Qcuu�,[��北 F��H�����~"�r���7�     `�uww�w��x衇�ꫯ*S___�X��\A�|z{{cǎq��7_��e������6mZ̘1# ��������t�� �0�@�Y�t����r�@�ܹ36l�     ��������wcΜ9q�=�D.�*������g��cǎp�e�bV�����������Z�r`X$I�k�B�嶶�o@p*J�X�!��G:ο��Q{�����     0<6m�G��|0Ə�}Y���r{��9�w��'O.����U>�����q�W����r�/.Y�d�O<�# *��,�b<��#���%I2+��e	֮][n�     �,T��o~3>�яƌ3���T*�m޼9��iǎ1{��
�����������.&N� ClfUU՗���?���� @���'OnM�dn@�;|�p�Y���`     ~'N��o}�[q�]wŜ9s"��c�ɓ'�U�;::����Ν;�[n�����ƬY�bʔ)0��J�Ϧs! *��;P���'I�
w�رX�re���     p�d��W^y%8>�`L�4)��~��x�����Q�����zCC�E}�1���3���t� ���B��b[[��`�pƼ������s.���/��      #Cp��7���w_\�������/��R�ڵ+��e���YG�K��*����E>������onn~���e} �a����t�����ӥ�T�ӧO�+�gU     �����'�{�kb���%��Ν;�U۳���'�¾cǎ�={vTWW_��d]�MK���1n�H0d&�J��|�S�����}�h �Q���1kٲe����/�˛*X�sŊq�ԩ      F��{�����}���e.�F��{�5kʁV`t˺`g!�[o���νY���"|CCC�?> �ȭ�y���wӑ�$��Y����>����
600P��~���      F�,d�v��r�r޼yQ[[�,Yq�M�6��͛�k`l8y�d<x0����K���mr������� "�P(�B[[�
�1H�����?V*�~%��e�����
     `t���o}�[q�7Ľ���'O.��;wƺu뢫�+��'�Ȑ�o�N�zI����moo��ӧ��P��r�^(ֵ���� c܁1��G�������eU@[�~}�۷/     ��+T�ݻ7�̙��~{TWW�/�f��l�0ve�����`�o�=Z��>k֬ �\.����s[ZZ��"��)�<��������K��h7n,?�     F����x��Wc˖-1{���;݇Ih�޻��#3�";�f�Zo�喬:�%މ'ʟYWW�|> Y}�T��e�>��� #܁1e���-�4/��������o     0�����k��V~�Ut���[c�8���¡C���[g��ʓ�����W_}��|^www8p ��띷��p_gg�o�ss ����1�P(<�N�<���޽���     ����ڵkcÆ�����&M
.]h}�7Tl���=�L�W\qŠ|^ooo��Ur�8qb �$I�������?�1@���9��P��,�֭�nZ     ����6m�-[���7�\�O�6-�0����cǎؼys;v, 2�{��ܐ�[Ǐ?(�900���ڬC} ���P(���ֶ9 F9w`����?=����+�&�B9r$֬Y�R)     �ʒ&�|���9sf�v�mq�M7Ÿq"g����~��ضm[y� �_��_�o��������3��|GGG�������`M���_Y�x�}O>�� ����^ww���tg@�:y�d�Z��\]     �l�.�ɺ�fUݳ�{V)�w�>}:v��o��V:t( ��ԩS�o߾��k�s�=Z�g���
�$I�C���-���(&��j�B�_���P����+V�PU     x�,4��o���ɓ�뮋믿>�������ƞ={���,��#.p�������������U������| �O
�����> ���;0j-]��C�\�*�ؾr��r�      �3��[�l)��S���_u�U����ƍ����c��a�l<xP��d�&�I�&ń	�s��f���/�ܫ��`0�r�Ǜ��׷��� ��ؼSƼB�0%��J��P��]�Y�={8     p�N�8�nؽ��������<s��Q[A����\a9�g���'O�`����ܹ3n��,8:���u���!��'� �X*�����<����x �2�����,�N:��@Y��_|1:      +kf��ld�j�f�*,kkkc���1y��i�.�Y��]IGGGy��!눱w�޸��k������&���;Ͻ��Ԙ^�=��? ���;0���O��?�P���Z8p       S����Ə_�Ϙ1#�M�S�L)/�9� ?����Y�4�:�؏=�.��$	��!�T���s�`��m��g���p�r���
�ﵵ��N �"����^p�O���PY���۷     �p���������&M�Tyf!�	&�g���rE�Luuu�*���fV�8q����������;N�>]Y�=�Z��h׮]�s`v�
G�)�gΜ �*���b��Rkk� %܁Q�S�������/�ˡ�C�n��ݱy��      	�
�� �4Y�<+L���X��3�?^��SWW��&!���e���x��O>�� ܁�"����{�|S@���u�l�      	�>{��믿~�~ƩS����Q__UUUp	n����B:��t$0�	��BSSӿN��*P�3����v�       ���)S��̙3��g����r����K�SMMM�\�|�o�'��x�b�$I~=��>}:V�\}}}      �Ȳ{����'����g!����?~| \�$I�K�Px���me �`����x���tz*�Ш8�C�+V�[�      0�d��w��������������������Hչ\�KK�.���?~$ F(w`$�UWW�n:_Pa�� k֬��Ǐ       #WV�l׮]q�7��I�$:::b�̙1u�� �H7���/��O�#	�H�����c��w*�����&       ��9R�Ϛ5kHNr?t�P�#xt�H?Y(�mmm�`pF����y�M�oT��7�w�      0z�޽;jjjbҤIC���n�Q[[�\. .Tz��L�X\��ں. Fw`�)
S�$�b�Pa�o�o��f       0�d�ճw��gώ���!�y]]]Q*����.�����{����D��U\��w����
(xko�t�=�t������T���n'&s9���I��'��v�ĘL�y�>g�L&ݭ�hk�-wD[��U�oUE����Ac� T�޻>���=�Z{����k����ފ �H
���/���O�""��\.��aZ@�o߾ظqc       P�Μ9�ur�4iR�������Y�رc{$T��)���X: ���;PT������1��5k�d+�      (]��oMMM�5�G~_[[[�ݻ7ƍ���p�>�����ҥK�8 ���;P4f�����cҶq���Jttt       �oϞ=1x��z�ٳg��ދ1c�����b���'/^��'�� E@�(
�?�xukk�_{���DZI���~7ۦ      ��v�ޱcG̘1#***z�wvvv��������A��"T>C�������˗�
�^&�����'
��}HZA���'N�       �Kjx�k׮��kz�w�`}sss�1"� afee���G��	���������>f���q���       �<9r$ZZZb���=�;S�����Yӵ�Ç�E����Ɨ�.]�Ћ܁^U__?�0�a@�y��سgO       P�ҳ���Guuu�������̺�\�|>�Ն���MMM[����f���
7RY8Ї�-�nu       �W�ܹ3�O����l\�رcY'��� ��!���%K��Q�� ��@�������0;�9p�@���      @���֖5C���k{�w�<y2��B�p涴�|�0�R �w�W,Z�����Ї?~<V�\�M       з�n����1f̘�ݭ���o߾;vl���/ .�c/555�� �a�@�[�x����?-������W^����       �oڻwo<8jjjz�w�����^r�������]����q�ҥK�@pzԒ%K*ZZZ��p8"��H�S�=m�      @ߕ��c�Νq�u�E��=����8�ɽ��* >¨B�����׾v6 z��;У8��}}Ȇ�СC       i��;vĔ)S"�����?{�lr3fL80 ~�|>�رc�p���C܁S__K����![�l�ݻw   py0 �F=u�K���H�%���;�/���K��𾢢�ܖ�iL?�t����]N�>��i��U|��t��9s&S�!u�;������I燎Bz=�7���ZS����3   �]'N����欓zoH�����ѣG��������������Ŧ��U�܁Q___S��P�}D
����   }]
�4(�w�]��t�ƮJ�1�S`=��u\�[��t��� }W�=U:N���]���:?u�T���f��  �Ҽ��{Q]]555�����閖���+�- �҇ğ?��#7?��S���	�=��\.75��8x�`lذ!   �ܤ�y
��T?�8=�O�λ*u�K!wz_������R����`S� |
�w?~<N�<��w�:�  ����Ν;c���0O;�������vРA_)��@7p�]CC��������ʕ+=�  �d�L?�R�NO��JwH.6(����S�y�T)�u�*u�7�  �i��r�2eJ�r����ԨQY��"<��ظb�ҥ �ȓ�[-Z�hra�À>"m���+�d#   ��F??�>dȐ����t����RP�k�ą�������5�׏;&  ��t�o߾?~|���to6lذ>|x |�|~٣�>�ݯ~��;����fɒ%�[ZZ��p84�HSW�Z�M>   @wK!��@:�СC���;��b�R��!>u�ARW�������) �ȑ,�~����5!x  ���߿?[����K��>z��ڍ�C+|��e]]ݝ˗/o�n �t����%�\>b���q���   ��!=l�
���j)�^[[{n�u��y0@R�;�C&�ۻB�)�~���lL!�� � <  ���ޝ;w�u�]UUU���O���r�n-|V�߅qI tw�[,^�������G�����;�   \�`?�{���]��pyTTT�[,2nܸ�~
����)��)����|zO   �	gϞ�B�S�N��^���s ������666~k�ҥ�
��L�����/ooo��¡e��	{��-[�   |P�6bĈ9rd�u=�Q��G
�w-6�ꪫ���)ܞ��������СC٘^O]  .��'OfϠ����K��R��ѣGg���AE>����=�؍��{�w( .#w�kkk�j.����.^�֭   ���M���	-m�����8=@���������t�k���}�u��8�U�+J]�
  ��hnn��.��zZt��)R��Mhkk[^�e$�\V���u�|�����z�Z�*:::  �򗺝�éR��ԉ=��SW�������S�Ly�{�O��B�)����=��S��4�  ���޽;�_�p�\.����p<�E�����G����
��D��l�������\+W�̶�  �|��j
����)Ȟ�S�=����p�Ң�q��eu�|>Ǐς�---Yuu�ooo  ���ٳ�s�Θ6mZZ��[{��H�# =�����Դ5 .wನ������Z8�lܸ1�  @���Ȟ§�{�q���M�)C��jҤI�{�ĉ�o߾,����=�S�  �{N�:{��+���#6u{Os)����ߖ,Yr[�l]\2Oj�ˢ�������-}�[o����  �4TUUe��Cޮ ���㣺�: �IMMML�2%�.i'���=�S�=���ѣG�n�  @yknn��0����E�Æ������---�Z5 .��;p�������߿?6o�   �������Ͷ�3fL6�0{z�{�[y��ٖ>�RM�>���O����{
�tu{?s�L   �e׮]Y�����ԭ=��]� �ĿY�hъ'�|�� ���%��������ph�+�ޱc�b͚5:c  �ԕ}�ر1nܸl�
چ�+R�媫�ʪK��J��S���K�  J[��iǎ٢׮E�)�n.(B�x�⛞x�c�1	�������0)�̵���ʕ+���=   �Y�{�#�0��W^&L���� ��t>|xV�]wݹ�O�8���޽{���5  �ґ�����'N�v�K�� E�����\	��I�������0�Ӏ2�Vï^�:N�<   t����]�Ǐ��%����)S�d�僡���{/N�:  @�:p�@6O"�����ijj�� �܁���G�2��-�^{�hii	   .�����ߴ%@wz ����od�(C�	�"�����W�-[�N \$O���#WQQ�qd@�۱cGV   \�f9r�{�1c����>|8���{��w�}7<��x  􎎎�l�{�ǎw@����rT?]�| \O���V__����Ǐ����[��  �ū����&L�+��2 ����ڬfΜ�����EsssxO��ﭭ�  ��cǎ�ƍc���P�hhhX�����p܁��x���;;;�S@�;y�d�Z�J7*  �T]]���S���W\qEֵ��0u}�w9r�H�ݽ+������� @wڵkW�5*&N� E�_X�t��p�܁�x�����Q8P�Җn+W�̺Q  ������#�S���Ç }S�H����̙3��{�ea�}��ecz  ��6l�Æ�
����ٟ,Y�d~��q�"�\����~c@K��֬Y�m�  ��0 ����i?~|TVV |���1iҤ���Kbsss��}�޽��;�����  �4�Z;=߾�{�10�x�r��[ZZ~�p�����.��ŋ�*�}1��mٲ%�*  ЗUWW��Ξj�ر�D �Ǒv�7n\Vs���^;q�Dx߹sg�ر#�=  ��K�GS'�[n�% ��/���?�lٲ�#��_������?+�(c�{�֭[  ���
��N��'O��C� t�����>}zVɑ#G����={� �"���Q�F�5�\ E�"����E�f=�䓇��p>RGGǲ�01��;v,֭[   }����4�� Л���̙3�s�w  �8���Z���f�� ElB.�����O��p~���������	(c���r�ʴ�#   �ѠA��+�8j;vl�r� �b���o��vְ  �����z������0�x�r��kll��K�~- ~ W3��裏�)_(c�|>��?y�d   ���UW]'N����:F�-�@I�`��СC�k׮x�w�:q�D  @_��{�_�>n��� (f�|~Y}}���-[�/ >��;����/�����͛7Gsss   ����ʸ��+�J]�S����" �\�1"��o�9;O�w��۶m˂�vk ��J;m߾=���� (b�r�����c�!܁������|�se,mg��[o  @�I��fO��S�=�З���7�tSV���{��,����o���  ��M�6eBkkk���hcc��K�.�� � w�y��G'����(cǎ�6  @����κ�O�:5��5p��  ����I��Lu�}�ŉ'�.���{�ӧO  �����X�jUv=\UU �*���熆�盚�v�y܁�Y�dIEKK�S�áe���-V�\i�b  �����W\qEΛ4iR�;6r�\  ���&�O��U
�477�Ν;���{z  �Mkkk�]�6n��� (bC���]�d�=�r��#��OKK�?/����Eq�[�.N�<   �f���Y��� ����7.����g�0R�}���cǎ8z�h  @�ؿ���[َ� �*���u���Ņï��p�ill�.���F@ۼys�۷/   �A���c�ĉq�5���ɓcĈ ������2eJV�������Jww  ���-[�9��#G@������а���is ��;���,Yҿ�����᠀2�w��lu:  @o:�K{
��` PR�'�-�����k׮����m��ĉ  �&-�\�fM�{�v���B�i]]���˗���	��������������ڵk  ��UVV��W_�uhO��p �_������Ļﾛ�S:t(  �T���ƺu���n�\. Ejv����Ua��y�@����T����e���-V�ZgϞ  ��0hР���k�@�.� P�***⪫��*u�<r�HtO��w�ޝu� �b���غukL�>= �U.������g�-[�&�>M���ŋ�����¡'픥|>�un?y�d   t�ԙ=�S�}�ĉY (O�{�ܹY�>}:v�ڕ��z�8s�L  @1ڲeK���Ƙ1c�H���r��C�~��O�g	�C��ٙ�t�D@�ڴiS�  �;�5*�z����ƍ ��8p`v=�*ur߻wo��=u�<t�P  @1Y�zu|�S�ʮc�Ԍ���_/��@�%�}X}}���_��={�d]�   .�ԕ�ꫯ�iӦe�����  蒮&L����w����Y�=uv��  z[{{{����q�}�E.��"�K�-���O>�b }��;�Q�?�xukk����'Nī��   ����2&N�3f��B� �1f̘�n��8v�X����7ߌw�}7��|  @oHצ6l�ٳg@��(�����/��'�sܡ�jmm�Ra�P�:::bժU��s  ��c���1y��>}z6�n�  �b�С1w�ܬ�?��Sw�ݻwGggg  @OڵkW�92ۭ�H]{����,���sܡjll�#��7�����g+�  .Fmmm\w�u1u��7n�-��n3dȐsa��e
��ڳg���  ���l=͉�Ř �(e�
����� �w�c������.j=GYڶm[��/  ��H�M��uj���+���WSSs��ɪ��5�~��x�7bǎ:� ���������ׯ_ �4i�����˖-;@�!�}LUU�o���)e�СC�iӦ   �aR��hj �͠A�b�̙Y	� ��B��?�#? EjREEŗ
�� �w�C�(ܘ���ӧOǪU�l�  |�����j J��a�4��}�vaw  �E������w�uW �|>�P��MMM��'�CQWW7��E�t�"�̤�9k֬�n�  �TWWg��TB� @)8p����[�n�-[���ݻ5�  �hnn�vL����	��<�Ȭ��z�x eO����������S�P��>p�@   ��ה)S�N�'O��
���wf͚�Չ'�{��^��曱gϞ  ��+ͣ�E�C���'@�4x���(��({��466ޑ�����޽{��y ��K� �jjjb�ܹY<x0�x�ؼys9r$  �bUVV��/���8r�� (6�|��௛�����	�C����\�b�p��>e����nݺ   ��Ĵi��뮋I�&	� }^
 �y�q�wĻﾛu�L��[[[  .Tj&��o~3~�'~"[P	Pdr�Z��#��zꩧ�P�ܡ�UUU�V>��Pf:::b����  ��\.������p{�( ���k�	&d��O}*v�ޝuuߺuk���  |��������Ф���o���-w(c���w�����2�q��8v�X   �oԨQ1s��,خk ��K�ܤ�nR}�ӟ��۷�믿;v����  ��M���x��g㳟�����S��j(�릦��(K�P�����ȟ.�ˠ�l۶-�:  �����1cFl7n\  pi���ӧOϪ��5�|�ͬ���ﾛ��  �|�s��#G⥗^�{�' �L�P�y�YO=��� ʎ�;���o�)e�����iӦ   �O
]M�6-��.�:C t�A��M7ݔաC���{��~��L   � 5�x��cذaq��7@��T���Ral���Cjll�'�����ӧO��իu �2�:��P�7�  zΈ#⮻�;�3v�ڕ��Sw����  ��Çǚ5k����ɓ���744�Ϧ���(+�Pf������?��o�e���3�iN!w  ��� U
��J�  �]�\.�E'���ߟ���777  }W�NL!�+Vď�؏e�* �H��}������/�d eC��Lkk�,��Rv����Ł  (]��S�f�����:{8 @�I��̝;7�4/���oܸ1=�  ����ʨ���o~�`��2dH ����{,��!�e���a^aXPf���[�n  ��TTTd]@g͚S�L�~��  �cԨQq��w�wܑ�Ӧ��v�|>  �������������������
�"���ߥK��@Yp�2�dɒ����?*J
PVRG�u��yX  %���&n�ᆸ���-� (m����믿>�'NĦM����G�	  ��aÆe;�<�����f�- �DE>��/=���O?��� J��;���Ŀ-3�Hggg�]�6Μ9  @���rq��W�M7�S�N�� �L�Ō��Ϗy��Ż��7oΪ��=  (_i����6�y��������PD�+ܯ����k�<w(��������2�̼����o  ��2$fΜ7�|s:4  �R�i	Y�s�=ٜn
��ٳ'  (Oig��cc��'�iG�b������ŋ��'�xbC %M�J������pXPF���o��V   �)ug��k����n�  Ā��|R<x0^}��x�ע��-  (/��vb�嗳�i��H����|������˗�fJ��;���c��R>��%�����ƺu�Ҫ�   �Kڂx֬YY����:  ��F����y�YW����GKKK  P>������s���>��=zt ��*++�X'��%�%����|>�ke���3֬Y��  �~��Ŕ)S�n�W_}u�r�  ��r~W��k�ƍcӦM���  ��4G��a8p ����ǂ���& �������e˖�@Ip�ҕ���X�ˣ�lٲ%۾  �}#F��:��x�ٶ�  �q�7.������_�W_}5�=  �����g��>���7�N�PTTT<Y�-T>��#�%��������e$u�y뭷  �=�[��3�.�W^ye  ��T]]��Ϗ[o�5�~��ذaC�ر#�yy �R�c��[ZZbŊ��|��@Q(�gޝ2vK�.�j %G�JP������Hkkk�[�.  �ޑ�F)�>{��<xp  @w����)S�du���ظqcv?u�T  PZ������իWǼy�����ߪ�����e��	���C	*|�.+��Dggg�Y�&[�  ��q���ܹs���)d  =mȐ!q�w��ߞ���ꫯ�Ν; �Ґ:����f]�׮]�O�6- ���B�A�>@Ip�S__��(#�7o��  �3����o��3fL  @1H.�O��U�3޴iSv?}�t  P�Ҝ�����СC����ǰa�b�ر��r�܏��ݲe��<��!�%���nT��w�Ⱦ}�b۶m  t����o�Y�f���  ��ȑ#�������믿�֭�#G�  �+�9���ĉ'���F,\�0;�m�\�+_��V|�+_�@Ip�RUU���|^k=�Fkkk�P  �^&L��s��ԩS���  P*�]�Ι3'�oߞ�)�ܹ3  (NC�����8u�Tr���>�����Fvtt����3�w(�������`)��ϱz����  �������믏ٳg��ѣ  JY.��)S�d���x��WcӦM���  ����hii�jŊ��|&���e�g}}�_,[��P�ܡ���.\�7�����СC  \^��Q
���Ⱥ] @�;vl|�ӟ�;�#֯_���ӎ�  �~��e����~;k~7o޼ �m�\ni}}�˖-;@Qp�PYY�
��2���l۶-  ��#u?���㦛n��S�FEEE  @�����O~�Y��{��^�Z�*�
 @�K�7�Ǐ��k�f��iӦ@/�����}a�� ���;�ŋ�������ę3gbݺu  \���ʸ���[o��Ç  �E�C�̙3��믏�;wƚ5k�1��  �'���ڲ��/�Æ�v��e_X�h�_<��LP�ܡ�-\��_>����o�2�&�����  ��7�|s̙3'  ��w6��k�:|�p�_�>6n���� @�H���.;�o|#ea��x zQ���������._��#)�Y(bcǎ},���	(o��V477  ��.�)�~�7f�� ���T���y������ի���� @Ϫ����5<�N��B�?��?�����jVUU�
�(J��H544\����]@�H�r�l�  �Ż��+��[o��S�f]) �3`���;wn̞=;�x�,� @�J�dC���n�+V���|�3Л����_�h���'����C�ZZ({2Q�Vck׮M�  \�d�<yr̟??&L�  �Ǘ:�Μ93�={��ʕ+c��� @�H����8s�Lv�~��l"@/\�W\V���"$�E����g����P&^}��8q�D   �_�~1cƌ,�>r��   .���t������9K�}���3  �^���Y��g�f����W_ ���)��t�ҿ���C�y��F����n@�صkW���;  �p��o�1�Ν���  t��c�ƃ>w�qG�[�.k֒v$ �{�]uR��������=�\��p����[
�G_������˗�h�C�ikk���06��<y2^{�   ~���fΜ9Y����2  ���������7o^rO]�Ϝ9  \~UUU1dȐ8v�Xv����=�0  zɨ����fa�� ���;�E��](i;�իW�v  ?@�y�-�Č3��E  @睊��;�3�N߰aC6����  \^麫��-N�>G��+V�g?����r�
�?�444�������(���T  ��IDATC�X�x����'���)�7o�nD ���<yr�v�m1a   �O�:��l���7fA��Ǐ  �O�E���%Ξ=;w�U�Ve�` �$���|衇f=��ӧ�u�P$:;;�ma�P���۶m  ��R�l��;b���  ���ʘ;wn̞=;�x�X�re8p   �tiW����8x�`���X�n]�92�N� �!��M����7��_��	�Chhh�Y~%��-��֭  �?���;vl   �'��fΜ�_}l߾=���� �������C��ѣG���>�cƌ	�ސ���eCC�_655m�W	�C��ji��J\ZU�v��,�  }Y
�̘1#n���1bD   �/-`�2eJV�w�W^y%v��  ||���q�̙,g����<�L,\�0 � e��Z�O*@�p�^����H>��'�lݺ5ZZZ  ��lO]S�=m�  ���'f�w����w��uv ��Is�)k��Ǐ�B�?��?�ͷ�;njjz*�^#����������2p���x�7  ����e֬YY�}Ȑ!  �W\qE,X�@� ���rR����������;��N|��^�;�/�_O<�N��Kܡ����NaP����c͚5ٍ&  �%UUUq�7ƭ��555  �M��_~��x�� �WYYC���G�f篿�z�=:f̘ �`Dgg�oƟ�W�C/�����0<P^{�8y�d  @_���c��y�� �sR�}���ܜutߺu��0  ���:5��������_��#GƘ1c�<����_�.]�� z��;�%K��oiiYZ8���ԍf���  }����o΂�  ��BX?�?!� p����"���gϞ�g�y&[@8hР �a��}�Һ����/_�@�p�^p���Qn(qi�����  �]�4w�ܘ={vֽ  �Bt��{�x��c��� ���墶�6ek��Ǐ���ۿ������� �a3+++S���Q��þ��/L����Հ�n$׭[��� �r���ϙ3'n�喬{;  ��1~��X�`A���dAw� ~����6lX9r$;߳gO�\�2n��� ������WK�.�@�p�����Da�	(q۶m�&� ��.�[����� ��f���YGwAw �n�������N���7lؐ�3eʔ �a�;;;�
�g�1�Ѓ$���X@�;z�hlٲ%  �ܤ�@)�>o޼4hP   t�����}�������� > uqO!�������矏#FdГr�܏466��ҥK�G =B�zH]]��|>�P�:;;c�ڵ�  墢�"f͚w�qG���t  ��ƍ��������{/^z�عsg  �}�\.���o�b������7�,��&��
�C�___�bٲe'�v��C�����
�5%n���q�ر  �r����_}l>|x   �����O��OǞ={���;�  dy�l��������#GbŊ���~6����
�2��@�p����0�0<P⚛�c۶m  �.=��6mZ�}��Q[[   �`	�?��Y'��>�V
 ��4(Μ9�N���ӵR�y��[n	�����X__��˖-{5�n%��/-]Z�ʀ���Z�~}  @)K��ɓ'�'?��3fL   �I�&��?[�n�o}�[Y�R ��lذaYn!U�z��9rd6�Ѓ��r�?X�d�m�����C7khhx�0�P�6l����  �*DR�}���  P����ӧ�ԩS��^��_~9N�8  }Q�6J�q8p :;��)M;ޤ�{
���[[ZZ)��%�n#��������[%n׮]���  ��	&�]w�'N  �RSQQ7�tS̜93֭[+W��3g� @_ӿ�,�~����<]}�ߌd���ߪ���˗/?@���ݨ���7
è�v��ɬ3  ��+��"n��2eJ   ����ʘ?~v_�jU�]�6::: �/4hP��dY�������/�< =hDUUU���-ܡ�,Z�hNa������2A @�1bD|򓟌iӦe��  �����w�s��ɂ��ׯ��� ���C�F{{{tO�n�W^ye\���S����/Z��'�|re ���;t�%K�T477/-�(a�&�СC  � u���[����  �rVSS��̝;7V�\7nL�  (w��Immm����[���K/ŨQ�b̘1�C*���t�������p�n�������%������o  ���ʸ�[b޼yQUU   }ɰa��ӟ�t�t�MY���� �rׯ_�>|���}gϞ�g�y&>���g;� �|>?g��ѿP8�� .+w��-ZT����S@	���5k��� ������p�q�]we�  ���c��c�Ν����gM �Y
����'Nd�Ǐ�+Vă>�uy�	�ϛߨ�����/_~ ��F�.��UF��M�6�ɓ'  �դI���{��,  �����~8�l�/����~ ��:4��ڲJv���֭��s�@QYY���b ���;\F��?(a��ͱcǎ  �b4jԨ,�>y��   �å��3gΌiӦe�W^y�\� �����f��t�R�z��9�ĉ���BCC�SMMM��,��2Y�dIEsssS.��P�:::bÆ  �fȐ!q��ǬY����"   �h���1������_��^{�\� �\���/�<x0;�����s���?��ln�T�r������׾v6�K&��IKK�#�/��%l�ƍq�ԩ  �b1p���7o^��l���1   >�������?s�̉o}�[�}��  ('ȮyN�8���>}:�}�����>���[>��3v�؟/.��y2���E�j�o����{/v��  PR��ԭ��;����   �ҍ5*,X;w��>5p
 �r1t��hoo�3g�d�����~��q�]w@O���_�����˗/?�%p�� �˥p��������j  @o+�_Ŵi��{��Ç   �ߤI�⡇��^{-����ɓ' ����f��Ξ=����q���ԩS���������� .��;\����م���6d�s @o�0aB�w�}1~�� �R��9O�v�߿v�l%�<I�]ۡ��K��~z����?>���N�|�܃���ά��Zz/UGG�}���z-�|:N?�� �%}�t�M1cƌx�Wb�ڵ>�����qR��{�^�v�I�w�������iU ��;\�%K�T4777�r�~%j��ݱw��  ��RSS�ul����{$� ���Yx<�S���]A��ϻ���?X\��<�>�?�����?�U \^����̙/��Rl޼9[� P���͐!C�����y{{{<�쳱`��s���QE.�kZ�dɭ���c��������������  �7����ٳ㮻�� ���F��)��V��0�����TT��˹ �+�
]�3g��?�����.@
�=����}Z�r��;� @�J�6�~0�/&���w��la@w���s����p��|,��1=��c#
�_
(a�ׯ�  @O�6mZ�{��V� �%�Ӣ�VW0�+��5��R�=��{�ߍ�B���?X)�]З�?>~�g~&�x�,�~�ĉ  (E����ye�3X�v�I�:ӧO��������ߛ��p���cjkk���0*�D�ر#���  ГF���w_\{�@���i=uU??���e��u���.)�����)�B�]������U�>����c�ԩ�jժX�r�` @�H��)䞺�����_|1ƌ����F�Rư!��&�CCC�����%��ɓ�iӦ  ����d��Ϗ[o�U�]�2���<R�`��+��$��N�QR����{W>���qS�x�R�����θ�bŊ�}��  (%i^bȐ!q�ر�<ݳ=��3�p������|�/^���'���E�-��?���*y���Y*  �n���̙3�{���� �����]A�d4hP6v���/������îs�<\W�=)Z[[��T�XGd�><,X۶m������#G� @����y�N\��o��q��@7���ٹ�0~�P� .��.\�����၀�&�8  ��Ə<�@6P��b��u���z�q*���ҤC)L�����dʔ)1y�䬑N
��� @)H�ZZZ��cmٲ%����������а�����`�L�Ex������N@�:~�xv�  �)��R��믿>M��R�=׻�� ��л>* �B�)����N�:����(�􆊊��;wn{��cӦM P��5Lmmm<x0��>y饗b̘11bĈ �f���?��/��'� �p���~�0L
(A����nݺl ���Y)�p�m�EUUU гҢ�^<xp\Ocuuu��;����ʬ>, ���=�ɓ'�~7t������ƬY����:� �4o=dȐ8v�Xv�?�쳱p�B;��m��ӧS�pI �73\�ŋO��������o��Ç  �������{�aÆ �����]!��s�o9����Q���^[[۹�{W���s��骫���z(֯_���w�]'  �U�J�K]�F��^x!x�� �N�|�W}�ѧ��կ��#	��:{��s�\u@	:z�hp ��m�ȑ�O��?��' �O
���z�ԁ��J��>J�L�a����)�~~��ĉ�9��UQQ���5cƌx��cӦM)�  �h�����3gϞ�ηnݚ-ڻ����ׯ�o�����466ޑ��}�P����5�D2  �S
^Λ7/n���ׯ_ ��uubO�R7�bO#@wH!����ϙ4���)�~���s��T *}�|�����o�9V�X{�� �b��F�8��x饗b�رQ[[ �haCC�MMM��C	��GX�dIE��+�C��(Io��V9r$  �r���k�S��T���WYY��������P����!���F�:�z�h�zO��S�=����2~�������x�ײ��v�  �M��:th=z4;O�8�<�L,\�0k�Ѝ~oɒ%7�#�ȷ1|�����9%������}/  �rHa�{�7fΜ �`ig�ԅ��A���� (5�3-}��J��ttt�/���ٻ������߭y���@`0`���Lf`��g����8�uo3t MO���4�l���9���֎��vl�" Fb�y@����_*�8@ڒ����z��,�>���[[k�~��竗�Y'J�҃33f̐I�&��{qq1�f ���MWWW�a���z9x�,X�@ `M�������C |)��W��ʊq�\?��t#����%   Z_(�����` �^HH�DFF����� ��6FGG���W���}������g�+VȔ)S��?�r)  �
�T���z�W�8qBRRRd��� C�Ǜ7o���;w�|	��W������6Z *//���   C[:5��������j��5�k�{ ��у�z�G���޵Q�M��ޛ����# |Gjj����RXX(�{   X������JMMM���O>�D����: ���� �&��/D��yyyS�N�lH7�N�>-   �@iS��y�d֬Yz�W ��|>̮

 ����ϸ�8s�!��&}��3g�L�<ٴ�_�pA   FZ߄���F�ם���{�ny��GY0d\.׷���vn۶�X ����p:���Q����G��ϰ    ���iZ�i��+t3,,�4��E� ��w���5J�x�	)++��>�HZ[[  `$�ڐ�����������Ç�}��' 0D��N�v�}��r	�?@�����k].�
l�ܹsRWW'   ��Ҁ����eܸq �J��}��}w�Z y��k�G{{�	�k�]���	 �0i�$��Ȑ���KQQ���  )�����m.��'cƌ���T�!2/77���۷�! � w�s�n�T]]�3��!��h���ӧ   �:b��{s��' x�����fv�BBB `�N�-�z%&&������v����`_z�pɒ%&�{�n���  ���� 111RSSc�����˓O>i�K `(��k~���Ͽ�o��o��������~���:Q ����G�2�   �E�gV�X�ߒ	 v�v���/̮�[� ����o'z���萦�&Z��KII�^x��u����7�  ']K�i�����O>��zH `���}�� ���p����x���Cl���   ��i tѢE2e� �
���Hd׻^r ��Ρ��-�����s���}��={�L�0���WTT  �p�����ó/^��Ǐ�̙3 ��7o��?w��yM ܁�8���o��}�:u�    �BǾkk�.���������  ��-�ڸ���闭����ziX�u���O>)���&讇U   ���=�D���2����$s��

���f`p�Svv���۷�!����#   �W���˗���� �NÉd���]�  ���p�CRz�3��=�766�K��z��=%%E���+�����
  �p��������1� N�S>��csO�
����k^���y}ǎG w��������l��
   �2�?c�Y�h�	 X���5��׸f��  
:$11�\J�MMM&�w��		1SȦN�*������  �p0�T��]!??_�,Y" 0���u_� a^@���r�V`3��r��)   ��.��\�R��� �����4���v�� F�h���wuu�fw�h蝆w`�i��/� ���BӢ
  0�BCC��Akk�����R��>q�D�!�(77���۷�#��#���u�ր����	`CG����n   >O���f͒0.�eDDD��7:�Y���] ���ѣG�Kx�A[T.\he��^[[+   CMױ4���jϞ=���$��� ��r��)//o��m�/�F�>���z���*��\�tI���   �����ڮ� 0���	�w ����2f�ٴi�<xP~�����  ��N����ܡ����]���� �B���&�}���a��Ӳ��b��#�����ɓ'   ��6!�{�2�|Z���GGG�0��	� �������&�WSS����
���m�:���;�]�v����  `��:��y��כ��z����ٳ ��_o޼��ٹs'c���ç������6Z �)..��N��   ����N[��6 0���L�]���!#  |Qhh������r�������" �N||�lذA
e���0  C&$$�<�=�>|XRRR��
`(�j��;�(v������Fy ��$W�\   @i�t�ܹ����v CM�g���$66��	  ���9��WFF�tww�Vw�kۣN��Y��:g���̔��_�]�&   CA����^/��)}��<��f� xXVNN�߱c�)|w�,�C�?�o���Vzzz���D    ���*���7M� ��6S��L\\����0  �'00�뛶���!���RWWgB����3����瞓�G�J~~�9`  �i:Ͱ����uz�>w,]�T ��4��3��Z D�>);;{���� 6��g�Ikk�   ��ic�>(3f�0� �I:bԨQf�N��O �Yzx,))�\}��k轥�E �Ȝ={�L�0Av��%�/_   O���7kgzhU���Izz�L�8Q ��V���ؾ}�n|w���[������#�(���8��   ���umm��� ���H�)�����3  ���2�Tgg�Y�z{{������O?-G��}����  <J�ht����={�!V][ Or�\?ߺu�t��#�!��SSS���lD[|�?ΨZ   �ʋ-���G�� �5iH���]׃�ݽ��^jkk���C �}��{L��| /^   O���2����jWW�|��G�n�:��xڝ���/���] B�>��_u?P�H �9{��O   ߔ��&�V����h���F)�k�]7��h ���w���5n�8p���3aw��u���O�2�O?��6w  �1��QSSc��]�f���; �$���yyy��m�X�� ���������>E �qV���   ߣ�s�Ε{�W��� n�~o�[\\-�  x���;v��4����z544Hoo� �jzh���6Fv��%�/_  �����7S�0�Ҁ���$&&
 xP����3��o���3�lْ�p8^�f�MDO�  ������C=$			 �J�h��/���  �S``�	������������% ��}ꩧ���P����  ���`����7n�g��>��L���v �?�����m۶]�p��������%��TTT�QV   �F������LpK�͵/�m�) ���ڢWff�����Vw�k��ӟ�9s星���{O���  `04இM;;;���I<(. �P�ө���p�O��ʚ�p8^�F:::��ɓ   ߡ��իWKJJ� �W�3��&   }���ͥ��Ѡ{}}�466��� ����6l� �������  �A���1%����&�!��� �-[����_'T�G�>����g�s`+������-   �~ڶ<c�Y�x1#K|���(=z�	�	  ��	�1cƘ���Ǆ�5�^[[+N�S ��v�	&�6w�9  ��!w}�փs���o�駟���P �w����Z /G�^///o���|D �����W�
   ��6+�Z�JƏ/ p3���j����_   JC�}�'N���t���6L�n�ر����˞={����  0ZL���������<[�\�R ��V���,۱c�Gx1��v���lD[ۏ;&   �~�&M�o~�" �t,..�Ϣ��̈́   OӃt�̡������M�]�4�×�ԃ+VHFF��޽ۄ�   nWDD�tuuIGG��?^JKKe��� �[�n��x���"���������z@ 9u��   ^.,,L�/_n� �m����&ԮwB�  `8锘��xsi��fw�w�SRR�>���r  �]:�����<S���Krr�)�  ����y�}�_x)��Z[�nr��� 6�   �5a���. |�v  `E77�v������{L�?.�~��ia  �U�lc������O>��kײ���a��Ϳعsg� ^��;�Vuuu���p� 6�r��"��  �}���dɒ%2}�t���  ;!���̙3%##C�{�=���  �[��������,W�^�cǎɬY� <dl```���S�wx��~������(���={ּ�   ����ч~ش� �-j�P����;�P;  ��χ������;|ƨQ���g����"ٳg�{  p�"""�$���),,���4�V ��-[��߯��z� ^��;�Rww�ܷ8l���M���   �E����{�,X��B ��y� Lbb�ij��  x}��g���ݫ��M؝	��f��?{�lJ{��w�D  �[�k�z@T�}��G�~�zS� ���E�/	�e�M	������t:s�������   x���pY�r�dff
 ��j�����xB�  �'���k�rװ�6��*!!A6m�${��#G�  ���;$�����M��<  �!Y���w��˿��Y�wx����-T ��z��\�vM   �=222d���f�( �շ1��v�� ���J�`�WGG�	�kK�N0��~ޗ,Y"��������<  �W	���(ijj��Ǐ�}�1c� x@`oo�߻���"��U����v:�O`:~�ĉ   ����/��͓��ό.������6�S   �C!!!���f���V�T��wB��6w�q�$%%�{�'�/_  ����_������]~���SO=��" Oy,''�;v�V /A�^��ri{;ui��ӧO�^  �%�����6m� �Opp�ijONN6�-   ���a������{OO� �@�X5�v��A9t�N�  �/3j�(���6�����p�B �歟�/�T�5��kdee-t�\��	}Y)//   �ߴi�d���4� ^&  @bcc���x  ��锫��hs�7NL�]/��;???3�-==]�}�]�q�   |}.���1��'O�4��z <`Avv�7_}�����-����`#Ǐש   ��Fg�O�2E x�`���F�U   �Y���S�����4ឪ�*S�Yjj������Hii�   |-�у������'���O?m� `��O�n�����$9l��;�Bvv�c�/�9�DEE����	   �+99Yy�Z�/fB�			$   :5'))�\���R]]m��ؑ��֬Y#&L�ݻwKww�   |��GvuuIkk�8p@/^, �����O���[ �#��[�~�����[lB_PN�:%   �'m���{e���4;6�A�ѣG�0Uxx� �n�<r��������_�Ν+  k	���tIKK���&�v�)�a*�h�ԩ��;�#555  �y���ӧOKFF��?^ `�����役m�6N������_t�\w
`'N�0/(   ����Hy����q ����/qqq&h�H�C x'��)eee&Юױc���dZZZ����3�N��K��5|��uikk�N�@�ƍe�޽�  ����766�<��ٳ�L��C� 0H.�k���M #�[{��C����J �����K�.	   ��;+WJHH� �G%$$H||<� /�k/d��ϗ������/RPP   {Щ;cǎ5Wss�TUU� Poo� v K�,���������C   �賂�]644Ⱦ}�d��� ��r��*//�l۶�Y �"�[�������"�����b  ���mDϜ9S �K``�ijOJJ���R���RRR��Ү#�oEuu�\�pAƍ'  ����2Wff����˵kפ��Q ;�4i�y7y��w���R   ���egg��={VƏ/&L ����ޗ��	`S�a[YYY1��+؄��h�   �C[S֮]k� �Cvu�o\\���{8�N)++��=zT������w� `O:�g����� �6�k؝flX]tt�<��3fҌ>�h9  ���]�ػw��3F��� ��p���K/������U�wؖ���[� 6���f6_  `ڐ�z�j			 ���֮�v~n��}�v�ݸq�#�\�g=��� ����`III��c�JSS�TUUImm�9X��X�`�ddd�6���  Т����,�駟��	 �����X�$�p�-mٲe���.[ �(..��   ��t����s����@ll�$%%�;?��w�pbaaa���իC��ȑ#���%AAA �?}�I>z�?��iu�����ɦM���ߖ+W�  @@@�ir���0%��&M �-yyy��m۶s�wؒ���ߺo��-�&����   �!k֬1� �Kè			fT�6v����^9s�LK�������v9y�̚5K  �E���{�^���&�M����:�N�і֢�"q�\  |[hh�9���~IMM��0�Q %���w���A �!��������݌=q�   ��t���G1�� �i��Ѧ�][9ik쭲��?�~��Aimm��;�!��; x��Vw	��tww`:Inɒ%���.���tvv
  �mQQQRWWg��^�Z `0�3yyy��m۶c�w؎��'�g6�#����   ֥!���O�ϟo6�XKHH�ik�`;m�}544�f��@�U��i�=;;[  �O� edd�q}}�	�k�;`&L�M�6ɯ~�+���  �t�"&&F.]�$gϞ��'
 �����;��3�B°����{�_�k�m�   X���|衇d����:t��v ��ͣǏ�oi/--��%V��g�ISS�DGG �7�f\\�����ڵk&L���#�H� ۆ�7���y�  ����߬�����رc%,,L `Vegg/z��W?�&��V�N�O�7f������3+   ����dY�f�6�B%11�l�h�& {���4a��{��{WW�X���h���%K �{4$���)�ƍ3�������Y�� +V����ٽ{�tww  �M:�R�W���#�V� �á-�s�	����N��Al@_���   �4s�LY�l����	��a�$$$�s	�H]]�=zԄ����o�o����; �8}�	Bz������Sb��4u�T3�ꗿ��y�  �)**��<w�9�	 ��@NNΪ;v����6z{{�c#���'O
   �G�W�\)�'O #K�����L[�n� ����3�N�z�������;t�  �G_N�8QƏ/555&L���&�H�w��7���o��  �o���1�ƌ#��� ��[�n��}q��G���������#��9s�4�   �Z�zݺu2j�(0r���M[�6
 ��C�eee���cǎ������իr��III  �����gV������_�f�����G}�d  |�>����ɾ}�d��� �0����Q��M,��;���r�~$�h���  `-ӦM3���i���M��0��M��XWmm�����Bijj_��??��� �у�z�4mt�~�:!c��3gJbb�����>�  ~O�C�]�&�ϟ7ӆ `��ٺu��W� F�������6S ())���^  �5�`�]w�% ������M+rxx� �=��ĉ���ӧO�/"� �!!!���)&�a���N��N�ڸq����RQQ!  ��DEEɁL��>�� �Q]]����?�0�����o#��b���  �5DFFʺu���/��$IIIf���	��h�lYYY����Hzz(�9|���w���'  |;v�yޭ���+W�Hss� �!,,L�P�����r�\  |Ghh����r (���[���K �"�KKHH��M��tT��   `��f���� �G�4�g��X����ڵ��ƍ�?��NN�:�� �m�g^}�ի����έ��`�顼y��C���  �!z�RY�;w�L�ʨ��y�}M �"��ںuk��K�/���gϚ�k   ���3gʲe�h`����%&&�`�6	yMMMRXX�h�z�����+� ���֓&M����W��2%Cm���i�&y뭷���V  �o6��RSS�4M ���W�7o�;w�l���ò���7��D�	`q���r��  �����9}�t0�$))�4�������^�6��vQ]RRb����h��[���  067n����KMM�\�rE���
`����Ȇ�׿�5�U  �}��u��K�
 ���J�r��	`A�aI/��rhWW����4��  `diS޺u�L�4��b~֒���� ����Jh��������*]������ �`�M:JHH0�U�ww}}� CA�]�������  ���9����L��p8������m۶5`1�aI���y��X,N�W�  0�RRRd͚5&�`�DFF�����8]� ë��A�9bBK���*�gi~QQ�,X�@  �}v5j��� �ݫ��	 ����6g�����w�}W:;;  x7=T�k:e300P ` F������X �!����Ύp�\�`q��\\\,   93gΔe˖�"���X�A�� �GIǏ�oi/--%7


� ��N	��;L��k�L�b�i����q�Fy뭷���N  �w����{��ҥK ��p���/����?�9c�`)�a9��W\.W� W^^.7n�   ?l�1c� �<m���?ml��ᡍ��!�o�>9v�tuu	��� jAAA���n���_�.W�\��><J*oذA~��_�ٳg  x7ͮ���ɤI�  ��������`!�a)999q.��e,����4�  `�EDDȺu�d̘1����Hbb�����������G�5�j�������
���2߅  5}��iI����9�ҥKf�����`Y�v�y���M� ��>��3��& p���/���n۾}�U,��;��/�W� w��)Ɔ  � ���p;�Ҁg����C#�ё� ��֊��M�H/=<O��z��}͚5 �p�gp=\��� ���&����"�`�gk���k�.���  �>��SY�r%k� "��riv�%,��;,#;;;�}�������  ��5s�LY�l���D�k���p �r:�f<t_��رc���%�6� �����qqq�jjj�+W���;0X�'O6����z��s  ��N:-p��� �������ꫯ��%p�e8=ĜX^II	�j   �HG�k�}ƌ�3bbb̸���h�Y��������BN���;=���: �H�gu����M�AwV||�lڴI�~�m���  ����QKM����p8��g`�a	�7oNv߾-���@]]�   `x���ˣ�>�B,�!������&����3����ĉ���ӧO�M[MϜ9c�N iQQQ2u�Tioo7��ׯ_`�BBBd����g�9|��   錄�.]j�X �6�inn�?n߾�� #��;,!00PO��
`a�����g�	   ��6�=��c4L�����t��� ����eee�����"���x����  K	��'��}Aw}.n�N�Y�x�$''���/���  ��>':t���gB���r��'���c��g{��
`q�y��l   z������Kpp� ���IMM���00p�����v>߸qC�������?/  X��'�;�ݯ^�j.�a ��N����7�|��[  ���~ש�3f� �M/�����w�4�q���?��aq:����\   0�fϞmZE� �k�E[ܾ��F3�Y��vu��5�o9~��tttHHH�  `E���fJSJJ�yV�|�2Aw�6}wܸq����0S  �w9����%( p������A�1�rssǸ��D �;y����
   ����\�t��}����顐��xr!�	�}�?s����K���(g����.9v���� �������{rr2AwHDD�<��3����ٳg  x=�?j�(��� ��������^;/�!���r��Rho�����˕+W   CGø�֭3�� n��0��Z��������4�z<xPZ[[��~6� ��栻>��E��J'�́�  ��>ʃ>h�������}Q�B�#楗^Js?D��Ks�\RRR"   :����K\\� �u����h��l��`/**2�e�TUU	�U:$���w  ;��=<>v�X�~��it������T�y��ITT��޽��F  x���f�}a�.�۴)''�;v�8#� ����ӣ'|���K�.ICC�   `hh�ܣ�>*��vnU@@��3�V�� �Xgg�����^ZZj�����\jkke��� ��h�]������իfR-��ӧO���X��/)mmm  �CEE�)b�.�۠c��^`������`a��{��)<���O���ͥ�!!!��J�I�?W:
��QGR���!���.���0wj�E�
 ��f̘!˗/���l�޹s�d߾}&�~��1�������U�V	  v�Aw����׮]���D	6l� o������	  ����f��Nl�[�!++�'���Z� Ì�P������rߘ�K+++3b�vhp=&&F���%,,L"""�/�{��[ZZ����Vijj���F�  ��@����eΜ9��i�])n�@��4ls��Qh�`{MM� ���-�  o��}��}Aw��U4���s�ɯ~�+�x�   ���?]�X�h%* n���}���F���0�rrr҅/<X���u5�UBCC%>>ތ��K{5�>�44���K�ϱ�L�C�� `$�a��zH&N�( ��6-&''�p;��ﴷ�KII�وӫ��ԴlC�����3�p8  o���έhit�����'�xB>��c3!	  ؟����{�G �=�����۷o/`�;����B{;,��ɓ�t:�Ydd�i��P�^��Vn.m��s�����6a��ׯ��W  ��N4y���%11Q |9mV��N����黹NX��k[;,'=0~��y���  �I_���%莯����˗���O?���3  ���+WL�!##C ���\��tߟ`pǰ����t:�����jkk��իh����i�H�lt���4��W�Ƽ�5�Wee%#i CF7�}�Qr�Ŵ����`;|������jnn`$�琀; �[�t��0;�N�/2{�l�O��;�Hgg�   {+..6S���[�Tvv�y��WO0L�cX9�ο>w�09���]jׅ���4,
o�x�8q�ٴ�����/ʥK���  x̤I�d���^�{���IOO7��_���&'N�0!���|ӖXIAA�<��3 �7Ӡ���kً6��qoo� 7?~�<���_�B���  ؗNe),,�E���V���5��B)�Ac����	�۳XXEE�p>H�2u�^�o������[@@�i���{�1M=�3���  1w�\s��[ l����9444T _��geee��EEE���9rD����� �	Z��䉉�f�X[�Y��t��L�]C   �jmm��Ǐ�|  |���yyy�m۶��1l���,L7�O�f��/	�q�ƙ����i�_������.�Ν���riii  n�6��X�B�O�. ���u�`{xx� �@�Q}��C��n[��萒��={�  �+�ֈ�F�ܯ_�.@}��	7���9�
  �K5��řI- �5��N�f@�`6ưx饗�zzzho���9sF:;;�O�'O�,��ɴ��m�6m�L�:մ������ �J�	�f���� hԨQ&$�Kx���F9|�p��w؝~�	� |Qpp�)������
�t*������KAA�   �:q�)e��k �Oeee����^�+�w���=��_X�6qi;5����jC�w�)111�ۧ�Ǝk���fs(Dnt�  }�`��?n6��^TT�y���������0�hX[�N� �BC[999 ����n]_�q�TTT����,\��|>>��q�\  �G��tMoѢED��W��������� C��;�\^^^��A�y,��ɓf3�GD&M�d�5p�Ѐ�6�i���ӧM؝�; @�=�x�	�7������T3��6���f�K�H[[� �J�}5�G� ���;�]w�e~/^�pAZZZ���l���{�  `S��WTT$��� ��x677�o�o�~A�!D�C��r���,�E555ɕ+W�E�333e���ۇ����5k�L�2�l�kK#�� �����Ms{XX� 󳠍���M����&W_����J _�Mf��e˖	  ��!���[jkkM�{{{���iِ���|�M>  ������ܹs&k _!��ri���B�1������_f/
`a����D����'ʴi����������3U^^n6� �A�>���(���	Biii2f�3�����)..�oi/--��>M� ��F�m���ՙFw}����w�g�yF�x�inn  `?'N�0�)o�5^�����;v\`�pǐr80�e�����j�wHJJ�o|�#�Tz�����ѣG���R  �M���X��2|���������_ ;�C�:��/�~��1��� �s��!  L�j�=66V�]�&�.]bҧ���ƍMȝ�O  ؏\��ŋKPP� ����3͆�
0D�c�����Q��X�>��:uJ`:�r���2v�X�5DGGˢE��fƑ#G���I  �E7�x��7o� �NZ�����[ҦM=������|��� _�/���:  �Ӄ��N��H�;SP� ����M���o�-�ϟ  `/���RTT$s��aR)���[�l���_��K	�2��W\.W� UQQ�xD��f̻�K�L�Bk�E%''��ի�a��'OJoo�  �O�Z�J�N�*�/�1��Ǐ7��]��TIIIK��ӧ��+(( � ��е�q��ɘ1cL�]�����!��{Lv��E�  6��pgϞ�;�C �K���^q�_`pǐx��c���r�(�YZZ*�������LS8�MC�z!##�I
 ����k֬1�^�WEDD���EaN�S����������- F��x�	  _/88X&N�h�PΝ;G���-���  `/�}�����H||� ��زy���ܹ� F�C������[� u������O``�̚5�,��^"##e�ҥ攷�j��	 �^��z������(�/�p����� cYae�����v��SXXh�gXZ �V�!�3fH]]��?��������3{~��9�  ���rɑ#GdѢE" �B������X������E9��\,JN����3z�h�;w�Y�=�B��0�Ѵ���j ؃��p{TT� �FC�����F�� �ikk�'NH~~��4�`h���ʩS�LH  ܞ��8���5S>/\�@	���称�0y�w�o ��h��������/ �Dv^^�?n۶�F "��s:��q�b�(݄���؇����N��I��;hc����H���[ ��4����Khh� �&))I222�$!�*��V'��5��QAAw  HCQ����/_�lgj3(|�N�}�g��7�4u �=���JYY�L�<Y ��������� D���+�����G �jjj2��B�I`]�w��
ӦM���9p��i� XϤI���|�>�7�������:$---`d��᷿�m  �����K��&4ߐ��lB�o��ٷ  �PZZj����> |��������o���Z� B���ё��`Q'O��	�Fe�������� �\�҄ܯ]�&  �9s�,[��	*�)QQQ2~�x���`$566�ѿ�=x�\�~] XÉ'�!=�  G���W:_�pAnܸ!�~qqq��sϙ&���*  ֧Y�$�h�"2 �H����b�	�!��1�7os?��X�.�UWW�a�ԩ&T��J���x���&$PRR" ��7{�l����b���� ���0�,�����%ǎ�oiב�N�S XOoo�9rD|�A  �m���]��驪�����ޒ�/
  �>}F�R��s�R���8�����~�m۶f<��;<&00�O�7� �$=I���>K�/C���ߢ��ӧ���C�IOO�  ��~/X�@�̙#�/�E�1c�HZZ����0�*++��:Ѩ��M �CAAw  ���ѣ%66�L��г,������ׯ�w�yGΜ9#  ���@bii�L�2E �sb�Ng���S<��;<b��́�����
in�p���(R��є�]���%�~�) f�]�l�iL|�'Ə/������:9z�h�]'��'�9  CC�'Ǝ+���f��f驪�׬Y#|����
  �O�O���Hrr� ����/?����$�������\.W� �-ЧO�X��v/^�X���З��˗��{SS�  ��n?��#2i�$������4��Pґ�����-��l�� ؟6��� �����w�q���U^^.7n�x']�Z�r���{��1  ֧E����v �Ibgg����w�֭[�jjj^��Ν;'�_��JJJ���j�ODD��X�B���KC ���@Y�v�i���n�����p����ӜN�i/��k0���K x���BY�n�  ���k�:mN׉/\� ������Z|�^u_   X��{��f=�� �q?����͛�u�Ν��aP�cЪ��u)M��t���ٳ�Ҧ3}������=���~�|��  </88X�qIII��%$$�Cz����Zd���7ϭL |GAAw  �Qbb���ř�b���t$�4g��7�����  �khh�S�N�]w�% p���������%� pǠ�,Jǿ��a]���2w�\N��+�����ˡC�L; �s����'�0�_�[EGGKff�������.%%%�-�O� �I�ur�  ��5n�8v?��	U��̚5˔2�ڵ�<o  �*//7�ur* ���[�n���zwJnn�
��5[ ��� ka� }����	�[���x��ϝ;' �����O>)111x#����ѣG0�(++��=z��� �ؠ�
S�0� ��&ӦM�������)�.S�N5��o������  �.]3�}'�f ��N�������w���(����+�m��p;p;�M�#I�� 0pڤ�����H���Ӧ���43	�����@�^��� _�����;  #(>>ެs\�|�\�~�1a�3}����  �0-9|��,X���C 7��p� pǀ�����r�
`A7nܐ+W��G�F��w� �!w=��W.^�( �ۗ��,�ׯ���P�Mll�9L"��hmm���"���7�v�����?��?  0r4D���.����ͽ��V�=RSSMQ�o�!���  ����AN�8!3f� �O����.޾}�' w�_
`Q�ޮc�a-�9o�<N�bP4�>w�\r�  ��]��c���΀7�����#P�[�ϒgΜ�oh?r�� ���ǥ����.  #K;�y�R__/�Ν����w�g�}V����ݔ\  k�I�ZD��Q ��N���7���������j,HO�^�vM`-��H���������'�|"UUU �z�]�f����)))f���L|me��:tHZZZ KGp;v��  ֠�����z����aV��r׽@  `MZ0j�(��� p8Ksrr�߱c�!n������\.�C :y��Z�IS����<E?O.�?�P ��N�*�V�" ���=��D|<h3��<(ׯ_ 
� ��:v�X���7M�555���&�����TWW  ����),,�|���>��6p�m����r��`A��\[[+����PY�x�	�i����ݻwK{{�  �جY�d�ҥfc���?##C�Ygg�i�ki/++�ї CM�s  �5�;��ɓ͔ٳgϲ������駟�7�xô�  �inn������ ��nٲe�믿Nk-nw�6??��>;� ��E{��ȢE��b#0T"""��L���48 ��fϞm�n��3f�	����>���&X�w�^s��� n���t��W  X�6��0�fO	�"O=�����r��%  ֣�\qqq���& |�#  @[�7	p)�dgg'�o��˗/�S���͛7Obccj�9{��$??_  �s�}��)�7�m'N4w����:9z��	��߿��� ,������C	  �.ݷHII1A�s��ICC����'��_���'  ����b5j�DEE	 ��r��޲e�߼����"�-���-D �ѱ󥥥�6m�Y(�����:u��:uJ ��͙3G.\(���D ����L"�MfD�z�{M� ������;  6j�0jkk��ٳL�1���裏ʯ~�+��  X�>g麮Nd��~ >-��=�g�{� ����eYYY1��f,�������*����d�>}� �m�̙�u��ի �J'�̝;W �=z�dffJPP��w��岲��@��cǤ��K ���;K�p   ���Nm�x�"k�6���'k׮���~[Μ9#  �ZZZZ�:�=��# |���zq˖-?~���ϋ[B�����?��%)���OZ�#<<܄����H�ϝ~���}� �f�����`g!!!2a�����mM���}��Iaa�455	 �M]]�����ĉ  ؇6���j����6��h�}͚5�k�.�� `AW�\���x��� >-������ ���;nI^^^������4ܮc�1�tq�&�����`�^���P �z�G�;�~;�gɔ�IMM5��joo�������ӧO x=�C�  {����Y�fIee�TTT��,�]KX�j��3!w  �����L�����jvv��^}�UZ+��㖸�X6��d,����4j��O�.�������	p�����Ah	!!$!$�6v$bl�1��l��b��	ә;�������oe��q��*ql�v�SI�;Nwgq�鎑Xll��Z@�I�3��&$��Y�t���s���S/�J�r^�}�����n�����
�% ����|�A͟?_@��mk�KNN��:<|������ ������  "������m�Bd�r��}�  ��։m��6%$$@���{}9p�K�A�w�����.��,$q��5�}���*++����:uꔺ�� ��6^W�\�ٳg�D��]PP���!�X��@�>/^�( �vv���l�  �\6��֗{zz��;t#���~�a�J	  �r��e�ݻ��� ����m|����jjj�.�xL__�����Y0�{�qBv�W��Ѿ�o�� ��6�V�Z�L� "�ĉ5}�t���	�����N�΍@{GG�  �X��BT�-  �|��n�l/����B�Q
a�W�w�  ��'N8�YV~ fM���z"p}U�-pǝ�� ��va�-X�@)))�ƾ����sBV Mn4QY�i�	����		 r]�~]MMM�ki����g �����;  �#>>�y��)���n�K�r_�l�sݵk�  �w�������`� �a��������|-[���|B����������䨰�P�W͘1CG��a@԰p��իUVV& ����iڴi�����ɓ�������8Y ��Y������  ��رc5w�\���;��F$�r�&w{�  �`e��μt�R%&&
@L�][[��m�~.�cp�-^��� jll��������Z��Y{�O~�]�vM �,�n�:�$�����6--M����N3�m4��׿Vgg�  �f�-�秵� ��b�2S�NUVV��9��/
����s���n  ���-��٣ŋ@l����M%���E�k���3�Gx̥K�t��	�}��������U^^��{�
 "�m�nذ��LD���|' @k{d�Ѱ���/����fZ	�.Y!�Ν;�r�J �蔒��ٳg���ÙJ!Sd���{�⦷�zK  �l
{KK�
 ����555�}��w�w|�߶��@��<x��B�&�Y�f	����jkk���� ��6�6nܨ���"55�im��D�����z�� �"� @t�6�<g��&���nL%&� �w�۷�y�������'��g�w��׾���k׮��c�ԓ'O
�;w���D
k�]�`��H
 ����=���M�& �3��ɓ5e��#�m�p�᱀;  ���ɚ3g��>��ڪ�ׯ�f�qqq���W�� ���x׮]Z�t� �|r�����sϵ
��ׯ=p#�c��ҤI�D���\����ĉ�H`�s֭[G�#==]EEE�?"Ӽy�M��� ���٩�G�� @�8q�ƍ�#G��ܹs��-\�й���  ������ݻ�x�b�s�����8p���� ��?��/9���?-�cz{{��˂v��D�����ԩS4� �<���~�z͘1C����u�ԩ�xv�#ۘ1cTYY�l&  �g-�� �-�>UQQA�{� � ��Xa�,..������RSS��<��g| w������.�x���PRR���4�ʾ��,{��!�WYX��Gq~^^����|WG�-D���*� 0Lp�ԧ>%  {��=33�	h�={V�.�����  p_cc�����% 1�FCo|��� ��ٴiSB��5s��uuu	�Wii��HW^^���f]�vM �5n_�z�f͚%���ٰ���ٸGt���ֳ�>+ @�점�s��K  {UVV���'��Z�w�s�=��o�-  �.���k�.-]�ԙ� ��nݺ����7�yE�o���ILL����"�cho����h`��3g��� /��|Z�b��
x���:��>��?v�X�?^ �����i����3g�  @�����t��=�����׎;  �u��U'�~��:�f bFv��׿�[��!CCC���xMgg��pw%$$���D@���VSS� ^p#�>{�l^��ӧ���l�Ă�_�B �����p  ��G�%K�8��  ��Ç�Qbϟ����M�3$@���<��2��?W��466
�+--��ѣDkq��}��	 �f���˗���edd������Q]]M� ��@�~�i  �m�---;y��������;  �:t�233���- ����uww����D�����
�S�N���WpW||����D��!s ��6����)��ڼ�N����<ƁƐŋ 0<Ѕ�   ��C�6]�6wo�u��z�ir߻w�  �{�~�v�ޭe˖9�u b�eX	��A�������e� ����f̘���M%�>}���� n���UUU�(--M3g�TRR�[&M��j8y�  ��`Ԟ={�t�R  |Ѝ6�Ç�ܹs�wX�}ŊN����  pO�v�ڥ{��)������ݶmۻB�#����^�y���8qB�ϟ�eyj����XS�-V@��w�}�$ó�L��|hm�]v��?��  ����'�  n���+**t��i���8���7B�ְoSy  �{l�͡C�TZZ* ����=p����C[�n��� ���=��}j��N Z��;??_����p���O|��&99�9����*Ķ��j� 0L;v�  ��L�8Q�ƍs��/\� x��Į^��9x��i  �e�I��������?][[��۶m;!�4�������%E��X���ŋ��hoG,())!� �,4z��
�I�&����Q�p,Z���.�" ��	�'O�T^^�   >Θ1cTYY�<7=z���a�ď<���n�` �{�y�-[�LIII����,���BL#��6mڔ�����!�h���$�/==]����]NN��}�@8,X�@��� /�����b�;V��|4k�,Ʊ�0544h�ƍ  ����L�wsk)�r��>��_�^?�я���,  ����g�eɒ%�� ���o|�������/1��{�KHH�L��/�C�ي�vo(**+
���
 Bi���N��%v�qƌ����QUUU�`����	� �;����y���رcΞ�g!�6�?��ZZZ  ���۫����\ �^�+W>�>'�,��� ��vk���l����@@����{ｧ��!@(TTTh�ʕN�			΁�����8p����- @�]��5i  w��MFF��of��p׍&�����  ��#G�8������~�ֺ���|��(�1�g�Y�!0G���<y��v��<y�ƌ# V���ƿ?~\ 0�fΜ�U�Vn�gdee9��rneΜ9JJJҕ+W ��u�.  �1n�8-X�@���:}�����x=��cz�����!  ��={�h�ҥJII�������������BL"��섋 ���[�O�. �X#w #m�ԩz�Gh�'�F�M-���p'��ܹs���o <kq'�  ��L`��{ss��]�&��ޓ�|�I������  ���A�ڵKK�,a��r>��2��c�USSS���!�tp���}�8�8'ĢI�&9�{!��`�O7n�脊��������)=�kUUU�`������SO	   X&L�رcu���={Vp��ѣ��O�W^��  \��۫������R �����ڹ۶m{W�9�,b����|>���S:$xÔ)S8劘dM8���jkk WVV��ѕ��(�m�|g��{���U]]- ��������Srr�   �e�LeeeNi��c	�HII�'?�I���˺x�  @����(##C�'O�������|A�9�c�֭[3>'�Cho���S�
�UӦM#�`���ӝQ�III�d�b3g�tހ`͘1�9����# @plR؞={t�}�	  `�l�q��˗/hM�W�\  ��{�:�E6�@t���������m۶�b
�488�9pI�!��{��L�8Q@����UBB�> �`�hob!n?~����ϫ?�ǚ�-Z����' �����;  16fΜ9Na�I�7�8���k  �k׮i�Νz����� �R��Аe^�T�)�rǘ�������-<��Ο?/x��{G�% V�����Ǐ eۆVff� ���2�H���'`�p�᫯�  �H�5���B������	x!�lOa�ƍ��~��  ��ڷo�s�@�zzӦM�����b��������$�C>,x���b����-�����+''G�[�����ę$ ����j ����U���</ �gS��ϟ���F'���:u�}�Q��������  �˦��3��ɓ *e&&&����y!fp�1>��V��X{��s�� �p �{֖�n�:���p�ĉ��6�� ���UPP�l  ������   FZbb�*++��7;X��+**��ի��o���  ��޽{5v�X���@�	<c�q��7�G!&p�!�7o��T	������TRR��Xg�6ҕ8 �׮]��7���k�̙γJ��N� ���;  %�ϧ��<���:������*++�իW���\   ��]��]�v����w�N D��g�yf鷾��7���O�2jԨ�<�ԩS�����Z?�Fnn.w �e��+V�PII� 7؁,�[KjUUUz��W ގ;444��  R�\:�|9rD���Bx����˗�g?  ^.\лﾫ�
@��m�;�A�=Flڴ)7pyB��Xs�%;;[ ~c	jll ܊5@̞=[��L��|��Ao�7ւ �����P  ���8��!##C����!;�ϒ%K~�"  ��ĉN�e�ԩu�n޼y�s�=�*D=�1"11�~��J?x��ӧio����,�| ��ŋ;m�@��3�	ť��������k�޽ �����;  �������СCN�8�g�ҥ�����  ��ֱm��M�UFl	\�!D=�1���.�����<���-����߰���/^�( ����
�w�}��$9-ڀ���	��0544�_��   �%99Ys��Q[[�:::��{k֬Q�ZZZ  �Ǧ��$�x@			U�ڲeK����/	Q��������e� ���줽݃&L�  f�w em��V�r6��p���3f�`�\g�+���J ����;N�i���  �Q�F����i1mjjҵkׄг��u�������N�8!  >�.]r
[.\( Qe����\�����ǆgx���dm� >����V�S�L�ڵk��) \���4k�,���p[yy�RSS�� @p���:S1   �m���?�u��!��5����+�����. ��f��_PP  Q�끏52���E�=����,\	�����={V𞌌�0k��l�kÆN�6.6M����C���`���  x� �kUYY�cǎ���]=����O꥗^����  �����w21��Q�x˖-˷o��S!jp�r>�����
����Â7�;V >�\ 7X[�O<�1c������&���'�k,�I� ����^_���  �[{�6m���ӝ��k׮	�e��l���_�իW  �chhH;w��ҥK��*�{�?�I4�g��ax�ec�Q��{۴iSn���c<�ܹs��󨴴4⁛�{9�|�� �.kW��'�����s�f�r�� /Z��Aq 0\MMM:s�Ə/   7effj޼yjll�ŋ�в�?kr��W588(  ��{�n-^�X�3j?{��N�<�|�^~~�.\(�#����?��MBT"��7~�$
��۽��j��٨2�@�5j�֯_���l�`����Ŋ��u�e�&MRGG�  ��Bk{��  �6;l_YY���V�:uJ���\=���я~�4� ��8}�����5c���nj� �Ϭ�ɚ��>���BTb�<J��֎�o������w�H|<� v٘fY��)S�8��^g-����  �khh �  <Ê,�e�/VZu��u!t������O�S ��ٿ���T�߻]����]�Lh� �x�����m۶�u�G����O.9<�n�!ޔ��& 7��c v-Y�D���B-!!A%%%L�AD���&� �T__/   ����ܹsu��A���	�cϽ��ڵk�  @xXv�~�.[�L����Uwj���Ǐ;�Z���< -�}�B�M�:ܣW� ��|��N�8!x���#�Ħ9s�8�M �Ǝ�,��"*"SUU����(u ^WW�Z[[5}�t  xIRR��nii��ӧ��Y�t�s����  �q���޽[���'K>j�W���#G�h����`hh��������M�(C�=
���,\
�{�!��mx�����" ����P˗/j����6m�|>��Hc������ ��Y�;w  �Ev�����������^_�غ��իu��%;vL   <:;;��Ԥ��bE��
��ѣG5s�L�3F����E]]]+�g!�p�N��ac�i�]�pF��x bKnn�֭[�l���,�eff
�d6邀; OCC�>��  ��rrr�}���Fg�#��"7lؠ�}�{���  {������,E�����g8;�h������m��C�=����N�yL�GX������Ӕqqqpsv�}��=������SBB��PIKKӬY�4z�h����J���w ���Pbb�   �ʊ`�Ν�r��F��=��z��u��E �г���]��t�Ҩh"?w�SB�P�GY��5���X��3�|�[�j��(��������ۜkk�w���	ܞ��-99��@b�	Bi�ĉ*,,dB �Ƽy����i
 ��ʕ+ڷo��ϟ/   /��teeeN`���Uyv���'�p��y�  <,`��s�5@+�\�p�y>koo��˗���v�ZZZTZZ*�F��~���!jp�"��]�`�� ���{���pn�Nkۋ!��d���ܞ��! l�5XDۈK�Ξ=[;w�  x���� @����s�؇rʮ0�&L��U����-S� ���ngRMII�"��������EEELȆW|�_�����/�`%�G����G�i<���7D���q� �˚�׮]�I�&	;$e�L@����&� ���Р��  D��c�j�ܹN������Ț<y�֬Y������  ={���̴����K��t�a3g��Y�����/Q��{ta����FkC� ���	�z�!�U �
`m6��Vp�˿�K �w��A'fA1  �HaS�***t��Q�8qBY�f�r��z�- �гCe�w�ֲe˜�"/�j������UXX�~<!p/o���O�(�e˖�˃<`hhHG�"c��۳�z ������4�B~~��M�&��' �;�9z{{ ����ڵ�9|	  Ilݣ��@���jjjr�k0r�P���}�] �����w�h��^��wl��B�����S$�T;�8c��x����{�=B�#�%�T��}� 8v��Ї�' ��}Dkն�)`����fee	��F�҂����L �����p  k	JNNv&�\�zU9��x��E�  �^OO�UZZ��s�~j�rS���a��ӧ;{������l"�(�u�֤����� �C{{d!��/a@t�8q�V�^M�6F����ϔ�������X�   ��zȜ9st��!'���a��֭�+���S�N	  ����Ǐ������;lJ��O�8�K�.)�Y���t�m~���[�n�?���o�"�(000���%S����G�i�XE��=�@�HOO�c�=���#)##Ù�k6b�� ����ᬫM�<Y   �������u��Q'���a�M6lЋ/�8  ���=w�ޭe˖)))i����ϟ�]�=�UV�:m�4rH����F�/!������_��0/�����	�p{jj������ςbZnn��L���Ǐ <kq'�  "���Xs�5�[�ihhH���4=����������A ��PCC��,Y2�B�M���x񢢙�����PSWW���/$��{����Y������ӧO;�Yh�n���|���v�Zegg)v ���XYYYb���p�᱀�O<!  �h`�p���jll�իW�����њ5k��믋<  B���Wt&�܍X
�TSSwxŌ���ן	��{���n�%^a-�<4g ��}D��K�jƌFʘ1cTZZ광�������_ ������ׯ3E  D��8g�:tH�Ν�o�̙�����_�J   �,����I�&��ˡ��b���N�`�6�֊�{D#��6mڔ����vj���G�<w�۳���UYY��
)*))Q|<���,p�<7@�l������+  @�HHHpZO[ZZt��)a�/^��g�j���  ���;�h�رPzt��e'���������N�^�������L}��g�	��������e� ��=rpn���\S�L�ʕ+�k�>}���|XZZ�3�`߾} �����;  �:��b���ӝ=E�܇��vR-P  BkppP�v�Ғ%Kt����^GG�Μ9#�!+H��x�|��Fe�Q��gBD"�����Fuwwo�v"���XDn���L�Ǐ�ƍ5j�(�e�EEE4N �P]]M� ���6��  �Svv����u��A�����5����륗^ҹs�  B���W��/���W�
�g-�g x�Wkkk���m�x�@�#Tww���e� hnn���"�����ָO��3f�=��c=z����5St�$��������� <;(de<w  �h����9s樱�Q.\�g��q'�΁  B�p����{{ֳ	>��&�������
��{��� ���ǅ�e�� ��	Y��hÆ���0\iiiN�=11Q n����	dZ0 ;`�{�n���  �V��b�G�Չ'����u���?��h ��9rD����6��o#3	�G ����6?�r�� hmmյkׄ�E�p{�'@dY�|��L�"`�llvQQ�sh�����k޼y���7 �W__O�  D=�ϧ��gcKK�<�{\�b�����Y   ^��ޮY�f9Sg �-���)~��g���B�=���?
\���Z ��ڄ��%���O��Q]]�8��IL�:U �NUUw ���  ĊI�&)))I��TkfϞ���.���;  ��߯��fgr�2_�c���C�(�#�O<���%p��1B�Q�fj���O��0s�L-Y�D�pX{Xqq�����Y� 0<G�UGG��  �Ni�����{�|P�ϟ�  x��s��M�\�����?۶m�B�=�������S���);D����5���&N��5k�8�d X			*//Wjj� �����.���) @�v�ܩ���   VX������6�ިQ��v�Z�������  �ۮ_���+--ಬ�����kB� �y6	��S�N�ҥKB�&��/pg��������,���c�9�d X)))*++�A.ԏ�c �W__O�  Ĝ�G�QWW�p�lm��J_z�%���	  �mmmm����x��p�WE�=��S#�lٲe���_%�la	��»��ES)ps�/_v�V �&;��n�:~�aXƏ����#�����; SCC�   &���̙3�����V��7N6l�k��洦  �i``@Ǐ������-[��ھ}{��G����W�~� ��H��g�
����	7Ǵ
��V�X���|��4i������`dTWW;�� x�ϟWSS�s   ���9m�v���ؚ�U���o  �m��͚6mep���{*p���G��������/� �ۣ�5T�9����͛�ٳg��o������# #˦":� ���ر��;  �iYYYJJJҁ���/ܝ��rutt��w�  ��,wq��)�#�/��^x��y�#Dww������p�5wvv
х�j��q �d�>���`��ǫ��Tcǎ�Ш��"� �T__�/}�K  �e)))�3g�rg���=��C:s挎?.   7Y�*wx����ԍ��+��p�~����0��F#3f>�\�pA n�����֯_�;e̘1*++Srr� ��ܿ���	 ��{��ʕ+Nk)  @,KLLt&9:t�	k���꣏>��~���x�   ���۫��gJ�M"��G�-[�L��|+��F������"���-ּ�q�F'�ܭq��i֬Y��@h͟?�	  ���A'�x�b  �:j�D�cǎ�F~��Æz�Wt��5  �ŊU	��m~�������m۶<�]������H� ����hhhH�>��`Z����������,_�\�����ĉ5c�1k���О={ ^}}=w  ��:u�3��ȑ#L�����r�J���  pKgg�.\����tn
�K�Q��O#��quuu����_��ׯ���M�N� h�����{�Νc�����R�ݚ>}���� ����	��0�رC[�n   ~/''�	�<x�F�P^^�ӧO�  \��ܬy��	p����ҦM�����?�'xw����^��Ā�l���[oo/w�#Ο?/ ސ���x@�ݰ��%%%?~� �_UU��}�Y �g{zz�  �cǎ՜9st��]�rE�3˖-SWW����  �{)--u,.����1p}Y�,�޷I����
��̙3*,,�߳ �و�68ae�N���;�c��	�7�A@�l��Ν;�z�j  �Ò��~r�IŸ=[c���_|љb  nCCCN�CYY� 7����%��a�=���fj�B��:;;Y�����a���,��~�z%''�S��`�b|o w٦������o
 ���z�   ��+**���Ě���r��588(  �pkkkSqq�����ݷe˖Y۷oo<����n�/��~j*�:;5��g-JLL 9�m���V�X���\w*%%E���<� Q]]M� �iǎN����   ����9s�v?u�p{���Z�r�~��   ��ݱc�4c�.�r��O"��Quuu�����(�e��n�~�Q��ӣI�&	�o��� ���:�K��7n�JKK' �`w ��9s�)�`�  ���a@{^�v���V��l��ӧ�{�n  ���wM�>�9��%���M�6�����FD�ݣ���
�<S�����b�^��o0�p�ԩS���S�:e�i6�%??_yyy:y�  �khh �  p�t���:t�%6w`�ҥ�M����  N}}}���p� e'$$<��H������ಁ�������~�����;Ǝ�u��qZw��


��������P �����볟��   p{YYY�d������ǳ5������_Թs�  N������fu	�{w�����ಶ�6}b�5V���;�@,�z��3@����kÆ�(a�NX�inn� xw �={�8e���  ��Y���ٳ����}���Z��ɾ���  @������ٳ�����߿j˖-��o�N��p���>�K᪡�!���
��F5Zk�ԩSĲS�N1�p��?����c�R%%%?~� xۢE��{��3 �������.\(   ܙ��͙3G�����˗�������+W��?��   ��ȑ#NQ�8��g���)x
wo�� ��8q��8C���� ���g���;w�JKK܎5����)==] ��Z��@��� ^CCw  ��dp�ɽ���i�ǳ����N�ڵK   �b�}}}JNN�?����ښ<�������.�-�e���.�Zs������o/P �+77W>����3f���˝�� "���p�ᩯ��3�<#   ܝ��8�X���I�����{���i����  �h477���R��
����\�U��344�� �����`î\��,��(B Y;	,����>�l4�����lFZ���R]]��|�; �СCΚ]FF�   pwF��L�҄�Ǐ7gO�V���~W�.]  @8;v���)΀[|>�ew	�{?<d�֭IO
pYKK��la��;b�@x�ĐիWkܸqn%33S�f�r6� D�9s�8!;P ��Аv�ޭ�˗   ��:u������T=��#�����<�  �ڵkל�{aa� =�y����{�f`� ��!������|${�˗/�ԩSBl������;�C ���+�@xY�oQQ��[���u�x6"��,�c� �W__O�  `�&M��L�	9�/�?d/^�_���  ���fPv7���|�\��@��C~;� pUkk+9pZ;;;5q�D���\�zU �c��ɺ��{܊}O�M�& ������; ��  0|YYY��������P��{�Gjkk  @����9����<n�m����Gp��������.�ś�G�
0��N��ƾ� �#%%E�>�('�qK�Ґ��/ ���v  ��6����5  0<cǎUee���߯����l������:��   B�����;�6���v�m��\G��#�~�S>{C\d�c4�kc�7o�Ă��A�@�X��6FRSS|���"�Q�������̙3 �����;  ��"�ٳgk߾}Lx��1c��Gѫ�����!  ������*##C�[�~���Z�u�=���.����s�C�[��g��������UXX( �� �d�M�2E��عߒ�gL4��b���E��O��O ���^O>��   02,�m!wkr�|���a6a�Лo�)  �Pknn�������M�6����Opw���^��
pQgg'6�G�!���a/I B�~�X�����8���jܸq������0�ܹ�9���>  �HILLTee�r�x��a,�ɓ'u��a  �RGG�������,�%����WW��_���V��������ۨ+ �e�egk��GY@���L������� ���՜9s  ��c�Sr?x�o�߳5݇~�)M;w�   BehhHmmmξ!���o�^�.#��~:;pyX�������K��X!D�C�	@hY3��u�q��G%$$���B)))ݲ��5m�4=zT ��544p  �Q�F9���l��{�G��ƍ��/:�   B��%%%�3���_��צ��_��q�5�]xA�l�� �E�����܌=4Ξ=[III��իW	Xa��Ci�ĉ>�=�����;@�� O}}���կ
   #�B�3g�tU�O�~o	Z�l�~�ӟ
   T����� .u������Cpw��|�/pQ���;&���w�Z*,�D#ko��9�б�#�%q3���Ns{bb� Ď��*���k o����t�RSS  �����TTT���x�8qB���s窣��y&  ����p��Аe{�g�Cs�K���駟.\H��UǏwN��r��a���9�x@4��G������ҪU�|TZZ��|���@+ �,X��y�`�9 �j�ڵKK�.   B����Y������+V8��===  �.8�������mٲe�����\AR�E���_��9�w���
�����d��c������� 4��{�����ƍ�4�ۘg �'%%E���ڻw�  �khh �  �����M<�o��Ǻu���K/9��   �`Y%�p���w�.!�������Op��r��n���1������#jXc��� t��g���>Ⱦ%%%5j� Į��*� 0L���  @x���8{d������7,l������_  @(�:uJ�/_v�s �|jӦM[���>!�H)����gu�2Q���p��\����f'�D�Ç;�k �QVV�|����Vqq��t��f����  xǏ�ɓ'���'   ��7�D2+Ϲ~�� g��رcb  !a�=ʾ3ܔ�.p}U;���� ]�z�9�܍}��9-�6v�d���N�
��7n��/_.��&M��<G ����Pjj�.]�$ @��q�F   <l���im�M��������C]]]  immmΡ���8n��|��%���.غuk����.jmme|�Z��zm�@$;t�s���5j�֮]�ѣG�aڴi�<y� �[��?��z�- �G�   ����TYY�CY�N����wք_|�E�>  ������vg�p��-[�L޾}{�V�]������G��rF��8p��Ӿ���$ Y��Ƈ�%K�8M����� |TUUw &��Z�4  @����h���N��
�b]VV��.]�����  i---��Q>��3���'�w�vd��'N�\��������	� ���wߥA2/Z�H�ӧOW^^� �f��� �.���Qeee  @xY���mߌ�Wi�ܹjkkӑ#G  0�l����9T���"�v�ì���thhh� ���
���f)33S@$9{�,?�INN֚5k�0� c_h�p+ֶ������N �W__O�  �%�G�Vee%!��Z�z����8!4  ��dY�pQqmm�m۶��{�}Q��Ν;���^�����g�-_�\@$ٽ{���0�,�n6�0���)���� ���AO=��   ��[���}���קX6f�=��#z��,!  ����ѡ˗/�'����/.�È�{=��q�˧���b�kY�1�"AKK����`�-X��	4����id�;Q]]M� ����s�T6U	   �HLLTEE!��ɓ';��o���   F��=z�I�pM�;��/~���/0�)L��QNNΊ��<_�K���.`�Xvnn��� x��}�w`�Y���`fΜ���l����Q�F�� �088���{�  �{,�^YY�ܭ]4��s�=:v�N�<)  ��b�Y�f9�
�2RSS��'��0������%Oh #���_{��q� /۵k��}0��裏�� �-&eee	 �Ƹq�4c�555	 ���z�   `k�r߿�.^��Xek��֭ӷ��m��  `$X��'4e�.�����0ٴi�X�ϷN�Kn�iFZ[[��M����<^���ᴄ y+V�Pff������Ǐ/ ���p��ihh   �!>>^N�{,����Ҵr�J����  )������߿r˖-�o�~Z9�a����D�2F�K:;;c~Bg�ΝZ�z�F�-�K���Z� ������������t 0,UUUz�� ^KK������#   �/..�	�[����l�Bh�  	���:w�3!pA����T�����#�>��"��Jvx,Y"�K��E__� �,[,X�j��l̰��322 �1�|%&&:�E ��w�k�
   �p#�~��'���/_�L�=s�   FB[[��Ν+�%�&����駟�\H}�5�`lN@(?~�i+,,����:v� �,5[h���;eee4# n�={�v��% @�|��;  ���XG;x��6��n�:gz۵k�  0\����3��/ .XP[[[�m۶�BHp��K���"�%vjmhhH@�Y e	JOOঋ/j���0�lZǤI���e�r���;v� `�TWWp�a�������   ���$���F�={V���mm��7�  �p]�~�)�1c� 7���O.��R�����}F�KlS��ѣ��Z~��_kŊ��E��=�կ~EӦMӢE���e��-��a6 #��۶m  xgΜq��	   �b!�Y�f�СC�s[,Z�`�3y�&B  ��p�[�~����fB��{�mٲeN�R!�%�O�֕+W��-�����{��k���1�@(�=Z�W��2����;����4�H�9s�ƍ�s��	 �;vp  ���{zzklm�֘���o����  �K�.���K���\0��g��ķ���_!C�=�>+�EvZ7�����pRaw��a�?�Y�j��f����
���
 B�6�.\����g ���A����   o��wII�����ݭX����5k������I�   �a�$�pK�yֲ��C��{��Ս
��~J�K�����j��E������-�ٳG F^ii�����4�njUUU�`�콸��ߙ�   o���M23�r/((Ђ��D  ��8}���\����$.�dmm��m۶�!A�=�Μ9�,p����G�r���~���z�-��7%%E@(��)��	�ȲP���˅�d��eee���ŋ 0<z���h�"  ��b=�~���;{ٱ��  �ˈX���.�|W��!A�=�_��
p��?v� 7�)�7�|S+W�Tbb��P���_��z�����ޝ@Gu�����v� �B,HhGb3H�ƀ���,��M��9�O�C��čk;��(MR7O�ڮ����cgm�ٗ6�0�j�Y	I� 	�u��m��u�B�3s��uΜ��s�8��{������M�իW+%%E��[s{ff� �yyy�2e��?. ��mܸ��;  @��[iԙ3g�'65��oֳ�>Ky  �*���i䶷	D�e�	���#��n��DHcc#aOD�s��9��+V��f��=�����ٳ0��Ν���B����	�p[MMw �Jp���>&   D?�������_�]�=77י���+�  `�,��Рɓ'��[>�Od=��#�F ��������4"�F�Ѣ����\]�p���
��ꫯ��ɓ0�����1���M���,��jkk���}O ��{�7�p�رc  ��ge��o�>����Ol�����Ny  �P9r��;"%�������°#�>r����p�ZZZD[�JLLԼy���[�r�!��b�ax\�#�L# R�y���O Cg�7oެU�V	   ����+**�g�g:�_��E?������  �P�:uJ�ϟ��ѣ�-
YV��� �2֮]��=@�X��6��hcbr�5k����}�v�߿_ FƢE����'�OYY��� �����} ���$=�   ����3f��]���#�.]�_���  ��G����J@\{�wNy�'�Ê������p H�rg_�@��E9k�:`(v�ޭ�{�
�Ș0a�jkk�)--UNN�  �jjj��U���~'   Ğ����X�_\s�5:x�;&  �������J�~
pY��]ܟ����0�����+ B���% ��رùrǕ���Ν;`dؔ�[n���~�p���� ��Z=�$��j477;S�N�*   Ė��������@@�y�{��SO���S   W���['N�Д)S�-
���;����;�~��!G�,���ӣٳg�l��\ #���رc)..&� �TWW+55U ���p  �M��������222�|�r���?  �PX�wDH�w�Q�nݺ]°!�>���G�" lq�ԩSb�޽{����y�f�R�l٢����ȱ�ˬY�)**҄	 ��&�̙3G��_�% ��mܸQ�'"   Ħ��'�k�.����ҡC���o  �JYn����=z� �����b,�aD�}����9|���Xs�����������]0t�N�����|��6��O�8Q �����; \��[�����	F   6�!p}[���ŋ�믿^Ǐ��  �PX��M��
���A��0,X�F6b |��������Z�t����k������  #kժUJOO���	��fp \�޽[�g�   b��YH�/!���4�x���~   �+e�l
%����;fݺu�aA�}�?�X@�466���K@�:y�~����s��o�	����F���0�***TVV&�GAA��L�" �f6ebܸq�8Q ��mܸ��;  ���w�ܩ��Ny]qq�L۳g�   �Dww�N�8�~(""X����0!�>�n!G��Ξ=�����Z�l���������/�6�H��v�
������|@�N������ 0t����l�   �����ʕ+��s��	  �J���[��@�÷�z�'�����	W���0�뮻lv�t`!���f^`���}޼y�>��U�9|��^{�5���
�Ȳ��M7ݤ������4u�T@� � Wo߾}N (33S   �}��ɪ��r�ܭ����u��������P($  ��eŊmmm����	999K���W�����cb��<��K�����vpc���JH�����g�y�f<xP �a� ӦM�!����"@,Y�`�s ��] �`0��[�j���  �7XiɌ3�&w�h�ܹڲe�   �đ#G��7����e�	��à��.����V`�ǎ�E��}��y-Y�Diii�7٩ٗ_~YgΜ w���p�cǪ���	�@,���Vaa�:$ ��Y� ��   �b�fr߽{�S"�e�^{�P;}��   .���ǝ����8.����nm���K. �>N�:e#&	� �r��^e���i޼yN��b(l����G ܳj�*g�+����n�jjj��Uz��W   ﱵ���
�ٳ����l���ի���ϋ)o  �ruww���^���\6���ee��c�pᇨ?!o��� ���mƞ8qB���'��� �y�f�q��*++5}�t���[�h% �,�a� �����YS�4��   ����r
.���'/�{ٹs�j˖-  �\V�H�b�b�W���U���Khii������Ucc� ��O?X[[�	&��>�������F��뮻N𾔔'�n�F ˮ��%%%9$ Cg����   ����VII�8 /[�t�<��g�
  �r�:uJ���JOO���s�=�~���v�J���×�"�رc����'v���_�R�7o��Cl�P������o
@d�Z��i���Y���ڹ@���Yv`g۶m w   o���u��:$�JLL��ի��/*
	  �rX����B��2zzzn
_�/��~p����6k����SS��̙���B!��(�M�6���C "c���*--��۫�����, �
��D� ��k���`0���8  ��&N��?~\^�����ڵK   ���E���
�
��Xܯ
��p�m�Ym��D���������ԫ���Çk�ܹ3f�]Ν;焑,� r����o�->>���IMM xIMM��x�	 ����M���s�b   ���N��4�744ȫ�/_�#G�8��   ��l�hN�0A��޳f͚���ן����UHMM��"�����'O�'?�����4s�L������եݻw���NC��Z�b�����&���J��� ��>�F��� �ƍ	�  ���Y�݂\^d�+W�Z��}�{  �o��wDBJbb�{���!!�~���D��E�����g/�|�M;v�٬-))q�l���^'Ծg�g&��+,,t��𶲲2efr��7�!������F �����_��_   �W\\��Ӵ��ʋ,�ok����  �`���5�A9�M��p"�Ct���]�x�f`#����nH�nݪ�{�:[����]`:䴶wtt@t��o�Q�6;ԕ��- ���Z� p�v�ܩ.0�	  ���***�}�ND��t��q�  ` �i9z����
�)
�p�]we��_=-\1�Ct���[�v66��:;;�c�<x�it�ck~���G�qHY@��u�]�������-77W �u555 \{�߶m��,Y"   x���ٮ]����.�5j��/_��^zI   �!��I�>~}S�b܇�D�5#�:uJ .�-��n�ۍjii)#���M�8|�����Gc;�


T]]-x���'M�$ ����|�3�ĉ ���p  ��rl!w��s��Ey����߿_o���   b�!�܍7N��>$�CB�}��޴���*`��B�� \kt��
dO�>�	��j|������o8������u�7:ch�M'Nt �'���׿�˿ 0tp  ���zqUU�r�����p�:v�'��  ���wD��5k֌[�~=��W���\�x��%U��,�n� ��B���`��cǪ��XӦMSB_��b#�������'O
@�[�l����o���Qaa� �ojkk	��U:r䈚�����+   ��M7�or�Z�Qzz��&����L   �)�6� .J��{o���pEH�͇D@KK�:::`x�9sF�6mҎ;���������f���z�->|X����L��ٳg�4z�h���������=..N�`P ���������  �����:!w�x�g�3g���_�,  �����A��n�+F��
�Y�ƚ�o<�#�F������9����|�?^~s��Y������ ��4�իW~�(ۀ���t �G����!�o �ƍ	�  �TFF���˵w�^y������SO=���  \�ѣG	�#V�s�=c~��3�e#�~����	p���khh��u�?��m�oҤI�8q�v����g��&��{jb�5f��{����v%/~�����%� W������I   ;v��O����K����d���׿  �����������l�E�===�_�Y�l�#�ܭ"�ĉΘ w���999���s����1�lاO�VKK�����g��ƍSMM��=���N�=99Y �wp�� :��v�����	   �d�]6������k��ƹ׭��  ��X�{UU� 7�B����!�~֬Y���ǎ�ȱ�s���X��.,�n�Rk����h�1R{{��q}��)'�n�v�����U�V�Fo���ii� 3k�,���m� �nӦM�  |n�ԩ���v&�zE�Z��g?  \�����dn���{�����.�+���ts("Y�utt8�T ����~n�~z����1c�QF�����B���{/��hA�.8��6J�B����	��fΜ�ɓ'�SRR�|�  ���WϞ=[7n `��s����   �o����>Skk����髯�*  �w����D���
pQb�������p��P�V`�ᬉ@t�0�5����tOIIqZ'�e�x�wv*�Z%���zzz����`�������J{�Ͷ-8Z��� �5j��.]*xϴi�XT�wa�����l߾�Y[�5
   ���M��]�v9eJ^�p�B�߿_g�P�	  ��ѣGً����ߖA&�~��_�5k֤�/7	��cǎ	@l��5��p[�b�r������� �P[[�G}T ���C�r_�`�   �o��񪬬�Ν;�C�^`�M+W��w��  ����Fg�̊*��B���1�֭���D��2%$$X�=M���T��N� ��3e�UTT�2v�X	 ��JJJ����ӧO 0t�6m"�   ��f̘�;v8���&d���9M�   �u��	�pQb\\�{���Ap�|6  ������otF��;222����\���3r޼y��O* ��mܸQ   @?�j!�]�v9�//�	�G�QWW�   ��ry�����e!�~��Q���7p�-444  ��.\�4}�;RRR�F���8 VSSC� �қo��S�Niܸq   �pX���}�����Z�x�~��_	  ��Z[[u��y�=Z��nX�fM�����	"�~���V�t.kllTww�   �΂��w$$$8�H6
 0���Z �N(�k����n�I   @���lM�>]�̝;�	���;  �;?~\���\����tK��-a@�/C �U@;vL   o�7�7ܠ��x����Ml0 �����j�ԩz뭷 �M�6p  ��������N���+����?��s�u  ���|�Mٶ{�-�P�2��A�}��v[J�r� �uuu���I   oWUU����;l�/c� ���4� pu6n��4���  �w�6m�3m���Y�n	�5k��m�&  ���C}v�c�:��n��?�����z�M�$�HMM�>|��2;o�K   �����k������� �rp����- �е������***   �N�~i�l�ΝS�[�t�8���v  ����p��RRSSm�&] �>�@ �`_�   o�b�
;�)x��ɓ��  ��̛7O			��� `�6m�D�   �*..N���ڱc�:::˒��u�u�饗^  ��544���G����-�L�} �p뭷Ƈ/�p����u��Y  ����WEE����>u�T �.--��d߹s�  C�q�F}�#   �n���5c�m߾�	~�2[c߻w�3�  �_0T}}��M�&�-�@���n�-�駟������,_�	p��  ��laժU��#ľ��t������aP[[K� ��֭[��ݭ��$   ����-�n�� �e+W��SO=�D8  �??~��;ܖ>jԨ��� ���,
p  ����Ǝ+�>Y۰�� \���}��_ `�.^���_~Y+V�   p)V�QRR����+��3�YOx�W  ����Ӻp�3=p��3��/����Y�������Y]]]  0l_�`��,�n#pi���SUU�,6ۢ3 `���/���\'N   p)999�����6[s���u��  ����Wii� �������~1^�]p��;���%_��l�	  @��˗+>>^�}�n���! ���ȹs�귿��  Cw��9=��z��'���(   �R


�)@---�U���j�*���΄u   c����e٧N�Z����p���W�����Scc�   Lqq������7u�T�� 0�l�8w �z{���c�=�����   0+����T[[�bU~~�3�h߾}  0���jmm՘1c�%
YV�?������p��,���˴	  �QOHp���Ə�)S� 02jkk �?��f͚ų   ���J�ر�	��*��=|�pL�7  ��U__O�n�?��'�/F��wq�]w��/e\f_�   f������b��ѣ�&~ �ș6m�rss���$ ��	�B���?�b�4i�   �KILLTEE�v���L*�EiiiZ�d�~�_  �X~��ف>�%���?��� ���>$�e===l�  GFFm�����l�� #���F?�� �zmmm��'?�g�yF���   .��eeeڻw�b�M0��~ss�   l���L�0A�[B�����@���}@����W0  ��+��Į��x'��� �a�O���9p�����Q��ԧ   d�ر*,,��Ç������׆��F   ��#��Y)�������;�~��6wu� ��#  @AA�JKK��f�vk/ ���� � 0����諸�Z7�|�   ��L�4I/^Tcc�b��ɓURR�7�xC   ���UB�Z�����.{�������w����`��"mr��i  ��koGl�>}���� pOvv�����o
 0|z�!���;��   �@������ٳg�lm�Z�{zz  �����	����pK(�?���
@���� �?~��9  �9s�(''G�]�T���' ��jkk	��0������߯�{N)))   .�&��d�;v8���&##C����+��"  ���z�p�e�	�����뮻�×�\f_�  ����Ҵx1���l̘1�6m�  �QSS�0 ��СC����/}�K   ���Jm߾]����5vx~Ϟ=:w�  ��577������i��?���G}��� ��6�@ཡP��Mશ����  �ϵ�^���d!6����r�� 6	%))I��� ����'N�����>   ��5��޽;榘'$$hٲe���7  ���'N���H�K����_�Ip�~�����p����  �-//O3f�b�mz؆�� "�6�gΜ�͛7 0�z�!������L   �@233U\\�(����m���  :v�w��2�������s�=������2;�  ������z��c�mx0� �CMMw !6!�������?���t   ���Յbr?|�ʕz�g  ���ٳjkkSFF� �,��;Ƭ[��U �ޯ�����\��ڪ��v  ����v��
5f� �Cmm��q F��X~�_З��e   ��6m�:::�}�X2~�xgJ����  ����^���\��:|� p�
�n�2�  �e��K�.bSNN�&M�$ @���YYYN�
 `d���М9s��X   �@lr�=�[P���S������߯�/
  ��>p��~�e&�.�������pQ����;  >�x�b��2D(������D ���k��F���/ 9����l��D*   ` 			���Ў;+������'  �.8�:V��du]]]R��-�#����4?..n� �����)u  0|ƍ�ٳg��C�B� ��S[[K� FXoo�x�������   0+�&�}��)�̚5�	���>  �/+�%�e��?������p���u� ��8qB  ��n���1����� �Np ���'O�s���y�   �����ɓcjʹ��X�B/���  �Y�oƌ�
�,�L�]������@p��^#� ����jʔ)B�),,�� ��ĉcn� b��/��g�}V��G   f�ԩ�p�Z[[+


�5�7�xC  ��:::t��i����@ �����9���뮂P(����ڍzzz  ��_�-[&Ğ���kҤI D���� ���\��՚={�   ���䟲�2m߾]�����]w�:���^  �=�pQ���>�k_������vҁ�v���v  �k�ܹ���bKzz���� ��������/ ������}�ݧ_|�M>   *!!A���ڱc�s/l����W  ���~UUUN��������/��,
�"�E��n�  �RRR�`�!�$&&�����
 �!���w>����  #�F4?���Z�n��   Tjj�JKK�o�>�
;L�g��;wN  ����t��)g�7���g��V>����5k2×%\�����2  |jѢE5j�[��˕��, @����p'��3 ��7o�7����_��   �����)S������<�t�R���K  �d-���@ 0��;���O��M�����M�K� �  🬬,͙3G�-EEE��Y @�����]p���fr   .KAA������ڪX`e([�lQcc�  ��X�o�̙L0�[���{��oʧ|p��
�����O'O��@  ��|�rtcLnn�&N�( @l����O>) �{���>���jÆ�Y  `P�@@eeeھ}�:;;���.[�L/���  ��������Iyyy\r���Ϛ5kC�Ѝ\d_p���  �bcV����ؑ����ӧ ��E%55U ��̙3�����o~Ӧ�
   ��3VVVjǎNa\����w&:tH  ��ŝ�;\t��5kRׯ_���.߮.'&&._�pQ}}�  ��X��u�]'Ď�***h��g��g��+��" ��v�ڥu��i�ڵ   c�KKK�o�>�[�?r�3�  �Kcc�SpK�\2*�gmE���|ȷ�B��-6�b�ͭ�  ���9�[��˕��$ @쫩�!� ���Okƌ�  �e���v��?~\���kUU�v��)  �/n��I��!..�p��@ p� �<y���  �a���.]*Ď��Beff
 ���� DF(��?�y�����  ��RPP���v���*�-Y�D�������  ��ĉ�w�M�	���;$��e�}�ڵ�`�P���  �˼y�4z�h!6�;�� 𘢢"�7N�N� �}�ϟ�<�'�|�)I   T PYY��o߮��NE���4g��q  �Oѭ�#-
��q�s֭[�U>�˿a��M\����&  �a��555BlHIIq6N  �b����׏�c "c�޽z��G����   cA1[�ݹs�3(�ٚÎ;t��  ��,`ss�&N�(�qqq7�/����;��j  ���ŋ���,D??���+>>^  �g� �^x�͘1C�W�   0����СC�f6�hѢE���.  �/�����&�<��|�w��k׎����ĉ  �������j!6+==]  o���u3E{� xݗ��%�`�ԩS   �cmmmN;j4�9s��mۦS�N	  �G�M�\0���o���}-�o�����v�B��×$.��$MMM  ��b�
%D������
 �]�Y?m�4>|X ������}�ݧg�}V)))   3}�t���;��������Z}���  ���L�I�� .>>~U���|ď������  ����'D�藚���� ��Z�	�@�<xP_��W���|F   �`���)@;v�pBd�ʂ��7p��Q  �hhh �7Y�����¯����^  ��������7Fh� ���ц �����9s�n��   ��������f����s�Y�  �?X�³�g������/ߴ-�*�~�]w�_&
p�5�777  �Ì3���#D?kn�� �?̙3G			LX�(�w�w���PQQ�   ���?^�ΝsBd�*//Oeeez���  ������4q"�T�bLsssm��_�	_�C��́@@�[���s  ��Bs�/��-0�7N  �HKKSUU��o�. @�]�xQ��{����o9��   �`�pd{{��V��~����  �É'��5�@�&p�������^  �fϞ���!��Ϩ��P  ����%� Q��ѣ�����zH   �`���T^^�<�Gk�\ff�3En���  �`f�p[||� �~=(��M���{����=O�K�G�   �KJJ҂��f-�6"��N �O555Z�n�  ��g?�����}��   0������h߾}�V.��ݻ���)  �}�AZ�������>��1��o�===���1�ƾ�= �?̟?_�F�����m �O3f���ѣu��y �����߫��ҹ_   ����I�&�ĉ�F�m�8���o  ������;\���wc��^>���{�M\d�G  ��Y�}�<E���|�3F  ��Q�s��e� �Lww���>mذA���   3m�4���E�!v[زe�� ��YN0:��H�B��&����zk|��z� �������Q  ��l�hRR�������;  555� 
����3���~�a   �{���rm۶M===�6���Z�h�~�ӟ
  x�ݏ477k	\���nKy��;�q�����ֆB�l.iii��i  0��]p֬YB���eee�d  � ��o�[�����G>"   `0�k��w�V4����k���3g�  x_CCw�%-55ui��sy�/�\c_X  ���,Y��_�R�,��HLL  ���@'N� ��#�<���
  ��O�<v옢M\\�3�G?��  ��566*:� �,M��#��5�P��r  |`�ر�1c��lc#33S  ���������� D���^}�S�r��-�   �ց�����ڪhc�77m��L�  �����Ln7n���n	_>!��|����
�f
p�=8wuu	  x�ҥK9}�F��ll  �N���� �555鳟��}�Q��   0�@ ���m۶M===�&��-Z�:  >a����}�c���O���<����U�W@�Kho ��&L��,�#:%$$�����<  ��jjj����
 D�W^yE�����?��?   0���$���jϞ=�6��������F  o;qK������ײ��cY0\E�n��  ���k	OG��ӧ+99Y  ����Lgsy��� D�u��iƌ��$   `0cƌѤI��`Y4���ŋ����  ��uvv���չ/FZ�>���qy���uuuq---������joo  �)S�h�ԩBt�&��� 0Kp��f�6>��hÆ��  �L�6�ٳokkS4),,t��?.  �mV�K�.Y�v����{�K����ӧ�	_X��k  �mٲeBtJMMu6
  Lmm��y� ���ӧ��OZ_���'   ` ֖^ZZ��۷���O�dɒ%��M  �m6M���B��B�Ђ��?�Q���XV���  x[qq�&N�(D��/++#� �,�g�Vrr���<[j ��e�}��_�w�!   `0�F�RQQ�8�h�?����  ���vg�LFF� ���V	pIGG�Ν;'  �M�^�x��l�"--M  \���$͚5K�6m  �=�䓚9s�.\(   `0���jmmUKK���ҥKu��Q�B!  ﲒ\�*��`0h�Oɣ<p_�v���o� �466
  x��?~�}������'  �Dmm-w ��`P�����a���  pYl"���vvv*Zؽ���<xP  ��,GH�n�֬Y��~�zO�W=p�+D.��W  �����ho�R��k  \��� b�Mϼ����6��D��  0���x���iǎ�&��~��!Z� �0�$��ѡ��T#,���dY�oɃ<p[%�%]]]:}��  �7UWW+++K�>�AA� 0֞2f�g� ��٣�\��s�   ��dddh�ԩz뭷-rrr�5����  x�����`��A�Jp�1�p�}!q�  o�����Z!����+33S  E мy����\ ���o}K3g�����   f���:{���K�,с,�$  �M��@ ����..���ͥ'�w�uWI�R(�%��  ����	QG�ѣG;w  ��b#� �ŊF>���;���&M   0;�n��[�nUoo���رcUYY�ݻw  x��ӧ��ݭ��$#,'��mf��]�ɀ��H�Mn�����  �����!�$$$����٘  �j0� bS[[�>��O�g�Qrr�   ��X��B�{��U�X�h��~hq ��,���Ԥ)S�i}}}�D�=f������+--M�A!  �UUU��������	�  �ń	TPP��G�
 [8��~X<��   ��Xkz^^�lr�̙3�}��rH  ����V
���<�s��������k���W�\������	�_�x�]��� @l�����6 rrr �p�i-� 6}�;�Quu�n��&   �),,t
�.\��h�p�B�޽ۙ  ����ٙ�b�`�-Z�v���{�<�s�S�N-_�D�5��k̘1����������-�nW�g�5�  Dko�D�Q�F9  '�[@ ���o�V���6m�   ��X����T;v�p��#-==�9��m�6  �`KK�rss��ľ�>+I⹀{�!dU ��9--�y]JOO���������� ��g�ٵ��Bt��N� ����󕐐��s �Q�~z�����g�UJJ�   ���^��<xP���"�%p  ��ɓ'	���@`��G�������������K�����л�-���<�  \�3f�}����+##C  7�خ��Ю]� �MN����/}�K   ������V�>}:�o�Y����;w�  ���F͜9S�<���T����xnooo� �������e�noo�� ��w���acZ-� �H���!� 1�'?��3��}�{�   ��������z�Y���ݻ)� �����ܹs���0¦�q���֭;,��T����oE��s�-�j��]�C��^6���!x��P($  �����bJKKmR�  )����o|C ����C9�eee   b{�r߷o_�ߊ�'a�����#  �=��N�n��&��B��
T||��-�v2�N��3���� �U����ǴiӔ��*  FRuu��lϿ ����ݭx@�?���0   ������ǫ��9�o�ٛػw/Et  x�ɓ')d�[,C�F'O�Ö�U�p�@xcAw���, ��:{��  �E���3f��g1q�D 0�� ��9s���/ ێ;�����ї��e   ��>}�Ν;��������4����  xKkk���KII0���ʺ����+(�L��c�Xq__�Tp�}���!���C���?  ����蒐���� �-555��#~�_h�ܹ��?�#   �C�,ߵkW�ߊ-Z�7�x�w  <���љ^��������u�<�3�`0�B "�� �E��>v�X!:XkNrr�  p� �[��8�����   $33ә&�����1n�8gm��7�  ��p�e�	�G�P(D��� ����蒓��  pSaa�rss���$ @�����<�^x�	,   ���ٳg#��m-���  �iiiq֫l�90�,K�� O�m���� ,��� � �A��G���$�� �H�?�^z�% ���ɓ���>�GyD�@@   ��XNii��o���a��-l��a  ��jnnv�� #)\�v����{�K1������ᇍqq/^  ���.\(D���bN� "�����; x��/���{N��*   ` ������ױc�"�>,X@�  �2�pAj0�	_���H||�
�3��  �X{��1c����ˣI Qp��_֙ �[{�1UUUi���   b���V���E�=L�<9*��  `x555	p�
p�+ *D�A �+e6�!�RRR���  DRvv����t��A ����O��w�^|�E�   ��7())����#�>l�,w  ����SgϞUVV���2���b>�^WW���ҲH "��.^�(  bEqq�ƍ'D^YY�Mf  �V[[K� <����z���n�:���	   ����TM�:U���{(((p�����  ��Z�	���׮];���;������E�@ M "����  �����`�V322 @4���o}�[ x��͛��o~Sk֬   0��'�̙3N�j��!��}�{  �q��I���
a	�`pi��#Ű������`��� @,�P�-P#���ӝ�  �b�ܹJJJRww�  ޳~�zUUUi��   .%8᳭[����7"�Hyyyjll  ����Vuuu)99Y��l5�H
?T��������6 +���տA`W  �EJJ�����e� �'곟��6lؠ���   �; _XX�D�=�����  �`���͚2e����luL�׬Y�����koowN� ,�0u�T!��g���*  �MMMw �0�D�����_�����   \Jnn�s�x�ԩ���ӧOWNN�ZZZ  ������;F\(�\�fM����cvPL��I��Bx��� ���NkxdeddhҤI  Y���_��  ޵m�6=��Z�v�   ���ܹs���q����kq��(  �p�&w2a��������Q�_! w��E���p Ą��,���
�c����<� �VEE�233��k �w=��Ӫ��Ҳe�   \JRR�Ӥ���G���=��8{��  @쳌]kk�Ǝ+`$�Xp���q��n"qb �+e��qqqB�ظ���4 ��^�k�ѯ~�+ �˚��������3a
   7n����u��i�o[��;w.�  x�ɓ'	��1]"���o�}|�R! ������w @��P��3�ȱ�A~~�  �v���l��?^��ԧ��O*11Q   ��X��M{���n�9s�^}�Ug�:  �}MMM�4Y`���}�����#�A1p���_� ���ݚ�� �hgM�		1{�	%%%6K  D;� ��={���Gս��+   �R���TXX���{�a�Y�f�w���  @�;{��:;;���"`�-���)\��9p7vJ���O  D���d͞=[��)S�(==]  Ă�� �cÆN`h�ʕ   .%77W---jmmu���;w�6o��y  0��Ž��@�H
�B׆/��������	@Duww;��_ �,�n!wDƨQ����/  bEcc�  �RWW��ӧk�ԩ   .�����c�΃�ﻏg����>���t l��C�?\���*Rq�I�I%2(LYA2�P\8�0"�!�0O\N=U~lClS�8���f��=��C�=��1�̷�*��s���{����j�;�#Vst�������W_�� .%%E����7�  �~�a��%.�ʀ�7ܐ�4��:���?p 8YLL�\q�����^�W  p� }������o�'�|�	�   X�+�������޽{����Z
)  ��tU�L�x<X���o�>|���2�����^xa��H?\���.�7w ������&������  ܄�; D���N��7�!w�u�    �)**2Bi�>nvv����ǭ  ��dddDrss����&�!�n���� ������]�o�� ���5\M���F�  n���/ �����P�������   X�6�����k��vɸ�t̃�;  �ahh��;,8v����2��\# ������7�  ���YYY���߿N2  �MtŲ��I D�����[��   �J������B���l}ܲ�2)..fr>  @�z
����V\�u�n�!?�i a���(sss�|�w �S}�c��.њ��!  �� ���ٻw�|��ߗ��   VRRR"��öO�����G  �mll���%$$`��o���������.�{������ѓ����]x �	������P`?=��?  nD� �����k_��|��_   `%��X��7���G�ЭTWW'���F(  ��?�d���R���z�	l�[���]�' ������A���  8�6� <��zLL�  �FgΜ  �O�Sٵk�|���   `%�⏆�z{{m{L��k�>��  �mpp��;,��x~?�yB\�u��/�6�4��a���y �irss���B`?m����  ܊�; �b���lݺU   XIyy��������m����"/���1�  �khhH ����k�e\p����- l.ooW� N��%��c���8���  ܌�; �bz����o�cǎIjj�    ��F���zy���m{L��c�y��  ����LLLHzz� *��[jy���%\p����_�)% L|>ߊ3�	� �&99�h׃����$6�U�  |D�  p���>����`25   V���&%%%r��i�S�/���GVa  �-��a5��M`C��
�_��s����)}~��� N�m�6B�a���%999 ���� X���?/Ǐ�?��?   `%���222b4��A���mm�  ����Z�����qq	W�~<ϵ l4��  '�e@������1�� p���9  V��C+���j   �r:FQ__/o���m��{�ny�7V,�  �p��YYZZ2���*�횀��={��- ,V�eN� �$4HIIث��B  ����g@ ����E��W�b4�gff
   p���)((0�X��j�ɓ'  ����3B�zX���[n�y�G�pM�=>>��.�Z{���;  Nq�W�
��� �Hp�� `-T:p�����   �媪�dddĘ i�]�vp ����wX����~`C��L~���@�LNN��u�xB�; �)���8����Z�x< @$ � ؈^xA�����_��_   p���8#����a�㕖�JQQ�5  p���alpu�����k�܁0���]uf�~��  N�%��6����  ���` �F=�����,�w�   �r���244$���<���۹� ��MLL��̌$%%	`!�d�]p߳gOF`�$ �b��vE{; �)233���F`m����  "I�  �>�O��N9~�����
   p9�x��ly���F��/~a�  �;�上�
,T{��7���v���+�111Z�# l�����ӫ~��; �)v��)^�W`���Z=V  "	Mg ���;�C{�1�I  �)))RVV&����?Vll�l۶M~��_  p���a��'�g��\pא- �i�]��VC� �			���"�OVV� ��D� �Y'N��#G��7�    ����ˍ����叵c�y饗��  Υ���~���p7C���{ ,&''��>w ����!w�C[	�� �H��� gϞ  6�;���qn��\   ��-_S��-���T������v  �377'���.�Uܒ�v|���[nI��|;�햖�֝EN� nzaXI`]-11Q  �4���4� ���w�y�;vL���   �������####�?���p ��t���iݳgOƑ#G���p��|lH� a���~���h�  �M$���{$''KII�  �Μ9#  k||\���o�����	   p1mq3��T^^.yyyF8  �������`����ث۟��9>���x~o��- kLMM�{� �k�.�}tBA�]  �D��� @(�z�-9t�|�K_   �b����
�|��叵s�N��O�W  ��_43˸<,v�pM��z� �������r�g� ����B��mTTT�Rh ��F�; �O>�����ɵ�^+   �Ŋ��ehh�XM�JMMM������̌   wY\\�s��INN� V��qq8Gܯ������*`���P�� 7���'UUU @$#� 0�6l<xP��뙔  �KhkMM�����>Nll������/�,  �}tBwX�c��������ΊC9:�^XX����2���ֽw @8���JCC��z�=&&F  �d� f9��|��_��}�{���    �2])UWL��:�����ĉ���  ����466
`����ԝ���P���_�D���iYZZZ�~� �˽{�^�����$//O  �t� f:y�<�����~   .�+��={V,{���L������N  �2::j'�J�U~��&�����6�ޮ� �E��p��t����Z  �i����  `������V�ԧ>%   �2]1U�����>�Ν;	� �B:fq��9)((�*^���m��?! l����� ᢁ봴4��JKK%11Q  �t�����  `�{��XRZ[:  �e����d���1�����X�U�{   w������믏y�g�āp����5���Vn�qm�� �}�v����㥼�\  ���� ����}���ѣL   �%����W_��}0tL�g?��   wa�l�����ؾ)�؀����=+��ljjj��%� ���L���XO�G�  ��̙3 �U:;;�k_��q   �%%%+����Z�MMM������ܜ   �������Y
`)�j����|��x<�>KKKƇ�F��?  v۱c�p�h���tc�R  �w ��~����ݻ�3���   ��|>�>�@��}ill4>��pӕT���,��j�---r��	  �-�eeeX����8�c����V�޾ѕ���U  v������f��tYT  �	w ���^ٲe�q  ��h�U.��f�p]I���J�{�=�c�Ν�ꫯ2� ��p���rd��K_�R���B� ���7*�  � ]��*..���  �p �A�C���'O=��]  X@�;O�:e�;::dbbb������;n���^��d����R]]m�6  �{h��X�7�P��c���q������� ��^��̒gV-� �Z�a֊�����
  ����  v��鑯~��r�}�	  ��q�g��v��]Y����O*++p���y��,�[[w  \fzzژ�IQ���z������82�.��"�����O�; �n���RTT$����X �6~  ��������O�T  �������5̮A]�k�=X��p
��8�U��i�>55u��   ^��N�V�x<�7��;`3���h  ��v��!��^�.((  �͹s�X� `�x@���e�֭  V�a���n#����nj8W�y�u�	�:�BCl�L�X��땖����-  �=FFF��	�92�����_�� �Ѱ�f�� vJHH`������x �hcU3  k�k�{���ǏKFF�  ��gd__�>צ���~�K��E`���8���Z^^n<�����*����m��   �A'�����>����8����>�/] �fjjj�?C� `'m����XG����9 D'� �p��C=Ąc @�Ҡ���i�WC��־��d�cwuuISS� NQ\\l'nv�����4`�y  �aff������`����k{`먥~p��| �"� p���6�ubbbX� լl `=��կ��'����˿  �����@��fg�W��O�N�u�շ�z˒��w  �E[�	��bW	�u]% l��7�3z�, �E�����X���B��� �hE�;  �y�imm�m۶	  �H��5P�h�п�4ڴ���####�ﻮ���S�  �C�	(�����&�D9�� N�}�v�u�����N �f� ᶴ�$_��W�رc���%  ���瓾�>ioo7����˩Z������'�w]�@_Of�z����,/���   w�w�b�qT�}Ϟ=��M� ���%lw �]RSS���^`���jc�S  �w ���������F�  �� ��ٵ����Uc��w&��IHH������5}ߺr��/�,�� �;���E��
`��[o������pT�=>>�ぃg�5�M4ܮ�@�5O� `����-���K3   B� ����<������ ��MNNJww������qq+��޽[ �)//���!���3u����RVV&==��/ �uh�;wXiqqQ[�s�言{�U�6:�+� v�`{[[�������  ��0�=? �
����lL����+  'YXX0��5Ю�p�,)�������(\��,_���L߷��p �=FFF���R i��iqG�'� �ЋM�tI0� �'fk���Jbb�  �ho 8�����.9~�����	  ��zΤav�kvqqQ"���>}�h��F�	���ebb���nٲE������ ��i�;`1G��;&�gϞ���
`=IՁ�`p ء��U`���xj  ��  ':w��q���c�ILL�  `����������
���3�M�T�����k���Om�ojj�W^yE  ��i���H���"�E��ٳ'�ȑ#�8tL�=>>����' [���:w �Ւ����������.  "� p�W_}U>,7�|�  `����3�����Q�
���)�\s� N�A���"ӯcl۶MN�8a��   �O��	��Bq			;�_�8&�.��"�6�댮`,--7  ���!4�YCOv���  |H�� ����_�U���	� L��Z�O�:��ϑ����277'			8���h�mqqѴ}fggKii����
  p���� �J����B��R~��J`]J0�ش� ����"�Fuu�x<  �� �dz����r��1)..  �1::z!Ю-���Gi�_O���8Qll�����S3���p �%�������܎	�8�D:�kaaA  ��.�Iø5��%33S  �� � p���	ٿ�<���'  �gjj�hf_����6��;�N�Pt5���Y����� ����i�> �5��Z��u�v�
^��c����v�m����U�r�<033���� ����a�2  >��; ��~�my��e�޽ �������k@[�s�]�9���p2��k\���Lۧ6�777ˉ'  8�ٳg	��2�sɢ[n����G�������M�{�崽=�Z� Vҋ���XC[]8� �Rz�L�! �-�;&۷o�뮻N  ��'O�l�k�����Q������������r��y�����J�  ��s���
����5�M�]�|���v�:x
�  +���Kbb��\111R^^.  �R�� ��{�V��(499)���F�]��f[q)�_q�8YUU���曦�OC�������/  ��tR&`%�߿+���p�=p�z��X"���瓙����A� `�����4�/  �R� �FL���'G���� D.����3��|��/6��7w8]FF����pkkk�  ���ޒ����nq G���`1�u2	w �U�b,�h�O�u  |�  7���o|�r�]w	  r����h�ZC��־��$��������tU3�[�l��{N  8������`�+�����g�y&�'�a��|��U���|`���������(  XA��00�^��z�  >��; ��~��ʶm��ӟ��  �ktt�B�]����s迃�X����d���RTTd��]!���N�}�]  �644D�VJ���ol�	�_"�wqH�=�|>���Ά������� X�ۛ���JKK���<  +#� p����u�V��� �;hpz9Ю���1�3�w�Ayy�p3kŇ��&�  ����8��R��f��;�x�� ����9��Rd  �TTTHFF��\�� `m�� �[iHr�޽��OJJJ�  �G��P{{{����R&�p��'?)�����Kii�tww��?WHMM���I  ΥY����Kzz� V�]��_��wpB�}7�H �MMM�����y �
���sis;�  X�  �;u�|�k_3�� �0::z������X!tlT�À�i�]'Ә�~��]%��_  �\:qvpp��;,���
k���믏	�v Ki;���l��!� �BBB����	̣��  �N�qϝ;'  ��O�Sٵk�|��� ���dJ'-�����d������t^�W��˥��Ô����p �t�C��L�
��V�m�ݖ���΄��ր{aaa���c�L�b�$��p X���Ibcþ�PD)))���$  ���v3Ε p����h�lhh ���vo�kS;��K��	��-


����F6 T������/CCC  �����233#���X nnnn{`�_���5I������#���9�� Vhmm�G'���	  X��P  �z�v߾}��SOIjj�  ̣�u=�0��{zzdqqQ���p��TUU�;�c�������?��   �҉m����a��1�n�ր�����lv�Z>�OfggM�w �����V�G�!� ��p Dm����`ij ��D:;;��ɓ���eJ#2�gxxX&&&$==] 7��Ζ��Ly_�:�/�K#o   �iiiIFFF��ׂ`�]�|�&_�~�n`)��f�D]r  3��n���)**  �>� �H������O?-���� �qZ����g4vkS{� J�۷o�-�����^y?)))RYYi�'  �:���������5�����={��$ ,555e�~t�Efg ���z���Q`���
��
  �G` �|�A�q���M  +�r(����M0�:u�q0�H�#��&L��ϗ��������L�  ��l����"57�tSΡC�F���a�'$$���|am�"�^����5e_�\ �������0GRR�q�  l� �H�e%����ǏKff�  >4::z!����)sss�G�+:!����:�r��ِ'����+��~	 �si�]�9f�E<��֮��'�x�̗����Xkzz���2w ��ho7�^��� ��#� �d���r��y衇X�@�Ҡ�6�/�����,o���"�">>^������/�����JCC����  �iaa���wX����h�{��]fo�L/��E? 0K\\���s���INN�  ��YZZ���a  ������}O���J  �
===F�]��uR+��0�>���m��ʌ������&�  8�N��wXdg�8lw����i �;��e� f���7D`���J  ���r  �:t�%�޽[  ���a���{�؆�V�ϭ���Z 7�����Rc%�P�>233ellL  �3i�]s��d�wX ���rK��� �Y��2w ������2.. ���&G  ����;�S�?.��� n799)���F�vGG�LLL`5}���	nRRR"�O�i�v���_|Q  �3i�]�i^�wX��_�bᣏ>:`���,p��  ,�\f"� 0��PUUU	�QQQ!  `s��� �h122b��>,� p����3�ڢ��U�,x6B��r����M�د���x�Ess�����  8��쬱j���4wX����l~l��%�8�[e=-tF��� �������I�}/--M  ���� �6���9rDn�� '���kSC�*֠n��$�7***2Z����އ�"[\\l�  8��Gi�=..N �DO�]>��`��#f�}i3  fХ,a���r  �G� ����H[[�\u�U N2::z!Ю[�K� 3tvv���
�6�-�����p ��4��x�枘�(���~XJ��p����~`���v �Y��C�B���III  �y� �H�L��9v��� �J[�O�:%���F�]����䤤��
�6������gނ���>��s�� �C鱪f47H�f�x<a)5�=���/~Q����e� �j�֭z�+��io  x� �j||\���o���l5 ������-�n7s%b�~��x��j(��,�)�<y2�}hP���֘�  �g9/855%�������[n�{�G��|P��111�}>�W XB[/̞5M� `�#tڴǬk  ���m�  Z���[�裏ʭ��* `me_�wvv�W���s��;�*??�hq�,�����;  ���h�w%$$\�f������S;�������) ,cv{�ZXX  B��윜Ahbbb���L  @pΞ=�D����  ��IDATn @�;z�����ʵ�^+ `m	�fv�wtt��Ą �F��:i�UJ�F����������A�Z��㹮 �C�y��5?H�f���{�`+ ̠�]II�q  �̙3 @��p�������8����r���^#��z���-@$;��M؀���JZZ��\F\\���Ԅ�  �р{vv������d����#�N�;`��hE�:w @����{�bcc���T  @����  |�۷o�<��L��.�k�]��j�����E����������w�	��u���;  δ\���j���zLf{����={�$6[�%t��� B��^���
B��cbb  �w  �ǻ�+>��t��MNNJww�����ɓ'effF�h�<���J�J[]���ebb"�����������  �,zζ��dd
4�N�&��馛r:4b��p�`���~9�E�ga�I9�h� D���&Ah�䳨�H  @h� p������"��ԧ@t�£��>#��-լ~|TWW�ш��mnUYY)o��fP?�����:y��  8���4?���fl3330����nl���m=�
��v
 K,/-b6��  ���z������ɂ  ��p ���^ill���*=t�G��5̮�vmk׶? �ӱ���^>3�jF�mll,��ohh � �C-�5G�Ǯqqq����i<2�;�%�hoWV�� ѥ���X����_AA�  ���B	 �G���}���ѣG%11Q D�����v����
����w��������A��>�����  �����Y'�&�5nk�����	�w �SmݺU���2�� 0����  �������O��9t�����B�=ض^ �C?3���:�L�]����ܹs��Y�Е{�z�-  �255u���a��v>�m�={�$���`:].rnnΒ}p �">>�&��� �y4�333#  `e���!۷o��|�3��|>����I{{��2}����0���4,���,��i�{0w���H�  ZXX0r��3Э�
cbb0I��7ޘu���Q;̶�{\\\���D��b��I� �Ph�Gl,���(--��  ����  X۽��+[�l1n �att��kC{GGc;��t\VWFhjj��RRR$//O���7����_�  �A��p_���������Ҏ�-m8����x���W�[\\4f]�v�ϡ�Y]  �����g|aa�   sh�  X�c���'O=��Z�<������}!�>11! 쥯?����Aܵ�GK�^�u  ΢�����&��E^����	 K茫�YW�� ]�r9��au������5��Zh�  K��UUU������� ��� �1===�կ~U��>~:����kj��]�k�Z���������A��744p ��fff.�yvv���;�Y�~�mYp�����tՄ���!Õ�Е���M�;  X555k��fd�����  �p `�}�Y��+��� �ұ=v�0��hu҉�� p���19{�����
�vZ�L�]��uş��)  Ρ��z^��A�j�]'�f<�l˂ے8:x�7p0�" G?�4|�����K����v  [�lO/3�  s���  ظo~����,����Z����]]]F ���k��;"���srrddddS?�Y���z��o~#  �94�777w!���a��1��={��9r���d[��Ν�	lR��p� ,m�����v  �A�;  ��%({��cǎIFF� 0���������ݸi���脔ݻw	***6pW:��;  Σ�����̌ &J���ol߲��l	�/..���M �B� ,�kH���  kp `��������C	c=@�|>�\hi?u��5 g}s-�@[ܳ��6=᪴�TRSSerrR  �sh�/;;���6����^�&h�H	�{<�6�:� �jhh��v  �155%�ϟ  �y��կ�������_�� �8	.�;;;�%�D�������ـ�N��1�'N  p����p�Y|>�f¿o���p�& \��I  �Ѐ�6�#8eee4�  `���~  ��ַ�%---�mC>�j4@���h��萉�	�twD���4��̔���M�\cc#w  ��ܟ��j-�Il�@hW��w��� ������x���䀢�"  �;s�  ���r�_��W�رc�����(===F�]C�z����@������"�N��l�]�5222d||\  �3蹩f������^XX0n�I B��xlɄ[p��۲��������-  6���^�� ��  �npp��?�補�"j�ɓ'�P���5� z���]�N�����Z����cC���   ��U�.>N�,�~�&Ȼ�曋���o[:�fy�}nn�Mf�w �f���JMM�`�ho �Z4� `��_~Y�x�	��������tww�v��?^ `�6c�:uJ������oo�g� �<:�b�a2mqww�ݮ*z ���f��� �ͨ��������� ��� `��{L�����+� ������h���X	������;"IVV����mjRWII�����  �3h����|W3�111����i6��Y����Ô> ��|  �e����� ��� `��'w�u�?~\���p3m_�cE�kHU��u� 6J�;�H��<������x�~�x�  �0;;k\�Y.���_��4 Tv���p�& \G�$ `3t�omm�`�ho �z� 0׹s��;�0��i��ی��^��M� X����+�zD����M7����p �A��)))���@�0���pK��f-.��� 6���J�K{;  ���3�  �\����p�馛p2����h 0�N�ٹs� ����|S-�/���  �Aχ/��o���+@����ٓ|��˂����z�^RN�p lVCC�`�JJJho �b�ޮl ���x�	ijj�k��F ��%���ɓ�����  ����4�➜���쀮�eH��  ����q=_�R���DB����ؾl�Xp�z�m��ty  6J�555������  X���_  �544|��A9v�.�b�6(kȴ����X ����0����6X���%� ���4QM�F�fXZZҌ�;��VN� w�� ���$'@������8  ���N  `���	ٿ�<�����6������m�;;;e||\  \�<����RZZ*@$��˓����i�]�}�  �������ū�S|�x<KK�-���-���  l�^��敔�  �w  ����o˷��-��,������kS��i[2 8��7pG��RKmq?y���eHz��  �Oϛ5���r�kz~�7J
���b����4�`�_�5�?�  ���I�}�


$!!A  ��� `�cǎɶm��� T:V��q�P���...
 8��W}� �����ó�����p �9.�/��;B���--A�,�~�7f6TR.��4	  �A�4���� �}� `$�s�=RSS#���l����@{WW�LOO ���21??/���D-:�1����ݿ��N~���
  �ҹ�����Q��={��9b�@�e����f��;q� ���o^NN�$''  �G�   {���}���ѣGY��� h__�h�`;�m �liiIN�:%���D-;�V����u�!yyy244$   �4�~9]�E�^�W�P���56�
������� 6������ �}t���ٳ  ����!��O�$w�y� �&W]]g��]��f�$��F��H�oEEE��ӳ��k�;w  �A�z>���,��֐;�|U๤Y�g�طe������ w"� ب��T���l\ff&K} `���ABS  ������K[[�|�ӟD��������N��� �T�^D���c啍\gщ/���  ��[�'%%]�u�p�	��ڱe�ߥ��w �Fi�ų|�>�� ��6� ����׿.[�n���jA����2�ٗ���� �bxxX&&&(9AD�������]k�r$-�  ~f�<����B�e�V�۲��X��`-� �����l\JJ�dee	  �w  �GO���+O>��qN�ȴ��(===F�]�����U�D3}?ܾ}� �HK|6z�EǐN�8!   �4���}�ז��d~~^����fŵ��A��o���b������t� ���INyy�`����  ؋�;  �M���� ��{� r���J{{�q�p��� "��H���(���r���u﫫 p �V���	�#D�7�|s巿��.�wlI����5{<�N4� 6����X��|�  ؋�;  �����Dv��%�'"p���I���6B�'O����� `e�^�+Y��@������~III� � �y��1��322�f�w�/�f�J4�  6���F�qz!�  ����/   ���>ill�������}}}FH�>0&�@8 `}���""QZZ�������Ě��z�R]]-��  ��ZZZ2��.��~M�#@�~���f�ת��&�J�� 6B��zQ'  �G�;  Π���퓧�zJRSS΢�u=n�0��ڵ�]� ���S�dZ����{���:�  8��/������YIII �dƭ
����˃ 6�����M���T  ����dppP  �3���ʁ���&��9����@�n  �tvv�'>�	"UNN�$''�[��eIZ�+� ���������N�!�$3nE�]�H6
 W���  �SSS#�]ʫ��P  �����eqqQ  �s�򗿔���g�g{��r�]occc �FOO���`/�����c���k����8  ���v&����L�3=�~�7V6i���� �����
6���Xbc�Z8	  ��̙3  �����FikkXGW��j?u��5 ��t�uww7���������ٵŝ�;  ���+KKKL�D������ߚ�Sӓ6111�~�_ �����  ����L����O�[׀;  ���~  Σ��������Ǎ�0���,�;;;ennN  ����ɼ^���!�����=��  ����1��5����!@�ǆ�����o ���L-  �qA~����$>>^  @x�� �sʁ��6&�#8SSSF�L�211!  gЉF�G$@$+**���^��u5:�Qoccc  �kfffŀ���,w��)p{���p�x<4�.���L  ����N�1���  �;  ���/����=���?/����!2�k3��0. �444$������*@��������uW���W_}U  @xi�===�#_׀���3Vh�aE9��[�+��v �Zmo��nNII  >� p�C�Ikk��رC�Q^�c�k�����XR �|�����9D����u����� p ��D�]���$))I� 5��CS��� W�%a X�6l0cwcJJJ  �w  �oiiI���'Ǐ���\�m����r��I�����i ��NN"��H/yyy2<<��}4�m�L�  ���}5~'���<x0>p�7k���GFF���K  k����/11Q���  ��r�)  p������;����Q9�~~~^�����6��׀
 p���秬��H����qqq�}t�  ��v|�Z�;�AqCCC5��o�ڡ�����/���k�;wN  X���p�mog� ���s\]N  ��+��"��/�"_��$�-O��0���O�:%>�O  �GW����"YJJ�dff���ت��1&�  ��^�А�JM��j+��
�Fqj�=&&�Q_  ����� �jtyI�@�����  �ho �}4����*W]u�D�����v���$8  ���?׌��g��{MM����?  ^�ԾR�}�{iii���6��?S�>����J���zBB�  ����j��
��;  /�  �����u�]r��q���7���6J��k��  �M?"q�p���l#,���վ�^�;  ��Z��	�#�!7s��=���{ ����  ֢KGb}���  ¯��_  ��h��������?�%�u	#ĨM�:َU� �ԩS�焛>׀`�B�ѱ����7  �g��h��
G7�l �t��Y�f ����3����rss%11Q  @��� �{���[r��!���[��4��.�wtt����  p������DQAW��������p  ��
���zr'��`��~mp���؟i�[o��`qq1G ����0w �������� &  �� p��G�Jkk�\{�����F`k9��ʨ �����:������u���
�>�� ��t�Z+pGRn��ֲ�~�ǌ��p���o�z���4���x ��h�֖��*���  ���;  ��������量�>lʗw5��M�z|�/  6K?K���@�h��n�]���KKK�I�   |4Į�վkaaA[ܝp���i��^���jZ  TVV
�F{;  �B�  �ӆ������?.���?��s�1���5����c4� *�|������"]RR�dee��h�w  �kfffլ��ܜ�|>���<o����/��'t�π;MOOM4  �$##C�����A���<  Πa8   �{�w䡇��o�ݒ�k�j9Ю[� �l:����K����EEEk��_  ���豫��u��Y��O�Y�2-ன{�w�U ��TUU	�V\\,L� �9���  D���~�~�S�
y_���F�������� �l:���;��'%&&����G����k�+���  ��&���	�#H�����`/� ��p_�.�UXX(  �9t�w  Y��^ٺu�TVVn��tI큁�-�N�2� ���s�Z
��@z�{z���  ��NB�B�Պ�V��lP�Y;2%�w�ޔ���R�J###� +��vEE�`u'  �9� y������o��G�m�k�V��@{gg���6  �m�gϞ5ګ�h��'�M.$� @x�糮r������dii�L!���M7�:th$��p���j�z��Jz!�` `%ڮ��	>��#  �,� �LV��������|}jj�Oi����C&&&  '�	X�-bcc���J�itU-Ybe  �gfff�<���ka@rr� ���x����P�cJ�=&&�Q�� �gqq�h�K  .�X]VV't  8P�  �����HZ[[���5(��)Ʃ  n���v��-@�(**Z1�/%%%���+   <�[�N��!���(N	��|���w��FF>\	BgG p9�k��  g�� �Ȣׯ���kjjNVTT�����=������18 p���.����YD������0J�.�cP� ��evvV� 5��S��Bp���  .����
kХ���  8w  �/''�_[[;T^^�bkk��u�]?�x<����v�mW�������v �����K__�>���ԾR����B  @��`_XX���%���)�r��[����ٳg%6֔� @�����Ef��&� �<���+�  gKJJ���ƙ����~�3�y�ꫯ>��K/�3�<#w�}�%�����_��U���5 �������U����R��Ct���F���ܜ   ��g��~��=h�{jj� �To�NBN�<x�;<<��C��hp ����Z�2=���  g��  w�I��������WTT��ꫯ~�s��ܩ�^{�����߿�>?�����ޑ��$ �%4�~��
-tLEK����.���������޽@�Y��������&_�H�-�rmh-���m:�v���}�:�����I��z��Cn�BZ�ݍ�a�ݙ3L]0g�3�͸CnHز�\d'Nb���t�:u���&Y��|?kiI�+�$��{�=�  D�
���Ԁ���<wLBQYYY|��7��r��������!`P*�~�� @_����Z�/   �p  z����͛�+**zk�?Y�b�[�%4E����'�y[�l��iӦ����z����i�  �p�̙P���Ѕjkohh���ϝN'w  f�
�_+;��[�I��������GS��)�e���D^{{{h����d `8�NMM�N5�  �����  D���4Y�`AKaa�o��?���~^RR�;�|�ʕS�o�ر�׫W�~��ɓ+U�  �Nm���-�7o� �������ijj���  f�
���7c���~���`�T�|f����5� �Q��ʟ�ٟ	  �qBql�U�Zx  `f�� ��Q�].Wo�v��p���/y�ҥK��9Z�y���w�y晇|��{Ξ=KR `����;t�������
���.�� 03T9����w�(�-��gL9�n�X��� 03� �B�}l�,  �^� �,����x<'Ǜ��z볫V�:VSSZv�����9n���[�������S �(W[[+�nRRRd������v�g�PS]����  D�
���5���L�td˧p��k�ЅB�� ém��n|��f���
  �^� ���L�8�RXX�ۅ��������E��ղC��؟k�ʕk׮��������  �XKKK薑�!�Nl6�Uw��;  3G���@('r�� �0�l���F�Z+7���11�� \�j��Z4�Ij�L� �� 0��n�v�\ǂ�_|��_���w��z������hRQQ�ֆ����l��� @4�z��h�"t��A�u``��ϘU ���Ο�������eppP���%..N�	����������B`8�����/  �p8����  ��I؋/
  ���9x�7��__�h�s˖-�9z�hh�Ν;%��޽{���˗�9sf�  ��CG��O�	�|�+?��ʒY�fIGG�  �����f�]Q-��1A�u��%�ݻ�{�0��{ss�+x�ZХK�BӋ�B ���ѥ���N� �����:�  ���p���

��t�M?޶mۯ-�a7��������?�.  D�����1lp�+�Nl6�Uw�P�K'N�  y���2{��k�F�Uf����U��0��{�G �P�w �p�$��n|R~~�  ��6��(  [RR�̛7���t�V�w�}/�}��=UUUr��ay���������n�zogg��1 @R!!u;g�t���
ȵ��_��*_"� ��P����`����1���{ (a41`L��]!� �j�JJJ��j����  �  |RLL����~���u:���s�=���p����������<���]�v�����  �Qmm-whI���
  ��	��s+���'�xY,����J������ �Ѩ�|R^^^(   �w  �$???0o�<_QQ�[.�Ɋ+޲X,�̌���TTT<�r��%�N��M  �B^�W��Nt���-uuu200z���.iiir��e  ����;�ש <wL�*Q����p� C"� ���|�
� ��G� ����d�?���������7��7�pC���+W���}��;�/_�t���l  ʜ>}:(JHH@'�TH�܇��Qר� y�����O����:pOMM`�f��=�w������#���; `Hpǒ�QdddHRR�  ��G� �un��r�o'ǫ_���-]����w�	-ߺu� t�ÿy���������	q @T������ ݂Џ�f��\�����_  @���x��M�@g��u��%���������Q�*� �b�Z	r�B�`  ����  3�z<������ŋ��Y������в�
F�}��?l���zj``@  �&^���;����j�moo=Ww  03ԬBף���y��ة�jC#y�V���o߾�ɼy�kZ�;x# g(�N{; `8N~��633S  @�S'V���  3Q��͟?�����.��g>��w�}w(�}��!���ڵk�U���<y� @���@WyyyW�*잞�.���  "k<wE��Ϛ5K�����*k~t2��P
�E� 0���yF���e�  �ܹs��;  F�Zϝ;�������q���˿|��{��<r�TVV
��g���<��+  D�.H[[�̞=[ �dggK]]ݕs:�����{�	  �,\���c�T�<��@ � �4pg� ��.((\M5�   chll  ���t�x㍵���.\��o��oj���C˞}�Y���X,���֞������8  Jx�^	��Uʗ��s弎�VE� �țH�;0A�ΚO%�� �D�; `$��*III�?Q����<  `� F���p���

��t�M?޶mۯU�Z�7>�������>  ���p��T�����*e
�=  ��9��/111�|���@�F�.&`�Y�e��p�h�����c� �!N�Sp��\f+ �H� ��P��xڂ���:�W��Η�.]�]UU%���{LY�v�za͚5QWW�W @n�B�^�t3k֬Э��CRRR$33S.^�(   �T�p<ň��]m�����H��w������ �!�C�'j�qVV�   � � ��骸����r�����r�-�=�����ա����̼��~���9���� ���꒦�&��l�H�����9s�p `pG8������b���IAD� 0�j�!�~�����N�  ����  fJ~~~`޼y�����.\���+W�����в���'�蔕�uKwww}KKK�  0ü^/wh+''G���eppP�v�����  Y*�>*�L���|�;�/��҄W�I�/^�蔩���!Cwf$� P�V�F��D5�   c�� I���2��˥����?��o~�n��>�����7>����������^�  0�T����� :R�|�|H�d�� @�7�>00�F�.�)&))Ie�?��'R������0�ZZZB�l`  Cho�ZJJ
�i `0�@@Ν;'  ��:��r�z�����Wo��}���w��y���[�
�驧�:�aÆ�}��G�]�S  0SN�:%}}}/��T��
�gdd���tvv
  ���4��ת�50111���{ p��g �s����=w ��0�F{;  �s�P  ��d��=O���xs����֬Y�~MMMh����{�������oll,  f�j�T!w��-��RSS�����eh�  D�D��1n*s>��M*�n�X��ᨋ�]]]��� C���ĩ��  ����(  L�j��?~���8�v���?x=x��W�:$0����Ž��g/]��$  ���K�ZS%D�{��]p  ��~����K\\�u_;�0<0�����A�J��Y---W��N�� 05�6--M�1��:��5  ]� &#!!An��n��u,x��]w�u`ɒ%mC��q�>�|�ɖu������������i� 3���V��^t�J����(g `��f��d&T^�cbb��H7����A`,��4� ��.����\  ���� ���l�,��x<�\�x����w�G�-۹s�@o{��}uÆ�>���\ ̄��f���Y�f	�#���̔���Pi��  �����U�M�k���ק2�yߤ�M��Y���Wp (4`�I||����  0� c���
����Gn��o۶���%��o0�ݻw�Y�b�N�>}�  a*(��z�S��� ���ɑ�/�J�Ξ=+   rzzz��Z� �9W3&N�Qb���kצ���g á� 0�?���S�F  w �uQ��v��<�������cɒ%�UUUr��ay�����~������6�?��\ @�p��T��joW�p  �Th=���f�Y�&�駟>7�7M8�>00� �D� 0���|L5�   c"� ����Q�������̙��o���e˖5;v,���?�� ��o�s�ڵ������[�  A*ச�)d���>~vv6%M  ̀���'�����܃R.`8~�_���B�	� �X�0 ���.���  ���; �%??�?o޼Ƣ���.\���+W���>�(�����L�����6n�X\�����  DJGG�477SP���_5���j�  �p�`K����>����z��={"�T����p���`�1w �B�ş�� �q���Jww�  �+99YJJJڂ��\�p�K��{�+�-� �v���؊+��>}�f  �jkk	�Ck�gϖ��L��ȐK�.	  �Z���wh]��p�8M�\}�w��R$ �����c�  %??_��v�j�
  0&���|�q�����N8�W/^��<p���Z~���֭[����������kjjJ  "����m��&��� U�D� �ȚH+�j|�c2�s�Mp �D����	Ҙ�  ���� `|6�m���48�7?��O�۸q��555�e`�����mݺ����η���9�  �������	G: �P����v9v�  ��Q��f��k�q*��&��>�x 3OM�>��;  ==}�$f�N�  �� �)x\(--=_PPp����'�x�5���W�:$@4	���]�z�����  ­��_N�>-EE.9L#!!A����k�	  ���>^�<	31NΞOh��ַ��R��p�7��A ������$IMM  `\��T8�n�v�\ǂ�_�u�]�,Y�VUUZ^^^.@4{�g�X�r�WO�:u�  ^���;��`��е���n  ����;�דG�8�Z�*a߾}�^�&�V����`M�w �p��:�HNN�   c#� ��f�.X�������3��̾�~��uG�-۹s� F������+�Μ9�-  ��
��_@g��١Ҧ��Z  �1р{OO����p1��=x��
���~� 05�YmH�p ���1ub  ��� @t���
����Gn��o۶���%��o`��ٿy����ڪ�7
�  a�twvv��T����p  ����&���⡯@ �2��	����LKK˕�111�$�  �G�;(5554�%  06�`�c*����t:�u8��w�}/�}��=UUUr��ay��0��۷�aÆ뺺��  ����^,X ��n��f�կ~%   2E��_����_�g�r���ד���~���jmm���v ��f��"(''G  ���&���v D�:�,..�u�\'ǫ��~�s˖-k���-߿� :ؽ{��=����$  ����%����9��  ���>ހ���^O� �aBt�._�|�1w ��9s"V�U  ���|> �W~~����4�%�,--=��}�ݚ��в�
��}��ݻ|�r�ٳg� �0Qw@w���b�ۥ��A  @d��zJJʄ^O��c�X�p��� �#�.���:!
  ����Q  �+99YJJJڂ��\�p�K��{�+�-� W�X,��۷���룖��8  �u�.P��y<�  D�
������ �F� 0�b���=�]NN�   �#� S����o�����o޿nݺ���j���.[�n �ۼy��6<����B__�  �ŝ�;t7�|y�7  D�D�sp�8�5�� �3<�;ѯ= �L��Ҵ�*&&F���  w ���6��xǛ,x��G=��S��~�30~�w�~qݺuKjkk�  �@��z�謤�D  @�L4�������_�����(++�	���y񸓮�V����)�P:;;C�!4������Dw*���  s��| �����@ii�����#%%%/<����X,0-�����|��ٳg�	 0����C�!U��*x,#������#   �&�Ȯ�C����\��q�� '� �ޮ� �p���  `4����n�v:�G���+o�馟>��]UUU�����`zeff~�������%A  �F}}}r��i	��	�+5����HN�8!   �dpppBYCp�5k� ���,��܃8Z�����c����~ М��n5Z8==]  �9p�?��l���������}�s{��o����ѣ 2���ׯ_�www�COO�E  �F^���;��v�	� Aj�eRRҸ_?��whIؼ=������w��@oj������١  `|�DiKK� ��233%%%�

�,X�������׃�;����7��/��۳g��ׯ_�RMMͲ@    Lp��{�Y��G  @��0	������燎�3�,:��p IKK���D�YNN�   sP��� �Dϕ���9��w�+_���^X�dIoUU�>|X�������gϞ�._���gΜ!� �6gϞ���.INN@W��  D�
�O��f�Z�uϥ��,K�x_K�09� �!��������T  �� `f�騸����r�p8�.\��+W6UWW���߿_ D����[�V��.�B Ljhh�y��	�+��j����  ~*�>Q����;��w #� �{���v  ����	 �M~~��ܹg���ϛ7��֭[߫�� �RQQѺv�ڥ����X �i��z	�Ck,���  ��Sa�H��!�@B���*��; �M��{vv�   ���$''KIII���|w�ܹ?��W��ӻ�{@ ^EE�/ׯ_�LMM�պ �T1�q��� ���6���7����~75x�! �������@_�ErssEW�����  0� �H��+,,�.**z?''�/^�ܺu�Z�������e�Ν�<��ٳvŊ_8}�� `�Եߖ��� �}��;  ����e``@bc'ҽͤ._�<���-�{�֢��x���|��U��p �����$11QtE{;  �C��Q�l�A����p8ޜ?��[�l����-{�������[z{{ϝ?>U  ����ZY�x� �
[	  �VW����wr�����Q����{p- ����v�� �)//OtF�  �!� Z���JKK�)))y�'����b	 -=����7n�Zgg�[�'� S�Jp��l6����Hp�J  @������	�G������=x���^7��{ �c�X��opW#����t������  ���޲��Y  $$$�ܹsۜN��㕛n��<�@WUUUhyyy� �ۮ]��m�ڵ������� �d�%*��u_hK��n�[���  ��
�O&�\Kp��>�׍+�3G$0����* `.:ܭV�   s9w�0�l6۠��i(..~m��Ż�/_~���k���شbŊ/�>}�3 �$����ٳg�nW0����  DH��ߣZ���kQ���yݸ�~����w ����rssEWYYY  ����	 DRfff����|AA�������Zcc���7��^xA `<rrrn���?��Ԕ.  L���%���w  *�>Q*ܮ������fZ܃6��<��6���W�p }���Ibb��H��9h �|T� �IC����9��w�+_���^X�dIoUU�>|X `2����֮]�����߶��s� 0)*�~�w
�+�  DNoo��GVc��w��W�* ���v��; �+//Ote�Z  �w �-&&F���{].�	������]���д���� �Gׯ_����k���  0Q�O��Б��
�._�,   �&��>��A���>޴<��A� 0��;  0� ���f�x<��M��}���콚��p۳gϓ�W��j}}��  �����ɓj�!tU\\,G�  ^��O��ژ�����ߟ�� �22�;��,  �5�>{�l�� �������d)))is:�����x�b�� f��O?}��+Ϝ9�#  L���%����n�  D��}N�&Z���߯��US� ��u����=���ל�纉׸��q%�D� �:X����� �y�|>�뉉�Q�~�.����x�ӟ���=��������~Z `��6�7o���������4�  &D���w  ��]��L�
������F��l����m�( �pW�������$11QtD�  sRS��;wN `46�m���48�7o��ƊM�6���� �F۷o��ƍWwvv>700   �ׅ���U����Qaa�  ��PA����'����lz����^s݀��b��0��w��@_��٢�ٳgs� �I5770 C�������

�������O��b� b׮]֬Y������  �v��7�,��l6[�:�
� ��R�H�zO6�w��� ] `^���@_*���x�
g�����[n�˖-멪�
-/// 0����%˗/?d  ����p���,�]  �_����@4\������9� �7��tuu]�fG� �E�  ���� z���p��5���<��;v�8u�رв ��yb���uwwt�ҥ8 `T�]e9(,���N'w  "`�M�*����CӀQ̹��p�`v� c�ޮp }�pOMM�:  s��0����@II�����#,8�������& 3ۼy��Gy䁎���� 0��ݡc���|tTTT$   �&��c�s����d�X�pχ �.�/_��9w Г�����!��ִ�  ]p�G]�(--ms:��:�W��Ο,]�����J>, ���;w��nݺ%����	  �Z�	�CW���  �o*�{{{	�cT�@�~�׌'�nW#) G{{�U�	���������I�� �yp�O���\�����_�v��������� �j�޽�Z�|y��3g
 ��P�;�C p  2Bm��e��e�:\���eee����9�P:::�zN� ��c�yjj*� 09�1�l�A����p8�,**z�?�AuMM�  >)##㶮���K�.%  �p�ԩPh(>>^ ݤ���f2nii  >*����?�}N���!kݺuI{�������?�f�XH�3��]��"� z�1�n�Z  ��:����$ �_rr�jio���;����C�^�X,~ \Wyyy�m��kWW�/zzz&^� ����`(��v�Б��$� @L6����>+�E�&�~��c-�f�=̴̙ f���; �w  `6�.]���}bbbT����r�p8�Ο?����t�ر����J ���?�O�ׯ�qMM��j�  c�z�ܡ���By��  ���5(%%e��MJJ`����L6�n�X���ttt\yL� ��[�}֬Y���(  ��@���l�����p�9���[�l����F  �cϞ=<��Cw744�  c����{�W ��;  ?��>Y�1���۵�_/�~�7�>��n���; �)!!!��	��  �w`f���JKK�q��/�����b�P+ a{��j={�d `��͡4ݮ	 
w  "C��g�0��k-�^�=�icioo��9w Гjo�ˉN���  ���� �/���ks:��:�W��Η�.]�]UUZ�}�v �WEEE��?����������d `\T����ʧ>�)t<^U͟���  ��T�{{{����!��Q��#� zRw�$&&Jr2Ef  ��@������������׃�;v�8U]]Z��~ D�SO=��M�6�=q���S FC��������|9s�  ��J���@h0���0����� ��� Pt��� ���/##�_\\����������vSS�  �ˎ;�?��C_nhhX   ���j�n3�Jaa!w  �l*�
ȫ�B`��܃?6�  c�� �X�V�	w  �@��:u�����n��gvv��.�����l@  Q�[n�lOOO�s�R �a�5����Knn� �Q���  >*�>���1۵^3�\!ip�w ��S�{ll�̞=[  ��p&NM�Z\\��r�N8�WKKK�ݸq��cǎ	 �X���ownڴiIGG�o:;;�� p��N�:r:�  �O��&�^`�npWC-r����p;���~RSS�������  ���Igg� �>��6��xǛ����_SS#  �۱cǿ�_������-~�_  ���v� �)**  ~�ŝ�;�����,v�Yf���Z���������� ��S{����%  ��hoƖ��$.���n��Z�/:t�e��B� LjϞ=[W�^�����[ �?:y��f=t���:.���  >S	��p| ��#�\�pA��F[8�M��Ǧ��`���W�p =�pW�  ��|>� ��:o[\\��r�N����O����Ν;ۏ?Z^YY)  s��̼����)��ĉ @�
��:uJ~@'����@>��C  ��7'K��U�=>>^���F�L4�n�X���ttt�6C����V��"==�6  4A�;tg��=O���xs���{�l��AMM�  �TVVַv��/��������� ���K�Z***"� @�M��]���%��ь�U�V��;`0*�>w ГN�  �@��IKK̝;�|AA����byy�/-K@  ������6l�Z[[����  p�җ�$�n�  ��J���܁�,�m�e�jp�M �Sgg�U�	��~��p������YYY  �@�f��㔔�tx<��9�W-Z��e�z���B˷o�.  ��{��k֬YRWW�� �^SSS�qJJ� :�3g�  ��j@]5������ �Y�fi3�Srr�$&&
  Ѓ���l�����nwmnn��N�s�SO=u��>  &�����|�\p�*  ��������.   ��p���`��1L�X��&B�;  33StA{;  z��f�_7����kAA�s���[5, 0�ſy��;��������
 @k���ܡ�������r�  �m��Y5S}��f���Z@�0����Ebbb ���:�] �]ww�\�|Y �Q3����9��w�+w�y�O�.]JM `�m߾���7����xn``@  ��z��Fe#l6��:uJ  @x��~�R�jq'���̪_+�n �2����v Г.�ou����*  @>�O #Pԋ��{].�	���j�~ߖ-[����C����/  �ˮ]��Y���uuu_ ������b�Z�ɜ9s� f��}������T��w�`��cc�� t���!:���
�V  ����(@���������,**z���`�Ν;O���  3���b�ʕ+Ϝ>}:_  ڪ��%��;  ������c�����]�n]RpEJ ������s�@O*��]�� ���#�$%%���d�۫�V�ˇ��X,���* `��mҺu��HOO�����9�@S^�W>���
��  ��T��1��+V�z��:F.5�\�r���p����; �'&&FfϞ-f������  胀;f���.**�)((x/;;��ܹ�����啕� @4ٻwoݣ�>�߻��^��1 ���ɓ288�5ch��;  �7�w���~*F
*�>����b�Vm� ������l @?���٩p;�9  �����$��6��xǛn�{oYY��  �x��'�n�����裏�
 @;j�ә3g��t
���.   ��c ��5S*0$&&&;xW7��܃���tt\=��� �G�u���%  @/4�#����s��=_PPp��v��}��a� ݞ={�����o9s�L�  ���p�N�,ǩ�����.   <���p�(Fͬ�p�����E � ���Lс.O  �'�1��y�������;���ʢE�^\�lYOUU�  `&�uww�_�x1A  Z����{�G ����ˇ~(   <�����3`.�e�w��0���j�
w Џ����dIH�z,  :QM�.]`������nwmnn��N�s�SO=u��>  ̬���q۶m�����===�[�F|>�tuu�Ϋ����� �����>��������7���� @?bv:� �՚���l�LTp��_\\��lo������> �����6n���?���@    =���'O�������9s�  �~�B�9�P��io =eee��p @?����Gbb�����9��w�V�Ͼ򕯼�t��A  �k׮�=��= h���p�VT�;  UH4888�|���B�qqq(c���p��0�����X �%>>��ӌwh%--M  �^Ԕ��h�v��Ž.����x5x�o˖-���ա�/���  �?�����j���pႹO" ����@'���  �k```��}}}�1w�̺���<�� ����U �����C!&  ��1\ff�����tqq�

�����_SS#  ��***Z׮]{_GG�/{zz�}"	 ���*---̎
m̙3't-I�� ��P��			S�pOII��rF�!w�Դ���W�p ��pr:��  h���ޒ����r]���UV���C�UZ,���o�-  `�***^{��G�����^M	 0?��x�bt��`srr���I  @x���R!y`���ޮp ���V�  @?���Z�
;

~�������ݻww?~<����R  ��<��V�^������ `z^���;����O� �0����jp�_�}ժU	~�?U Fgg�U�	��~233����㙞
  Mp7?��6��x���edd<u����   �SXX����� 0���z����ŀ�v�=zT  @xLG��
ɳ��a������������io�w ���:4� �O�����%---0w���G�n��۷o�2  Y?�p��M������o���\M ��鑳gϊ��@s��  >��ந���D���8�]o�3�	��QM�E  z1{ <��;  ZR�vr�����N�����[\\\�hѢ�-[�SUU%  `��ر�oذa{MM�V՚ 0/��K��P�   |�+ச�	�c��b�~�}pp0�p,`,��~���%!!A�,==]  �~h�6����~��]����z~~�S���;SWW'   ��޽{��ի�T__�  LK���.t���+   |���rF��w�����<&� �IKK3KMMUS	  Џ��Czz���v�l6�[����<�MMM  �_OO���̙�x���, �ҙ3g�����e9�����M0+   ᡚף�s`�Ȯ"��ǚw 2��=66V  z�={����  ��襦-))i����j����o|��.]ʕc  ����ߴi����~���N� ���'OJii� f���YYYr��y  �o���4�c�Ѳ�4�&���y�1� ���322  艀{􈉉����^��u��p�j�۟)++�p�ر����J  Ƶcǎ�͛7?z�ĉ]���9���p�6rss	� &j�d P��)��� ��	��
�[��tww_yL� �c�w�]�m�z  06�3+33��r�|���o�ݱcǱ��  �}��ݫW������; `:uuu�B܇� ��Z�����s�CW�{�EV5��qtuu]yL� ����&f���:�  ���DNRR��\�Kv���j��|�С��X��w�  ����~���˗7�={���d.\� �����Prrr  ��j^�����6e���'�@�/����B�!�@?f�gdd  Г*`8w� |bbb������t�>;;����ܹ�����啕�  �b�X�۶m������/_�B LF���|���w  �kx^q*T�PFˮ�vb��;` ���Uí�8 ���ٳŬ� ���/�ucz������������m6۾g�}��i� �p�?�xͣ�>�����G�u� �^/wh!77W  @�LW0��@b�X�f3<�N{; �GM�4�>E�����  ����	�.---��x|6�������G�_SS�   \˓O>�������G}M  ���j�4U��w ���������Ɔnd� c��a��L��uww_y�� �'==]̊�v  ����(�8un��tvy<�w���+KKK_X�zu�   L��ݻ��:d �)�k��x;??_ 3���
�#Q�Y �Iz���5�*&&F���
�~��t��~h{��AY#pU�}ժU	�&Y w ���ٳŬ� �7�㗗���v�ksss_��������l]]�   L��b	�[������Z[[� `
�ŝ�;�Ne'����Y��52�fQ!���������ЍYI��1]wE���{DP���ߟ����w�઀{ooo��8��Վ @/fnp7sx  \����n��g��޲Z�Ͼ��U\�  �w�޺-[�|�������� `|*�~�w`v999܁(6�Tó:�dx�}d ��;>�pW����D���U������L`(4����OII^ �7��'��:�[\\|�n�WY�֗��o��ҥK�c  DDyy��?��#_?q���)  �;u�T(D/����;�褂���}:�~W�����S�k��C� �f��%�;Ze��^y>|a�z����8zzz�<f ����&fdֿ  ?��Յ����^��u"''�&%%�{���/?~<����R   "i�Ν��ʕ+o=u�K  ��s���D 3#�D��ƎE��6o��x~
�o|W7un��Md��!��!��ꪒ���~��w�`hp ��5���.  @o�M!����w�\����7���v���~MM�   D����ۭVk���7 ���p�����
���������3���P������
���t��	�c�*i����{�p�tM� 2���fϞ-fdֿ  ���V���3KJJ��u�n�WY�֗:Ti�X��   D�]�v5=��#��������Hv �����	`v܁�5��k�����h�ۡ��� �P<��=QY���14��%e�wF�2p�< �'99Y����lRRRB'  ���lT�Oaaa����}vv�?عsg����C�+++   ��_~��#����VP� �u��9�|��ig��@�RAV#
Ꭴ������=|��JV��l�T����}����3������� �1��4N� �=�������nwmnn���������?<IK  0��;w�\�z����K `X�����OZ ����
�(���,��'C�+��������C���;����(�[�����#�� �[oooh���; �g���bF���  ����Ĉ���s��=��������g<�oMMM  `6��ɟ���>��ܜ"  C�z��aj*T�_�� �e(���R7�I��
���F0���Ѿ#�OpA�;`���Wp ��5n��>  ?�4��cq�����>x{��o>�z��^  0�'�|�e˖-����랞j���c*dH{,�,''��;e���>*��������C�������M���<�{ =�,i�D��:�`===W� �1c<%%eڦ�  ������~��]����zFF�S<�B�K/�$   �(//cӦM;N�8�(��x:::����<���X���C����Z�Gk�V���л�� �B�@$M���w(�lp�@t����4 �3����   �����~��u&//�����~��?���h�  �؎;6�Y��+uuu� ����� ���~ч��Ԩ��7��q��}�Mᙱ�0� ��|��Հ�z����|d"��;` ��4��~f͚%f���.   3pOLL����Kv���j��\RR�rYY�_   0*��y[WWWS��� ��Ԍd��~� fe�Z@t!�>*�����4��>��}�����>����������! �����cv8 @?f����  LLgg����E쿧�@���z


���������=���?.   ���~�{ӦM_moo���Uk ` 'O���-f��I�'m��Վ=Z۶jvW��U�}x���=p-�c��<i�0��jG��d @/��~rr���
�g  ��H��gff�].��f��������?��{^�W   09;v��ߛ6mz��>��j �
%�:uJ����QVV� �.���1s����w�Gv�'�e����APjYYY����W�V�J����* 2pg� �G�������  ��7ퟙ��(��ŗ�v{��j}����ХK�   �gǎ�_�z������
 �0jkk	�ô222@�P�akC��T��H*�0v��>�����\�xqV�>4����($� �����p ���s�IOO  ��hpW'���N�ﳳ���j�>�q��q  @�����1g��ٳg� 0���:�*��g�^�������Žx�$���O�23덛�U���R�&vڦ�vf�IӝM��Ĳ%�-��(R�\�i�N'u�qֻ�$Rwf���ݤʦ�e˔�IH$A��$J .� q���6`�� ���|f���H���?��;W\Q.s��3gGߧ������d�����>{
<�"pg%��̬��� ��	� �����w  Zj�~����۷�^{�v�5���?��?8�"= ����<}�}�}�R�|gxx���8y�d�&��q��o����g���l�S�����9q�|������k�O�:/'�;Qm0��)f�;@~e-p��=��m ���k֬�}�{�{����/�������_�� h�Gy������^z��}���C�x�����Ȣ+��R�	!pϷx���E�q�{��b307�]��|�}�_#q?���W�u0?��t�O�@��Mp�Sȟ��k�z� �}
����͛�j���O�l��/{zz�  ���#�<~�m��boo�� ��W_��Y1p�A�΅T���v��}.v?;z�!����77�9��5��̷b����=�d|��a�;@~e�Q�w `Ή'�?_�~�����{����?��<���}�x�* @�}�K_�����O���_ H��CV	�!9�,E��7)<s���禾��k�V�r��Ԭ��d>p�V�kLp����v�)��W\�$k�= �Ҽ��[a۶m�?����ߵ����}���'O  ҧP(T�뮏�]��{CCCƯ$X�R	o��f���$�=]]]H��EʰTs�������{���������011Q��0Y�������O��i77�}�n4 �%K�[[[Csss  �'.T;v�>).Nf7�x��>���  ���/|����������`
@��ss�;Yt�UW�����6��R�V�[�q�׾��b�=>>^ާ����\��5�xw�[�}���=�5�H�����v�|����5k�@^����ǘ=^8���{��&���  [>������o�����d  ��y�>�� Ys�W����J#�/���]ggg};W��b����܏�:=�M��
�����j��&N��!�9	��'�������@������G������/����*1 @=�����O��v\�! �HG��Ǉ�R)@���� p�b��---��܁�qx�ܔ��#��s�x��r���=�A˜k��^{A�@j���_�X,���@�ą������8��ĉ�g���p   s
���g>��[����ӧ� �3w>�e˖ Y������{Lc,�4�[���շs��v��b�>����y�ZY�7�į[s���{��pV�$�	� �����ǲ4� �(N����1j��ڗz��T*�  Ȥ������{~}ll�O;E�����dM��[.��-r��wa5��s�ù�C�v�}�v������g�Jܼ�����7�=�=�U��g�;@~uvv�����- �3888��m�&��U;.  d֣�>����sϧ^|�� H�x���O|"@���Pq��o�����1"���R�V[�����R�bq�kn�{��"��y�n�Z�)���à����w����)"pȯ,�kָ� �`ll,>|x>h?}���>SSSG  ��裏�������L__��D9~�x}@PD�\y�wh��ĔgX��7"p������kߙ���������q%b�˵7��!&�j����wH���=i߀Xyw `���þ��z������2'&&^  d�ڵk?x�UWy뭷Z ������{��dI܁���H1pokki��ƛ�nݺw�Z��ώ�禾Ǐ�q�|V����|���Mp���܋�b  _����(. �q�1{��:T_]mMMM�_   �y�����0<<�֎;�Ĉ�w�F��%V��q�c���=�"�kFΞ�?���\c�RV"p�7%�k�܍τ�߀�7��� �%+�{��ؓH �qFFF�ѣG��J���?O�\�}�'�  ȅ�����Ν;����?��FM����:dMWWW G�N#�%�nii�o��V���>�ǟ[�8}%���n�s띁�o��o�k��`>p :::B�Y��J XMq�رc��qR���@HRH��ښ�1*  ,Ȟ={n������? H�ӧO���~��k2媫�
@��i����b$���\�Q��c�>7�}��Z��=�_����@.5��o�F���M�����+��(��;@~��e�D�; ���ǈ=��1j���K�Bnss�H   w���?x�5�{��7�1� �:���,�z��Z� "/ܗ�\.׷���w�|��47�}.x��x�ߧ���p��E����Z�v U� ������Gc �oppp>h��c&ӢT*�  ȝG}tp�Ν�222�g���B ����O��OȊ�k��qΜ1�����[�B�ZZZ�۹���������=��YNnLȷ���ȁz�^{1t,�XY1pw�@���Gea�_*���, `q�a8p�@}��{��  �Ҟ={��w��Ń�/��X��/�k��*����Eྼ��aʸ҃}�r�>��t���CV&��pqߟ�-$���'O����~�ȑ�\����  ����Żn��z{{�z ���4��Ǐ��7�O����h^����o�b�#~,���4H��������/Y��I� ��������YT��:  ȵ�7~httt�fm �������hmm�?!9V�H�F�L����@~����0p���5�Rd��) �/w Ⱦ����d��:t(T*���b�?  r���o����v��k��� @�ě��g6@V�)�o��V V���F�L�8�7�.
���}�������b�h�CY	�;;�_	 s��j___=h��B��i�ܓ���
  ��c�=��{���^z��Y�/��������� Y p���h&��S\���r�ȥzT47��# �w���)�{��} ��x�p���z����/򷷷O?��3  j}�ў�o���C�}0 ��j5>|8�ȏ�H�,�tah�3w�k0�����	���;�w���B�'d @ތ����G�փ�����e!  �Ú5k>v��ן<~��U����w���)h��sMh,�{z���YhdX����s��	�"w��jmmi'�@����(�x!���^'N�\X�T  p����3<���V*�熇�]h���Ya�;�����h$�{z�����X�
� ��� ����Cڙ�@�E���������i�&�,\�P8  �?����wߝ/��җ_��S�N������� �\�����$���B�>q�;�t�wc4!E� ����/œ�,D� ��sA{�&&&KS�V�  ��#�<�{��v�'{{{. �����O��OH��k�`u��LRě-J�R ]�Cr�޴�ߵ�B�# ��N��SkkkH���NwF�Zccc�����A��ӧ�cbb�P  ������6�>�� ���"p'Lp��'N%)bk'pO����k���� � ���	�1p���V���ɓ�������a`` X?Y�B��  .੧����������˧O�V% ��8�=��^C�	�a��SI
��t�Ǡq��N2���^J#H�;@~����4��t�����q:١C����T`e��p�7�e  ������}��n�����q������u�H�5k�`u9n')��K'�O���?�k:��|��QZZZB���@Ҍ����G�փ����044X]mmmgzzz�� pI?���v�m�v��� ���k&w�N��kn�2$��=��Gr�>=�t��t��S���Ӵ��~�'��~q�ñc��A{��'�Ņv�v�3  `�~��~�?��O�9rdc `U�5��~����&X]�b�D$�^��d�;��7@>����4���G� ��b�#�x!6F�}}}��T*  X�r���u����>}�9 ���zJ���l�Kzutt���&�#���$�}z���S�P�CZ�q�Sw X����A��Ç���X �
��  �K_�ұ]�v�ڋ/�������x}�ȑ#��}o���C�b�^�T���$��.��K�ivv��{{ R�Z����Cw 8�����׃���8q"�*}  i���O�w�}_{�~= ��⺋���[�f��V���$I���]n՛���=ݵ����� ���_q� �C<'���'���I����W  ,�#�<�~�w�CG�� XQq�.�����$n�H/���j��S:�  $WKKKH�xcV{���t����A{ooo���dÙ3g�K  �%Z�f͇����#�N�r�`���ahh(�]�6@Z��G�J���+��_����@�|?p��_����/ 5Loȧ���V�����(������sA{��J���0==�  ��Gy�������J��NMMY�XA�?�c? ��:�W=u�$q�E�MOO�󧥧��Xڼys���x �!N)�S�w �������W�������T����e��'�	  p�����x�����[�G ���f#p'�:::����$�	��f��OCCC-���q�� �����o1n�@�?mmmNr X?��gjnz���� ���Oً7�FZ��J�`5X�'i��f��O��ڛ���~H���� @>�9p��G ����p�������:�!>R�t  �e������y��7�x�xV�0::^���~�� i�����'F%i�&���/�b�^*�˭�j5 �� �v��(Nrioo ����T�������)_0����   ��{��뮻>U�T�bbb�xa����I+�;�1*Ic�{����Ssssk�Z�z���ؘ���UKKKH���N�+ȉ�ǈ=��1j���-:q	�  ����������_~��;�`���χ?�� i$p��!p'i\�J����@�
��z�^,�����|jnniw �kppp>h����SSS�  ��c�=v�m���s���? XVq�AK�R������4^����O�m/555��^ �!ȯ�����$sA{�N�>`�Μ9�   +`�ڵ���>900�6 �lb�#�m۶H���� ���jI�t��}�,��uo-��	@jLLL �\.�4��[�Z'O���ڏ9R�9X���  `���LԶ��T*�ett���Q\'��F���XY1B���L?�{����R�^�$ �w��(ȯ����F�gppp>h�������[[[��W��  �����g��]����S$�O\3�����	���$��M駙̟�����V:�ccc��jnni�|w�$���h}2�\�>44`�Վ<� ���/|a�����:�� ���O�	���Ҥ��- +K�N	��Ͼ%�{�7H���� @>555�4>u��v�d���ǎ��qR���@p�;�����t  �U�f͚����\ �lq)�)�����&wXy"T�(�ĭP(����)���X� Lpȯ4No�LoH��h#�x�1F�}}}�i�B��f  �U���3�{����n
 \6�;id0�<�H�H{�|zٷ�O}�{�w�@:�򫥥%���B�Ɖ������v>A����   �d׮]/ֶ�=������7���(��J��'&����.���/8�&���j ���S��w�!�t� �W\lK���� �ꘚ�
������q�։'$Y�5�Z  �U�{��߿��>����� �e�T*�ԩS�k�	�&���wX!T������?�B����
w��J����� �ʈ7��c��9r��	Rejjj  �U����7n�?v��� �e�kRw�&>}xxx8 �O�J����nq���A��Z�}��Mp�t��W'���b� X>����A{�&&&�� �c  �U��SO����|ddd��9V�� $�O}��&q�;�2Lp'����1ilgX��	��H�x#���d  ����w���� �<�&�Ç��O��---�?��?�  � ===�������U���'
��h�T
��>+Ǳ5I&pO�8�]�������_qH��x�@~�1p��X������W�������dRkk��  �P===t�w��W^y�o �djj*;v,lݺ5@Z�~+G�N��8�t��ɗ��ٲ�Rb||< �_---!mLpX����z���C��/B֕��J  ��'�����|�3}�s���%��Zw��wX9�S������ɝr)V�B! �&pȷ4>fI�p~###��ѣ�A{���%J�қ  ���������`��� q����D����ʈ񰀘$��L?S��X,��i166 ȯ����&��TN�X	q"{�b_�h500� �j�  �����C=��?���O���LX�'Nԯe���H���� ,?��I:qt����N�+w�!�� ����=No��  ��9v��c���8�ݢ�S�Z}-  @B<�����Ν;���� X��v������/@��+CxJҙ��~���K�<�wH�;@��J��&1pȓ�����=~����#/  H�={��Ƨ?��9rd[ `Q⚘���(�eR��$��=��gr�\���MW-9%pȷb��ģH������O�:p�@=h��;�(�!  @�477�ꫯ�;u�Ѯ �wH��=5�BxJ�	��/~㖶~�%���B��d3 �Ҷ�f�;�5q���ɓ�Sڏ9b!����y��'�8   a��S�v���J��簾�\@X�ӧO���z+\u�U��wX333��u�l���{>
�R���.��� �&''�\������dA��>����֏ˁ������ @b�޽���ڵ�}�����k� ���V�	�$��l��������R�Wnll, �oi��O&���@ڌ���'�ǋq�
�J% ˯v�0   �v���ٚ�j�� ,H��?���.mC� bp*&�F����\)�b��D������v -�4����z�/�X܂UP*�N  H����hdd��믿� ����V�VC�X�d����3��4��)���M���i0>> �7�;���z��c�/�Ÿ�"��b�x<  @��s�=C���/V*��/ .jjj*?~<lܸ1@����ϵ����l0�=W�w �������	G�����h�3g�	  �{�����;w~��矿[piqN�Nҙ��O�N����\)�
�Bɂ$���X  ���H���� �(qRT�bZ��~�ĉ $�����  RbϞ=��~��7:t�' ���>��H2�a�	�I�l6�s��v�&B�	�H�b[{{{ X-q1j``��Ǩ=Nk���V�V�S  ������N�<�& �.�ɮ7�pC���$�	���=�or�^J9r��������w`���q���@:����'�x�  R��_����ݻo����hz��B�Sgׯ__�ڷm��lْ�'ђo%�aY�h��!ҠZ����&W�wH�x����T  ���Ǹ�P(��o�<|��|�~��� �S�X�	.  ��k׮};w������? �������۷���� i$p��%6%-��eC�:ƛ�\���ݑ$��� Di	�����劋�������I�� #ZZZF  �Ԟ={���;�W^�H ȸ����d���}�ڵ��\6�S�	i�Zcv�k� p�� ������- ,���`=f��:�)F�Q�R�   )�}��O?~�� �!1�ݸqc=h��ڻ��=��L�����q��w��s��vg$�`&�	܁�	G���+�J ��vL3   �n���ݻwlxxx�\6�v ����ǘ=F�6m�7��:�sX^w�����ɍb�v�R���2��(-�{{{{ 8����p�رz�'�XH����9   �v����C=t�s�=����8�����ڷn�jM�\�����&�g����(�fggMp�3����w eb�#��Ǩ����"'ov9   |��~�]w���/�� ����Æ�A{ۯ�� yW.��|\�!-���{n�m�� $�	� Di܋�b}�ȯ���������n��evv�?  Ȉڹ�/mܸ���cǮ 	��ׯ_??�}˖-��~�wX>q"��ؤ��=;�Q�Mp�����y�)����T����o��f ��x�^���  2⩧��ٹs�G���^�T*j9�!������۷���� \�	�|LoA���!��]��|K�t���� d[<>=y�����#G���,X{{��O<a� �Lٳgϡ��?~����#��:::�����k�`��|D���	����;7Lp�$�q�`���C6���arr2 ,Ess�H  �ڹs��z��w��^z���eV*�¦M��A{����ݝ���BRŧ�Cd
4��27�&�C���� H�;d���h}2�\�>44 �Css��  2����[o��p͖ pb�#��Ǩ=��1r�G|rr��M���'p!�q"��>3� p���&wH������W�������VD�P  �aW^y�N�>}xpp�9 ,Bgggؼys=h߱cG���ʱ�C�N���gK�Q�M��W���6H����  i!p��x�7����Q{��-@��P(  �a==='v���k###ONOO�inn6l��qR�u�]  m\_E��E�!�Lp -�岓H����p���z������ ��&&&  ȸݻw?�s�ί�߿��(
�����Ǩ=Nkojj
 �V1.5�4�z͖�"�
&�C���@Z���255����A�k��N�8 mzz�[  r`Ϟ=��g>���ɷ ���������� �
�ہF��	�d&��wh�8q```��Ǩ=NkwR$I�X7�x�_  ȉR��3W_}uߩS�,�AN�����[����֭ �Uw���lq-<Lp�$3��(>�4�ZZZ�����MLL��jkk;���3   '��S�v��{�J��OMM%�X�R�6m�T�������T���r��T�V�g�;$��Ԕ�A RãUa�ś��O�> Ңv�0   gv����>��C_�����9�!����1��;�a{�� �4M@#���E�!���� ����_����ɓ������رc��V�\  �C>����~�/:t�@�tvv�͛7�c�o�1�Y�&  �R��u�l�ʅ�	�Pw �D��cppp~J{ooo��� YP*�N  ȩ-[�|hhh��o���Dknn6l��qR{www(����P�w���`�;$���4����⍎��#G���CCC ��  ȩ[o��r��������wm$��1b�1{�������  \���42�=[�rA�I5>>  ��vl`a���ñc��A{��>00`1ȅ����   9�w�ޯ������ ����5�Ǐmmm X8�ہF�V����Z�L+��Hw �"���œ��ǘ=F�}}}��\����  �s{����;����?�U����n�Z��nݺ  ,�k]@���ӗ�M�	566  ZZZ�C����A��Ç��W,�,�"   ����6l���W��
���ׯ�Og߱cGظq�Ɏ ����왙��g��J@Z�ɻ������_�c�~�ĉ ���������H   BOO���ݻ?>88�����b �EWWW=h�ڷo�n�����U`��@���l�Cŝ���d �4hmm�'q�{```~J��#G�?��j�
�� ���ڵk�����/�������3l޼y>h_�vm  V���42�={��'p� �w�`ppp>h���u3"�"477  ���������^~������rظqc=h��ڻ��EJ � q��O��c��/�>�;$�ؘ�v ����,�Of�ڇ�� K����z   �e۶m7U*���Ǐ_�w�R��c���M�6�RI�  �fz;�&�g�3@H �; i��� ��b\___=h����G�,�B��  �w��[����/~xxx�{�J�)@�uuu��[�n��� HA)�&�g��H�@Z����EZ�c�W^y����	��155�  ���;^y����o��_�7qxʆ;�[��ds=���5d��=��@w Ζ���CZ�����G�֧�:t(T*� �ʛ���  �z����=���+/�����a�b1�_�~~J��-[�? ���H
7�g��h||< ��$�---�jjj*���׃�8�}`` ��� VW�x�?  �^}��Onܸ��رc�dH��>�o߾ݚ2 �����2�={�&�g��H���b�̓8����$�Wb�c���i���h�����W��  pQO=��LOO�G���^�T*��Z���1h���Ú5k@��kn����	܁��d��H�x"%p�\��<��{kkk�F���G�Q ����2  �����}��G�����M8DZ���q��z�'�www��	$�ﱰt�D��0�=��0v� �K\,�
�F��j���A{�H�����   ,�=����w�}��^��$P��c�c��oڴ)�J� =�t�?���0�'�p;�$�dy8ӄ�1u��I�b����OHO�<9�9r�̀ )����z   �G��[o���Ço� �����}ǎ�����- ����T �����g��=��0cc����%5�mnn���T������7LNN ҩX,  ��]��z���n	�����Q{گ�� �]X���q�$��%O��._YH�; ���=^�p�3�att�>�=�
�J% ���ӯ  `����===�6<<�T�:�J�������=F�[�l1�,�;,��i�mȦj��߳L�	#p�|��X��bxK/�;v���I�avv6 �=�}�  X������C��g�}�7,������}����{��p�,��;)��l�g��F���$�\.X��ǈ=��1j��� �qJm��   ,ك>�[���g?�ꫯ��2ttt�'���k׮ y��,M��733 �Lp�&��l�C�� 8W�M��bFFF�ѣGÁ���� �Pkkk��_��   \�ڱ�߸�꫏�:u�-��J��iӦz�'�www�z �	�T�z�'2�f����j�{�	�!a�_ �O�I��ι�?�{������z+ �o���  �l�>��`OOϯT*��gjjJ��uuu�;vԷ����w:c�;,��iW,�3c�{�9���w
�[��I�]�&�s�'N�}�� �j�
C  X===�s�����O����ΰy����������+� \�&�F�Nڙ��MU�3M�	266 �|��`����l۷o 0�T*�  �e�gϞ[o����:t�G��d7l�P�o��p�u� G�KsF�Nʙ��M�l�C����$��9W|r� 
��   ,�;v|�R��|��׍�΁8e�����Ǩ=Nkojj
 ,�H��{��3�=�fff�%p� p>I<(�s>�B۳�> `vv��   ,�[n�e������J�����
��$������ ��H�fFDJ�	ܳ�j�{�	�!ALp�B��`P.��K������  ��>���}�ػ�������tkoo[�n��׭[ X9���X�x�9#p'��bC~�5k���?��Oܜ�-/��&p��p!I[0���������R��D�����  ��x�����;��W^��@�İfÆaǎ�����nk� �H����dA���;;;�}Ŝ8q|jj���(���&~_:ܳM�	"p�B�vP~�	�->2��������jii�}�'  `�lܸ�###'�����N����z�'�o߾=�3 C���}C4j����G�s�k�q;�\�~v ?����7Ŀ�F}}YYwH�; ��E�;/�	�򭭭m2   +��[o�ܻw���u5?A��͛7׃�o�1�Y�& �&�������྘a��R�����ǹ��?$p�.�;$���G �|�vG�	C\L�p�W�W��jmm�  `������ٳ��g�y�qaC���8Q��.�?tww7,��℺�x�7dAR&�/E���!�qkooǯŖ���}n���v9��I&�;$����;� �����\H��O�ݼ�_�R��   ���;w~鮻���_~�c�U���ǘ=F�6m�OZ ��uaѼoȂ4Lp_�����v����!�����{���g-�
�3�Y6$���X �Iڢ�	�\L<�޲eK8x�`  �j��  �j�m�vs�R8~��U����5�Ǐmmm��q�8g�d@�'�/E�����/���υ�g��i�+p�.�;$�������Ib�;�/�	��kff�p   V�-��2���pxx��J���l1`?;h��; �'p�ŉOOc�
��[�~1��"N|?w�{c�s����/H���=��w .&�0$�	�\J��@~MNN�  �U���}��޽{��}����$�I#�����G��	���` X9X8���
��J��v���qv�>7�=	S߫���CB��� ���M�hnnp1�y�{�ڵk���P  Μ9��   ��������{������_\R��>�o߾�`��f��q���_���;���������������	�*p�,�;$�	� \L�&���� ��u�����~7 �/��ٯ}�k�  �!ZZZ>�y��cG��.����sA{� @��aqLp'+������!���������������c�n9�^����CB�����ɐ1n/
.%^(��O{{{��� �����>���|�R���zp\�ܸqc}�*Nj��	�swX�;Ya����^��|/4�=>5"��Q�gV�4 I�Dp1�@>)�#�`!�E�xҺ�P ҭ��u8   ����w������i����#��.��M�6�'	��aq����{�,f���v��K���l N嵣�b�c���|w���tvv����=���_ �G�T:  �������ܹs��ۿ�����5�oݺ5>U* ��LLL`��4eȂ��������Ź����w97�=64sề{�%p� p1I
�M<b1�E�;@�ԎN   ����>����䫯�zCȈ���6�םb�~�u� X(�a�bD*%+LpO��5��qscs>�� ��� \L|�GR���b�����7 �1;;�Z   �}�{�O�>}����j	)#�����Oi߲eK�� �O�wȊF�C�'!4j�<����� \J��7nI�pc�;�/8�׌0�����8  ��������{zz~�R�<ߞ]]]�A����CKK*�| hbb" ��Y���<�wX<u$�������
�����c��΢ĸ}�ƍ�������/  H����������|�;�����>(a.h_�vm ��o�St����%�&w`�� w brr2��	�,V�0)pȇ8��R�|3   ���C��g?�ٛ^}���6���7m�T_7��ڻ��C�P ����8n!K9A}vv6 ��N� p)q�{���b���� Ⱦ����?��?v�  jݺu�ꫯ>q�ԩ���}c�#��ǵ����j�f���NV��F�Pk�;,�UH w	��I pg���������� @�����   �zzzN����J�����V������7o��;v�� I�'N��NV�ņ��&���ܡ��ݎI	H6�I�x7��-[/� ȶ����  �h��{�?��C���g��m9�����aÆ��=Nj��� $����v��с�	�4wh0��X���ɐ�R��w��+�  H�|��;��x�R�q�A|r_����O�����  ���pw����)wXu4�;�X��,"�Y�x���+
G  �
���?844t��s��LWW�|�����  i111��9#p'C����`��I�`�`��0��\.X�u�օ���:�:u* �]333  �
���>��c��|���oLLL���ioo[�n��� ����pw���C�Lp���C�	�X����F����\�8�K��m����  �w�}�7~������{0N���6m���q-���;>�) @�3`��dI�'��aiJ�`N� X�$�&�s9��g�y& �M�b1l߾��  @j�������o����t�Wn�q�! d���D fff&@V4:p�7�gu�#� X(�;ig�Gw�dSGG�tOOO�X  ��z��=s��Gk����s��R���?��?  ���0�Z��ydI�o��~���C���� X�$,�	ܹ---���ǎ dOm?�  h���333?S����MOO�x�c! @Ό����Μ9 KLp�t�C�o^��� "	�{�㉹L۷o�dTKK��  h�'�|�i۶m?V(�A���L���  ��Mp���5��Mp��Q(AŻ�ݡ�BMLL4��`�;��nO?�t  {J��@   b߾}7�ś���� �w
��	�ɚF����ܡ���b$�����˵aÆ8��Sl 2�P(	  ��x��;'''?P��S?ض ࢆ��piw��������C��X�$|�h��ͤ_�X[�l	 d˙3g  `E<��ӥ5k����	퓓��}4� A�#p'k���K�P� �Pq�u<�p��Y۷o�d�����   ,�}���P,o�A���mm  ��R���fffdI�	�J
%h �; ���wtt4��o��p�7 �%ހ7==�  X�g�yf}SS�\�~sm�.  �"�IxZ2$]��.�%k�0ȯ��!��΅��Xw��ꫯ�֭�O� dC[[ۙ?��?	  ��}��hkmm�P�ӛ~��xm+ `����]���C�$�s���	ܡ�� ,V�'K4	�Y&q��w�� @6���9� ���w���j�������õ�5  +.���	�ɢ$tn����C�{� �411���?	��"�m�&pȐr�<  �wy�g�׎�?R������OV��� �ꆇ�pi333�&	������\ȩ��I� ,Z�o���,�K���y��(��'  ����133�3������? ���0&��EwH�ƿs!���<���kd����v�mmma���a``  �~�ㄣ  r��'�lڶmۏ
�z�>33�����  $J�R	��	��"�;�S�߹�Sw �bbb�a����������̙3�  �ľ}�n(�7�E�+  �f�;\ZpgffdM�j���i�;r��xH/�ɒ���_ ������   ��o}���柫}z������>n	 @����Lo'�����"p`)���I�mӦM�\.���� @�U�տ  �O?�ti͚5�	�����8 )644����E�s���5��a�;,��h����  �����X,XNq1a��͡��7 �^���3_��W�  �b���X,���jۚ  d�	�piw�()��fgg�8�x�B	�X�F�MMM��7� pH���v�(  u�����j���ڧ7������Ǎ �,�;\���,�Cz%��9$p`)&&&�{�Y	۶m �[ss��   	��϶���>��o��������?� X�J% W;F�5wH�d�{!g��SSS +� O|
�տ���?���k����add$ �N�r��   	3;;[|��~�P(�\�Vo�}�q{K  r�w�4�ɢ��R+�^���X�j������U��Mpg%ě5����� ҩ�/?   �}������~�����O]ըa @r���v���u�A֔���_�xwh����  K��4"p/�V�7� pH���ك  `���333?S���l?a* p����P;f����NV�<�R˻�w .G�>�v��U�}���R��8I�h�t�^  �U��O6m۶��
�B=h����h���O�  R��v�4�;Y����wX�d�{!gLp�r�)����`%\q��ꫯo��f  ]�J�j�/  ��}���P,o�A�~sm[  �R����dURw��`��1���Ѩ)wVR��.pH�����W���c  �ɳ�>{uSS���>�ivv�j7 �����o���d���+�^���w�(����7 ����>  �2<��ӥ5k���ڧ�*
��}�볳��  �L�piw��\.�$���	ܡLp�r�ɢ���� �u�����]r�1y3Il�,i�$BYH�
�BxJy <m @�m����L)��I�C��v��]6���v�ɰS��3�n�]�¶�d)v;~�eY~���I��s�"�m�/z�W����̜�7�t��s�9���/[�l��y'� �����x  �4���u
�����4�����U P&w�����Z$p���C�MLLĹs�0swjQSSS,]�4�����hll<  p�ׯ��(=MA�GJ�o~����� ���py)n�R��]w����� fj��B��ДWgg�� c���  ~J[�Px_�iW�����YzT� �B��g�ej���K�v�̙ ��8}���|]�;�bŊx��쨫��  �^�X,�]������ɠ�����5 @���	ܩe���'p�
�0[)pO��T:8�Sn7�xc���y��!��% �\����(
])j_�n�/�.  ��ѣG�4�;���w�,�;T�ٳg f#�� x����uuV������-���6m
 ������ @.���Ο?�2~2�=m�
 �*7>>Ǐ���Ԫt����:Y�;L_u��B���'O��x�n�;����)pȈ����w��m @M���/�ߞ&�����������c� ����ied���Ԫj�ޞ�a��Pai�. ���ӧ+�5Mp��� ����v.  �)/�������ݗ�b�xo�*;a `����k\Z�n�JP��)p�O�&p`.�	�f�;�p��W��ŋ''� P�ZZZN  ��v��7����[z�U,��xK�s�� �Z!p��3��Z�����q6L��*��ٳ �5ܡR:;;���? �nMMM� �LY�zukKK�ݥ�]�ow�ES ��%p���S˪i����O�t��9o��N���׫����;@6
�= @�����(�w몫�KS��/��U �V����U���'p�2������?>y�t��1N ̙J�uuu����1�=�.v��V�]�=  �:�ׯ��(=MA�GK�K��;�x ��1�.ϠNjY�	�iw�it������]� ����Z���K�.�={�f.\�  ̻����B���Ӯ��������d @ɑ#G�4�;����&���P{S'p�8w����Ȟ��M�7| TR������JJS�� ����� �������켽��n2h/m�/m� ��H]piz'jY������
�q̞S�>:: 0�Μ9Q(jQggg���? �Sccc��  *�����P(t���}q  pE�� ..]oNԪ����&&�������==�?> �ڤ��/X��"_OHO��t�M�'�XP������ (�W_}u����W��~��my  0-���i� .��vj]�MpO�0uwr�c���?��8y����U__˖-��[� է���D  0gV�Zհp���ޘ�~���{J��u%  cRb:5\���ZW�܁����Y�+7���1Ĝ8�Z< �v���}-�d1:;;� U���q$  ������B���z���Ҷ(  �3G�	���Ժj܁��Ss�����T���̙3 ��ԩS�Z&�3:::����а7  �����_w��b�x_��vc  P6�.M�N��C�	�ɴ��1�������l`>�}`�ܙ�^{m,Z����� LMCCÎ  �V�^����rw�i���566��ңe�  *dd�"�p9wjYj�+�-�L]u��e�_�)nJ �1�'O���ܪd�[W��+�c������/ �elllc  �3���:>V,(��?/m- ��8t�P �6>>P�Lo���S�R�������>11 �O��Nttt��йs�� �X�f������/=�z=j��` ��p��� ..��]�ew�>�;�.E�N���4�8q�b_�w�Kgg����l գ��>�� @����������흥cV'N  ��	�pi.\�ew�>�;u���i�� L��ӧcll,���Lpg�,X� ���ZSV �H�w��s�=�@ ȅ�����������&������]% � �;\���Z'p���Sv)`߽{�� �X�q,Mq��kjY��.p�---� �����u
��7��Ҷ8  Ȕ���O_.N�N����ݪ�0=w�.Mj߱cG  s/���S�R�z�� �:477� @������C��]�b�å�e @���9BB�4�;���w�<�;e��� @y�	�P�-[N�T����} �a�V�jX�p�m�hB���b�53 �r�С .�u7j�����:��� ��Ҋ�A��o�� �_�P�  ����Qz��z��˥ma  P��w����������E+����)�&�; ���������T����� P����������X,����M @n���&n'4��}wʮ��9 ����)p�_�� ��ĉ/ @�Y�zukKK�ݥ�iB{����;K�u @.���v��Z'p���SvigQWWg� (�'N��7����q��� `�
���[�>  �Y�X,�[��uuu�MLL�Wz|_�M� `�	�piw�w�$L����Kq{ccc��� 0�R�;666��-��?�����/_6l �ςƞ|�I� ��X�nݲ��}������J�פ���[  ��>��	ܩu�<A�	�yw*���Y� e�.�)��\sM@�����̳��Ki  300�>>>���Ӯ���w  \A�S�;��	ܩu)nw3<d����H��ɓ' �{Ǐ��)p`~���	 �2���/��^WW7������h�  �r����!Q��	ܩu�U�O�NEX� �'Mp/7'��-�%K����H 0?� �����(
]�G�����  f!���MLLLnP��P�T�� �'Mp/7�wQ-:::� ���`W  �B�������v����  ̡C�pq���---d����pW �ϱc�򢳳3֬Y ̛� 0����ZN�:�k�ϟ��?��?����Q,  e"p�K��ZE�w*�N ʧܡZ,_�<
�����ɓ'_ �+x���9v���������ui�=���p_��㦛n
  (��pqw򠩩)���Sw (�'N�Ez_�t�� *+�`t��� �O�7���ܺk׮/<x��m۶���g��������;  e'p�K�uZE�w*�]Q P>gΜ����hllȃ+V��A[[���/��T  ���SO-ܲe�C�c�O����ݿ[8�H"��ԧ  �����\�	���j������ ��)�i�j,Y�$ :::bժU@e����  ���b�_������ݽ{��_��׮;}z�o���'����  ������رc\���<hii�jTWW��	ܩ�; ��k��&p'7���7O��L'������� ȍ���CCC�9<<�u�u�-;t�Pa��y���x��W��xG  @9�ݻwr8���~>��"��;�v�$o� �<R�yQ(b���y�� �r� P������iǎ�>|�W�����G�Gm�8����#p �l����ř�N�k��X�~�������ܹs �=�;y���)p������  jF��>�k;v����ݻ��g�g�FGG��uS���/})  ��w������P;�T�� �G�N�ttt �U,�Y �;��;w9r�����]�������B��7�_�>N�>���  sM��&p'�9pOC����S1---q���  �^��r,I��dɒ����رc@e�={v  �Ly��'o޳g����?�s��_xꩧ���||<M��{�'  `����pqw� 5�@m�S1MMM ��ٳg'���ֲ����D@�IS�׮] �_�*r�ܹ ��}���^�q�Ƈ���?=44t�7��cccQmzzz�  �ž}��8�;yP�܁��S1�
� ��8z���-����)p�������˿< @�y���9v����������-=y�dկw���  0�Ҫ��N�
�g�ռҊZP�Lp��!p�b� ���k�ō7�X��6��j��4Q8����Z[[� P���ov�ر�s۷o��͛7����>[�k׮�ɚ�:� @>���&n'/�9pO׶���S1w (������j�V,����c���@y��� `^<��S�l�����𧇆��x�'�²�}}}�+��+  seϞ=\\-G�T���5C�N��y @y�3p7!�j����ʯ���@  ���]����������޽����ם:u*jMOO�� �9e�;\�����(B��S1&�@y��N���������jll
 �l��w����pף�>��СC��q)pO�
����
 @��ݻ7����w�w*�� �+��0l�;���o���� ʧ�^`K  s�k_�ڛv����ѣGܵk�ۿ��o6�����Ǐ�֭[��[o  �w�4�;yP__�X�~������	� �L����ĉq��W��kO��N�J'(R�}�� �|FGG� 0c�V�jx���?288���������l�u2�]� �\Hײ�����	�Ƀj���I`��TTsss�;w. ��8z�hYw7�Q�:::� e�N�����! �i�������۷����]>��Ç���k���}�s  �u�С�g�@4#�P[�TTډ��|�9˗/���uj�bŊ����� �<J����' ����?��e�6m�����;v�x��ɟ4�a��^~��8{�l���  ��޽{�8��ɋj܁��SQv" P^i�{9� O5���kc��q�ԩ `�� �g|���^�q�Ƈ���?=44t�W��Յ����ԥ_)r�{�  0{��� �2>>�-&�CM�SQ-w (��^{�,�k�;�,���쌁�� `�577 `��?|ϩS�~k߾}�|�k_��ĉ�L�ROO�� �Y+�G��Lp'/Z�PS�T�eF������N������Iss� ����?��Ρ���lӦMo��g]W�c)p ��ڻwo 'p'/Z߅��D,e' �u�������9}]ܩvi�{���� s���~w @N<��s_|�Ň���?=44t���,�����cdd$�,Y  0S{��	��ג-&�CM�SQ&�@y����ѣq�����
ܩvW]u�dq��� `n
�m 5�������������ݽ{��_��W�;u�TP9�\ƚ5k�#�H  �L����m�c�w򢹹9����O�NE��� e�N��u������fi���`�� �!O<�Ļ�4<<���c�-;x�`!�W===w  fl�޽�5�%���[�\H-�6j�������;r�HY^W�N�K�{�" �[� Ȱ�|�;׭^��K۶m��Ν;���F��������;  0c�v�
��Lo'/���j>�P�L����J;�B���Y (�rM�vg?�nٲe����D�jii)��_��� �Y�jU���?�������޽��/~�ם9s&�^�f��;wN޸  �544�ŹnF^���F5���	ܩ�4��� (�r�������j���K�.u"`���� Ȁ����}Ͼ}��0<<����.+�LI+r	� �	�����E����	ܩ8�; �ױc�bll,��uMp'R!p�;mmm� �П��޲y���lpp���O���qk������
  �.�;\���x@���5G�Nť� (�4i}dd$n��9]�v)p������x( �
��_�U{oo�g���?=44t�׿������A�x饗"�7M�s �T��G�	��Lp'/ZMp��#p���L �������,X�ti�6l� �9���8 0��b����?�q���o۶�G}��'N��ܹs��+�Ļ���  ��J�ۭ��~6��E��5��O�Nŵ�� ew���[5��,H'�-[7n f���~[ @�|�[��ܺu�g���?�ַ��m��A����
� ����� .� 3�ڇ�
�a��T�� �/Mp�kN�����w�9R��� P&�=���_|����O����/򫧧'~��;  `��w��Lo'O�=p�O�N�ٙ @�>|x�_S�NV�X�" �Ǐ_ 0G�������?:88��ݻw��/�忼��ɓoشiS;v,����  ���å	�ɋ���hl�� �B �#p��� P~�O��������5�dE
!/^G� f������� ��O<����/w=��c�<�j�411}}}q�}�  L���P 'p'/��#���0=w*�U� 122"p'�:;;���? ��� LSww�����ݼy�6m�����7�R�S���+p `J�9�N�
����E��j�����������u� ��СCq�-����	���;�쵵�� ��U�V5<���ٽ{�o���#�,N+��L���  S�k׮ .M�N^ܡ6	ܙi�"p��J�� dIGG��I�b� �Lcc� �������;��������|p��Ç]�c��߿?v��7�|s  ������jjVT#/ZZZ��	�a��̋�?~< ��9|�𜾞 dI:��t��سgO 03MMM~�0�O��Ooټy����?688������&7�RN===w  �hhh(���:7y����N��'pg^da� Y���
�9y='AȚ4�]�0s���;�\���^�������O����}�9�����x��  .G��fun��w�Mw�E�� �W:i�VLY�x񜼞����������̔�Kl r�X,�����kǎ����~�nqՍy�f͚��.c pqi����p 'p'O�Lp���� �B� �q�С9ܝ!kn��hjj
�&ffll�/ �Y��ַ:w����={��?��z�-[��^@�8}�t���q�m�  \̾}�����pm��H+�777G����9aͼ�@e����[���9y-�ɚ���X�lYlݺ5 ��4-���/ 5����v��ի??88���;w����o�V===w  .i׮]\����Hb��:�;L���y��eA �>|x�^+-�Y���)p���>���nȰ�����~��)fxhhh��>��kN�8������/9  �bJ�9\�����J��&��#pg^�q�T�X �|�2pw�,J�; �W:n? dΓO>���۷yxx��Xv��W�Ȭ���ǩS�ҍw  ?�w���2�&��h3hj���y������8w�\  �s�رHK�766���҉Ț7��M�hѢ8~�x 0u---#@�������;w�L������-�ݨ�{���^�{�'  �	���.#O�Lp��%pgޤ)�w (�����n�a֯%� ��/_/��r 0u���{���z���^xᓛ6mzh׮]�y�G�>}:�V���� �gΜ�pqw�$+�{L���y�v.G� ��:4'�{���Rv�Ț���;�4���o ���?�������?��t�砌�H�;  ���۷O^�.��2�$���L���y��� d]�`q�m���k�Ƚ��> K:;;'O8�0-��y������_��������G�G��˒WCCC�o߾���  ްm۶ .�w��w�]w�� *����s�Z�n�;Y�`�����k��g�֝={v] P���m����[�l�����;�����GGG��5k���?��  �7�ر#�K������[�a��̛��= Y��޹
�-gGV�)�w��)
q�5׼ �Ewww��;~��}fpp�����Ƒ�W��zzz�  �[�n���*p��Y�ӵ`z�̛6�; T���D:t(n��Y���!dU
�W�^ \�UW]5��O0��~��oذ�CCC�?��+�n�ڐ.8W���;ynÅ`  �3g�h����:�@^d�?4��O�μi�@Ť}s����dѲeˢ����� SP:^? �Jww����G�><<��ݻw��_����x
f����e˖�����  ��۷�w�2\#OZ[[#+�0}w�MSS�� *���s�:��dUz�y��7�Ν;��+�	 �eժU�?��G?�{���/\w��� �FOO�� �I۶m��\�%O�4`��t0}w�U�ɜ8q" ��ڿ������dYgg��`
���� W���O�}Æ_غu�G����t��*�I
�y�   �;\���<�J�������'pg^�����FFF&Of�)ֳ!p'�R���������� ?�{����իW?�cǎ�o߾��=�X���P/��r�={6SK� P�� .͹
�$K�;0}w�U
��򛘘�C�ō7�8��qB�,����'��>}: ��B��) �իW�����ܴi�C�v�zϯ�گ->u�T ��n�_�n]��}�  ��̙3q��� .m||< R4����P��#̄��y��� Ԃ�:p7��,K'9�/_6l .mtttm ���?��{������}���'n,G�U���G� �s۶m�b��ť��;y��ìLF���ܙW���I��l��N�uvv
�.#�dݳgOO �ğ���/{��W??<<������}��lL+`�'�  ������4�rɓ,��J��F�μj3� *F�?	���������wN@�h������M�6=�e˖�_��W���P�v��###�dɒ   ��w��\�%O���#+Lp���3������;r�H���Ecc�_#}>d٢E�&c�E ����N@����жm�>[z������Ç�T,���7>�я  �d�;\���<�Rwh�;̌��y����o� �&&&������7�yƯa�M-����\BKK�k�q�<����844t�����e۶m�)�����G� �S�N����\�k���j���y�v6Ǐ �����?��=�!�Ȳ���X�fM 𳚚��@���_��կ���#�����Ν;��Gm�����y	 �|ڱcG�y.O�N�d)p/
L���y���&p�
�����HZ��j���'Ҫ �S�P�V�Z�����dpp�w��w~�w�;q�D ��ȑ#�aӊ+ �|پ}{ �'p'/ҍﭭ��w��;�.KwS@�8p`֯166&p'Ӛ��'W2ؽ{w �O
�MP��~��oذ�CCC�?��#�l׮]�
AN�)�w ��ٶm[ �6>>n�r#����nuV���3�t7 d�k��������4��H�;d]GG���"����
|��߿�^��Ν;?188���{��2 I��o��o  ��V�.-�Y�k�;̌��y�`��  *#ݵ����|��3~Q	� M������ ��JDΜ9�b ̃������n޼��]�v���O~rѩS�৭]�v�7� �-��p.V)�Z�.y�&�g�	�03w�]�v8 �u��{K�.����8�| ����������@���SO=�����?288x�<p�\���ܹs100w�yg  ��6m��\�k��	�w�]����Rr0 �1�	cccY�N",_�<6o� �D[[ۙ (���?�g�/���`�r뭷�ضm[���D LWoo��  GR�\���<�C>ܙw�xKKK�={6 ��۷o߬>��jEgg���imm= sh``��{���'6m��Ю]����O~r�3�f���'}��   �l��幆K��!�T����@e;v,N�>=�>ܩ����ظ? f����~pp�C۶m�l�������C���K7+=z4/^  Զ���֭[�����<H�xkkkd��fF�NUH����H  ��gϞx�[�:���S+�,YW_}��M L�C0M�<����844t�O<�[���� (�9����}��  Զ��A�
��v�cȋ���ek���fF�NU�ڲ! �u{��q�ny;jI��v��  ���~s \�~��k��>�s��O��_|��G[GGG��zzz�  9�V�.��[�$����fF�NUh�@E�	�3e�;����S��b��r ��U�V5�^���6m����;w~�S��Ԓ'N�|K�;  �O�W&p'O,XY���gm�<T�;UA� �u����P���qڟk:#�$�鄂e"N�8� %O?���7l��������򕯼e˖-�Pe�����Sq�-�  �kӦM\���x@^d�34�fN�NU�ڝU �uq����馛���i@�|bԂ��ָ���'��<kkk�����?�K����ox�>�s��O���{�f���,���� ԰�G�N^�.�y�$k���fN�NUH�cӖ&� ��w���I�g777Ԃ+V܁�koo?@n����}����7m��Ю]���O}j�ɓ' kzzz��  j���05w�D��!p�j��O�� ���������Ԍ�������@�����f���SO=�����?288x�<p�� �֬Y3r44�� P�6o�����ȃ���̝���e망����.p�
J�{:�QW7��Ū+Ԓ�o�9���btt4 򪹹�` 5����~S__�#7n������϶m��011 ��̙3�aÆ���� ��c�;\����I��F�3'p�jdq Yv���x���k����	�P+���'#��۷@^555�i�����~����iӦ�v�����zh��ӧ�����
� jP��=\���<Y�`Ad��fN�N��@�)�3	�M���tvv:Q�ZCCÖ 2������_�����gv����~���:t( 򦧧'���/  ��t�kEa��;y"p�|�S5� Py)p�;�1���SkR��s�P��y晷|qhh���z�-[�n�/��g6l�S�Ne�"7  ��iӦ �L�N�d�/���	ܩN>@��}&�Ԛk��v��h�" �����k�:?�������Ν;?Q���裏�x/�O����U-��{�  j���F�N�,0�rE�N�hii���FKL@���kq�̙hkk���j�5uuu�S� oJ���g�yfG �nժUk׮�Ȏ;>�s�λz�%###������ j��͛��t�/�A}}�d_�5w�9�;U%�eu���  *�X,ƾ}�bŊ������Ԛ���;�K�����7O?���7l��������򕯼e˖-����� ��q�С8r�H �7111�A���O-��;̜���"p��ۻw����]:Y�`�Z�&���"���<ikk;@Ŭ_��������v��w|������o�����޽{���ҥK ��۴iS W���B^��0���y`f�T���  ��������Zq�UWŒ%K�����'���� ʦ����P(����+m����,=��QC+W� fo͚5��� @�m޼9�+��'�Zn3'p��������?�i��ϟ�Ss�w�;�7MMM��3����������M�����o�o�ᆸ��'�0s===w ��q�� �L�N�d�+���	ܩ*� Pq��ǁ��o���	�PkR����<���������u
��ף�_*m?7��OS�� ��&���~  ���ӧcpp0�+��'Y��^WW�<̂���"p���w��i�i�;Ԛe˖ECC��@��~�`Z^y�ť�*=�����b��1��K�{www 0sǏ�͛7�/��/  ٵ~����+s=��H�x[[[d��fG�NUI1Qss�` *,�w�y�>gtt4��455ś���صkW �Źs��pY�V�jX�p�m�Oh�p��=����w�bq֯�ދ��`�Ҋ\w �lK�;05���y���i�YS__��	ܩ:i9�; T֞={&Ü�
ܩU���w 7������ַ6�3���:
�B��Q��Kۢr}����x����������?��   ��05iP�\^�,H=a���#p��;�FFF ��ӧOǑ#Gbɒ%S��;����#~��@����a�[�v�����-=�*���o���_�r��`�^~��8s�L&�-  ��ɓ��Y	�<I=a���#p��du� Y744$p���K�N�)� �u��w'rj��խ---w��v���Q,�m��]w���?�� `����bݺuq��w  ٳaÆ����������w�'�;UG� �c����w�k�����Ԧ���X�lYlܸ1 j]kk례����(
]��c�b1E�-Q%~�q�ةS������� dT
܁�1��<�j�n�;̎���#p���&���S��8�4���C�tvv
܁\hll�ak֬���}���Ӯb��@������Qm�Ŏw����w�w�����  �400���ɋt޴��5�HK�#p�괷�O�r�� TV��~������9Y=���Y�bE �ASSӶ�200�>>>���Ӯ׷w�źȈ�+W
�fiǎ122K�,	  ���ɓ��S#p'/Ұܴw	�av�T�􋽭��r� 0҉C�;D\}�ձx��8z�h Բ��:�>�i�����������'�������"��� `v�*===��  ٱ~�z�a��q���x@\u�U�Ui�<0sw�R�1	��򆆆��;��ǟ;w.�VuvvF Բ.�dL___G�P�z#j/m��F�r�-�t��ػwo 0sw ��I�;05���'i�{V���#p�*��}��� T�����t��h	ܩew��544Ķm�\9����J�;?Xz��@�X���Gˣ���=��~�������NN4���  y��+�05w��w�/�;Ui� T���h8p n���)}���Z���1C�(�]u�U��We[�ΪU�.\x��ϟ?O�yc^��+W���ґ#Gbǎ�bŊ  ���<yrr05w�$ˁ�	�0;w�R�����r�~����Z���2���w�� �Emmm'�D___G�P�z=j��Җ��i�{��VV`�^|�E�; @F��펃a���EZ����5�(R���ܩJY��
 �n�������wJk�;�.�w�V577�'�NLL�Sz�U,�E��`ҢE���[o��7 3���?�p  P�֯_�ԍ�[��|�rCX__��ܩJo�}u���  *+ż��T�FGG''j��Z���?�я�����	��իW�����.=MڻJ�7�Yz�.j�ʕw�YZ�v���s��� @u۰aC Sg�;y�pav��P��	ܩZ�,�; T����d�~��7O�����.W��7�9���&o� �5�ʤX,֮]{G]]�d�^��yik	�䮻�����s 0s�|�+��w�yg  P��?CCCLM>�6ȃ,�&���	ܩZiu�С  *o���w���xX�lYlݺ5 jMSS��X̩�k��RWWw_��}�֭�P���`Fn��v�́���; @�[�~}�Q>��1��<Ir�J��'p�j-X�  �����:w�\@-����5itt���Yho�dB{�����hll�;�#V�^ �\
�{�  �z���:�;y"p�|�S������ۻwo���M�5W"p�֥��֤����ڀi���/�o��������?Pzl
�b�ʕw�YڲeK=z4/^  T�,2�!p'/��ۣ�!�y��f/���yw �?����eˮ��wjݛ���X�hQ?~< jłƞ|��р+����(
]�G�������H�; ���o��e��8  �>G��֪����z;(p���S�������)-� @��S	�ϟ?P�/_/��r Ԋ���S���{MSSӇJO���b���"�"�dɒ	 f���G� P�֭[�b1����.�,���	ܩjiG�" ̏]�v�>��+~�	��AGG���)---���jժ�������������B0�J�M⮻���?�G 0s/��b  P�^z� �g||< Lp�T������8x���t������VҒ߅��ڕ&����$�V����r������ޭ�����K[�G�԰�+W
�f)��H7�Oe�:  *'][z�W����VE^d}��~fO�NU���X �e���={&��+I!|kkk@�Z�`A\w�uq��� �ۃ�������Ӯb����㛃LH���� f���W� Pe�o�Ǐ`�.\�����9]�a��T��߉ Y�&�	��'�ς��MMM��500�>>>������&&&�+={�I�\s��{�t������O�� @�X�n] �#p'/���g���07�T5�`~N��Ν;P�:::�����ŗ��Q��YX�v�uuu]���9M���E ~"Mq��N__�d�&� P^z��)�.�;y�hѢ�2��an8�GUkii����ɩ� @�9r$�;W_}�e?N�N���S��!�u)x޷o_�i���7
��JOX�n݇J�]�	jR
ܟ{� `�Μ96l��o�=  ���ٖ-[�רȋ������S��K� �'Mq��;.�1w� ��7�|s�ܹ3 ��t�}�g�9dʫ�������+KO�^����;���hjj���� `�zzz�  U��_���� �G�N^,\�0�L�sC�N�KK���� 0?R�+p����������v:�z�V�jX�p�{���R�~�����SztV<��
���v[��� 3���|�+ ��[�vm �S,�B.�Uh�@"p��e}� Ⱥ���ɓ%�;;{�l@���o��o ���ڎU�����P(t�����JV�\)p��6ĉ'2� ��	�����N^���g>��Ü�S��l��566{��[n���N������Kj���_?yR��iÏ��jll�T����%���,=�*��\z�%�"R������ fnbb"^z���?  ̟�{�Ɓ��;y�hѢ�:�;�U�vZ �u����ܓ3gθ1�����[�|���?��jii�̋U�V5\u�U+���LS��(���+x�[��/��G� 3���+p �gk׮`�Ҋې���anܩzilkkk�={6 ���s�θ��{/�1i_�P�Ntvv
܁L+
������(�;磌�KS��/=^0M���;�o��o��{�� ��%p��1�����a��wf�O��v\w �?��'N\6`��&/R��e��ͮ"����믻p��JOS������7�.�3�r�J�;�,�޽{c�ҥ @�@� ��;y��w�uw2!�8 ����n��/p'/�͗K�,���� ȚX����s�����P(����+m���,=*ٙs)p`�z{{���D  Py7nt=	fH�N���EcccdY�����!p'j��, Ⱥ+�gΜ	ȋ���;�I����O>��`ƺ���;;;o�����K��K[s@�]��q�-����P 0sw ����K/0}�Ժ4h,�Lo��#p'���  �׮]�&O�
���}��Q,ݍL.�X�"֬Y Y�������(��z=j����s�஻���R
�/w~ ��Y�n] �gz;yQCp�0w�dB�y�X.Es ��8�|�����w�Ov�����ݭ�[��[�	r��Kb��qb'،cOg�;��U��o3��LU֙Tř�cc���n�!�Z@H��:�����b��H����ǣ�KX�����s���9.|�?�ާ����- �/^\�!�e Y����v�^|�Ů�kJ���/���:��J�t�@ P��Ǐ�K/��\sM  0q�;V>-�tw�"�S�Hr�V��Ȅuvv�ɓ' �<����IZq�S����`��x�� KοO~�~���+���_,��544���?6ԙ[n��|��MM��� &XZo7j�q-�����2�;�������ڽ{w�q���S�>}��"�����@洴���֯_ycc�]�����W��aȽ4 q��Ɩ-[���7���  `�lܸ1���)�4��FƲN��#p'3R�~���  &ϛo��N�*�5�����E�t��xꩧ K��۷GAmڴivCCç���]ccc�;�㢀����Ti�֭�k ���C�k�.���jG�Nf�� �\���={��W#��ٳg�b�������� Ȋ����T�k֬i���}dd䳿Xi����2W*��������������D  0��m�'O��2�)���S�Hr�V����; ԇݻw`�n��"ill�%K�Ď; +����G��_����?�u����Y�mkhд�/�]w]�f������� &Ⱥu��LZoO#d�wӦM�<���#p'3��ۣ��%Ν; ��I���ץ%��s�GW\q��Ȍ������_���ȑu���mnn����566����~��,}�^�|y�Z�* ����`  01�P9��E�o����jG�N��u�#G� 0yΞ=��y���?s�Ltvv��_ Y���u&2n�֭�###���û~�u��ؘ�v
���_�P�W_}5>��� ��ٷo_���TF�N������N��%p'SғZw �|�&��"f͚U>.�w�	�z���~,2�?�A�W\qCCCC9h����-W*���%�/|� ������SyXoO�P[w2%�C ��K����������E�V�7m� �����Pd����/oll��B�~�kz �bѢE1��8p�@ P���A�; �8K����	�)��4�S��q����Ȕ�<� Y���N�����fZp�"��+�@&����:��/�8w��g���]ccc�=�� >R<��@�Rlu��G444  ���%�ܹ3��	�)������)S�N���� `r���˗����)���"E ��������V��������CCC�<�cs �D�P��G��+��W^ye  P{�ׯ�w@ҽ�������K�n�j�+�LIq{WWW?~< �ɵk�.�;����}}}q��� �g---['��~����O�/���;��@UR�n�zw �q�nݺ *'n�:::�����;ԖW�3m�4�; ԁ�_=Ξ=mmm���阼s����P�i�]�Ի�����ڴi�솆�O��û���>�ǅ�Twww|�c��۷ �K�����  �5<<[�l	�r�+�]j�B���E���H Ⱥ��ꫯ�5�\�����w
%��>�l ԫ��������۾���Y������w���]���ill�!�qu�m�	���q������  �v�n���_����"�S���@��ɜ�; ԍ]�v�o�~�ԩ\=ieѢE�:�� �����l���[�l�ftt���y����_mL�������� �r���_�z� @�P�;E������A�5&p's� P?���S����Gm���$]�H��+�� �����j��6m�,~����gFGGg0�>��GGGG�% *700 p �����X�~} ���w)
���<��f��W���1���e u ���۷/���_�y�;E�^w�^�������֭[;GFFn��G��ky u���9n���X�zu P������� ��ؽ{w9r$���ɻ���܄�S�Ps^UdR:�D� �a׮]���ɴΑ�������@=iii��Q����M�/����w9h�#�O�k�RI�P��_~9�~��1cF  P���� �3::Z��<K`^ܡ���Ȥ����o 0��b�����b�ٳg˧�@Q̙3'�����ɓPoZZZ^~��_�~�卍�w]���M SR�@u�u����~�� ��	ܡz��)����ȋ��� jK�N&���- ȺS�N���c������i�]�N���<Ҋ�֭[�޴���s�������x������qq ��>�����Ç��� j��ѣ�{�� �#p��O���w�=�*2I� �e׮]����3g��_.p�J���p����'>�M�6���Ʊ��� r�[n��z( �\
� �^�\�N��322�g���1u����;ԞW����V�:{�l  �/��ԧ~��҂;MZPMK�.��)-��n��IK�.M��駿@n�J%�;@��I{��ŋ  �[�n] ճ�Nޥ����ESSS �%p'�zzz� P'�~��򑓿�؞ܡh����ٳ��7������Y�.���e�X���=dPimT� P�S�N9�jD�Nޥ�=O,�C�yU�Y�M.-�  �!���r��D��S�p1�j��O��ͱp��rО~����+��@q��������ʥ������ �ʬ]�V�5�D��)pO����@�	�ɬi9{� �.�4�R�W~�������P$)8MQ@����)bO1{�=fѢE�@�ߐ>����aÆrD� @eV�^@�FFF��G�M�>=��u^Yd�� ��o�Q>z����K�Y�NѤ���E�@5҅�A��%K���# >L
������@�҃�/��B�x� ��I���l�@��c"�����_y!p���Ef������144 ��K+;w�����)p��iii��޽{�b]��#�)l�7o^ \��n�ɵ2�H'r	� .]�5<<@���]����;��,2-��>|8 ���ꫯ
���
܁���s��}o�=���~�R)n���?�֭ *�¬o�� ��Y�zu �!p'�R�'w^Yd�� �K
z�bd�k��'OQ
V�x� �ei��Bоt����/j�T*	����/���ǣ��;  �8�O��M�6Pw�.o�{sss �'p'�zzz �###�gϞ���>V����˹s碥�%�H�ϟ��@quvv���/��[
�����@�FGGc�ƍq�w  g���1<<@m�{��W��_b�ƇW�����  v���^����W�NѤ3)jݾ}{ ő.`.Z����������� 媫�*�q�ر �rw �K��s�Pccc�ɵtbZSSS�E�$p���E��5�̥eX �>��꫿��~��)�QH)p�C�͞=;�-[V~ͧ��EL`2566ƭ���>�h P��k�  ��ٳ�iӦ j�z;y�:�$O�>�w]ɼ̽�� ԇ�(��+���W_]��)p�"Z�ti �����]vY9hOK�S�N�zR*�� Uڿ8p �ϟ  |�������P �a�����8^sss �C�N楧�� P_v���^�~���"Jg�g�cǎ�]�D�����/�<�͛ �,� Topp0���0  �p�=�\ �#p'���;�ƏW���cK  v��]^�hmm-/����ECCC@Ѥ��^dGz����+��)jOk펗����7/^{�� *700 p ��^�ƍ��;y��������;��.2O� �gdd$^y啸�kbtt��➷oT�b�8V��/}_y!hO_mmm�e���w�*�[��|M���1  x6l��g�P;w�,����ƏW�����8s�L  �㥗^*��ɓ'�Ғ%K�k���~ttt�_�����	P*�����~ P��Ǐ������k�  ��s�=@m	��3�;p)��ȅ3fā �{��)�v���N�8���E�~�ϛ7�gU�dius���lٲ�R{___��������7V������ ��܁�I�H�/ȫ����ƏW����DC P_�ŗ�;w���__^p��Z�t�Ϫ0	�
H���B{z���@Q�ӓR��e˖ �r��o~3  �M)n?s�L �c��<kjj����ȓ4������!p'��t ���;����Ƭ�RH)�}��_]]]q�e��_sW^ye�.�\�R�$p����?�O�����  �W�^�:��	ȫ4`���<����+�\Ho�)�K� P?����N�*/H���G(���������������+�i����σT �$��� Tnxx86n���~{  ����I�֭��,��g��ݼ����
#қ�ԩS���� ԏ���صkW�p�q��	�;���Ҫ�Ν;�\��SĞb��/Z�ȅC�q�זO�p��:���w �_�y���P[w�L�\*�0r#���a �gǎ����ɓE�b\�;\�t��Bоdɒ��� .Nz�n���jժ �r ���&��;y���=�6��;�1cƌx�� �/��9��i��*Ź�Gkii�Ĳe��_y��	0�J��� �J�w�ÇGooo  ���u��P{w�j�ԩ���-����
#7҂; P������������$��ٳ���'�}�� ����0w���V�/^�}��R�@��_�b  �v��
��FFF��U!��:h�l�ƕ���H�P
!R8 ԗ;v�M7�T^����
(��n޼9���E�A�ҥK���5 .����ǁ��	� ����z*�ڳ�N�͘1#򦡡��;�3�0r#��)r?v�X  �e���q���8q�����ST����e��_y���� L����x���ʥ�=-)���  E�z��[�P{w�,����a�	�ɕ���� �O�	�V��R/U�{S�xI�.�U,Z���k>=����'�D�RI�P���~;v��W]uU  �3�<�������H@��|;::"o�����*#WR��ꫯ PR���O~2��Ҋuooo:t( OR��"����=��.�ԏ[o��|� �:w ��V�Z����N^�q�=����gr%� @}:x�`��n(6PD)���]]]q�e���e˖E{{{ P�����~���_ *788���7 ��������J �C�N^͜93����?�2r%g��5
 ������Ν;�;�(G6PDi�z���Y���,(?��~ϛ7/ ȎR�$p��ƍ���= �"���'�G��Wy����O�N��:, PRTs��I�;��x�����.RR��������=��u�@v������ʝ;w.�l���� PD�>�l �cdd$ �R>u���#�;�?�;�����@}:|�p�ڵ��/����E���ݻ��������W[[[ ��_}���ӧO �� ���K/�0`F"�RǗF��&�35550���N^�5��X�fM|�(�ܩ)t\�d�{A��i��|JkB7�tS<��s@� ���z� Ə����k�g�&����IQFccc��� P�n�Z�H�����RH�r�ʀ�v���k0-�����r5��W*�� Uz�����C; @������ի?w�j�������I����ıc� �?'O���k����PDs�΍���8u�T�x�>}z9f_�lY9l�p@q���ꌍ�źu��s��\  ŦM��w�	`��ɣtO*5|y�~L�4r)=�%p���j�*�;����,Y۶m���������1��W^��� Iz੷�7> Tn``@� J���/�;y�F��z��w�wr)�j  �i���q������(�ܩ����X�`A��T
���r{����z뭱bŊ �r)p (��gϖO��O:)jtt4 ofΜye�&�W��w �~��ի㳟�l@�*������=�:Jk�MMM ���_�P�7�|3���S>�  �֬YS�܁�c����s�g�&���\Jk�mmm���:����)�����5kV9r$ࣤ#/������ �J��==,��� �\Zq� E��SO0���QgJ�C󨱱��L�;���;x�`  �i���q�С�;wn@�PY���I�/�)p�ZH�_y啱s�� �r)p��׾  y��;��֭[_w�(��J!xYo��#p'�� P��j��O?_��W�h�ҥ�nݺ�t�/=�s!j_�xqn/�0�J����J6l���a7��\K�pFFF_w�(u{y�������[y~���x��'�օ�ytt4(��\q!hO;��� L�������� �rgΜ�m۶ō7�  y��c�0���Q��=�����[�:@�:p�@���˱lٲ��IA���^򯳳��PÅ����' `2,_���9dhh( ������ ȭt�׾}�w�&�z���+�;L�;�u����ѣ ԯ��.p��҂��=��ŭ������羾�hhh �l��n�!�ʭ]�6���o @�\�2��722cccyra�6��0q���̙3� P�y��ַ��A
)-y?��SA��x=E�)fOQ��E�b��rP�J����J۷o�w�}��L @�;w�|���ɣY�fE^��������j'c�  ��IDAT#�R� Է'N��������f������CCCA���A��%K���#  ����ꌎ��ƍ�ӟ�t  ���ի�ԩS�?�;y��^�hL,�;���0ӓS�����j�*�;����Ka�;�����,(�)l�7o^ @-[�,f̘o��v P����; �;+W�`b����IZ7�6mZ��&���\Ko*S�N��Ǐ P�֭[W~����(�K��SzX���ｕ�ŋ�J ��K�q��zk<��#@�֬Y  yr�Сضm[ Â;y�N?N��J�K�N�w�; Է�N��3���w�P4)��~�o���K�Fkkk @�J%�;@�<���� @<���1::����7�f͊<K�=G�N��}Ϟ= Է'�|R�N!�=)�>v�X0�:;;�������� �"H�; ��/�� �u)l�'�8i�$uzyf�&������' ��Ν;���_��MZ߸qc0��L��-*���{___��J�2gΜ�C^{�� *'p �b˖-��[o01�z���X@^�����;�*�OL����G�utt��N�> @}{�����f@Ѥ�Z�>~fϞ˖-+�{Nq��O �si�]�P�u�֕�N  ��=`���$���yT*�_l0��]}
!��
���=����o|��^NZOD,u�FWWW\v�e�������S� �R����}/ �܉'b���q�� @V��4���L�;y���<�0���S����_ �����h��o�=�H��ۣ��/<\����X�`A9hO̛7/ ���|����� �I�2� @��Z�*����8�ǐ7w���B��@ Oy��;���l���Ik�遀��oi����) �K����]w]l޼9 �\
ܿ��o @V�v��522�i�*�'*�a�	�)������s� �o�?�|9��LѤP��g���������W[[[  �+�Jw�*�k�N�*?8 �5���J�޽;��e��<�5kV�]j��%p�0f̘�
 ������ʕ+��{�(�E�y(�tttĒ%K�ڧM� @���o��o�ʥ0eӦMN� 2)ݓ&V�j��<�9sf�Y:]ڂ;L<�;���H� ��(̯�����P��{���ZN566�ܹscٲeq�UWE___�b 0�������w�}7 ������ Ȝ���x���X��ɛ�/�O�2�}K�w
c��� dñc�bpp0~��;�H�Ry���ӧ��_^��^�ti��� 0��Cf˗/�'�|2 �\
� �f͚5q��� &���<ioo/�̜g�n`�	�)��D����! ���G�S8)�γ���������gt `�J%�;@���������  Ȋ�+W0�K�IFg����xw
#�Q͜9�|� ��7ovc�3gN9��bN�سp��rО������ u(� T/�F��/~1  ��СC����0���Iw�09�ʬY�� �����启��E����g��B��?E��!E�-*�� Է�������@�� @f<����{1������`��;�09�J
���H��׾��hjj
(��g)p�>}�{A��%K���# ��I+�?�я�ʥ�=Eb�DY �z6<<O<�D �cdd$ zzzr���Y��B�N�L�6�� �IH Ȇ�G��ƍ��[o(��K��/����E=JG��e˖��R� d���z��N�ڵ��� @={��g˟]����uzyQ��Yq;L�;��VSұ(�  y��;�����gώ7�|3�A�=w���V�/^l� r(}�N��n�T'����z����,��a��<I�4�.��C�N�� [6l�o��V!�9�RL>��{Ze���E����  �m�ԩq��WǶm���ƽ��  �jϞ=�cǎ &����hjj�iӦE�Yp��#p�p�q �-iA�'��?��?(���տ����Y^fO�+��2��� (�R�$p�ҦM�bhhȃ� @����� &����H#�E8�ق;L�;����2e�� �!�<�H���Q!�A�$�����5��-ZT��R{___444 Pl)p�_�� �;w�\l޼��{* @�9}�t<���L�yQ��Y�;L�;��¸3fěo� @69r�|sx���E�.�,X� ���[��^��SĞb����=E�  ����/��r�ԩ �r���w �.=��q�̙ &�����5kV�]������
)��
� [}�Q�;��B�j�������⪫��e˖E{{{  |�� �M7��>�l P��������? @�I'��kdd$ ������"��z;L.�;�T�'�  o����o�]>�� ��?���߿��������7o^  \���~�;@�v��G���3g @�x�jvj(P���>66�u�gώ"hnn`��)�ƥE*�� @v�5��+W�W��Հ"�?~ttt��ӧ���744D___9fOQ{ZkwD P�R� T'+�֭���� P/�����)�E����K�N!�(E�o��f  �����W��/��>�.Y�$^|���~n������+� PK�Fooo>|8 �\:�N� ԋcǎ��ի�\i��.���A�Na�7Z�; dˑ#Gb`` ~�w~'�~�~+�ڻ�� `�����O�� �r�� @�H'�Z����uH���"�N!sss �G�Na͙3'�o� @��X�B�Na\w�u�/ ��$p�^�ٽ{w�d ��4::�>�h �O�N̞=;�`ʔ)�!2`��)�iӦ���  ;�m�{��%K�  P{��v[��M�  �\Zq� �m���q��� &���<H��EP��z�ww
+#��(;x�`  ���C����1  ��K�W^ye����@��O��O `2��g?`򍍍���H@��1ٞ��(�;L>�;�&p�lZ�jU�ٟ�YL�:5  ��+�Jw�*mذ!Ν;�8 0i:�7o`�Yo'Rk�Fe����0��Zz� �'�~����_�r   �������w�ʝ9s&�m�7�tS  L��~8FGG�|w�H���&���BK��mmmq���  �%���/})  ��c������P P����; 0)���c�ʕ��;yP�������L.�;�7gΜx�� ȖÇǺu�T*  P[i���o,�� T.�>���ݿ ���jժ8~�x �A�N�uww�1��z;��;���,�@6�X�B�  㤿�_�P��۷ǻ�=== 0��=�~���dY�-
�;��;�W�7_ ț�[�ƾ}���.  ���ä����� �r����aÆ��g>  e˖-�gϞ �w�.��������kkk����8y�d  �����ώ� �qp�UW�̙3��ѣ@��iw `"=���ԏ��k����2eJL�>=�B��A���'�� �MO<�D|��(?�  �NCCC�r�-��#� �[�vm  L���ƍ���ɺY�f��A��lnn`�	��9s�8� 2jhh���s�=  �V�T�T)Ef��� �xK�햢���ɺ����v�w��/������� Ȟ+V����hll  �vR�@��+_�J  ��S�NœO>@}��u��+
�;��;����6mZ;v, ��9t�Plڴ)n���   j'�3-Y��� U� !��u�̙ ���,����(
�;��;�B�Y'p��J+�w  ����.p�����cdd$��� `<��=�P �G�N����F�ܡ~��R����/ �Mi�}����`��   j'���w_ P�'N������ ��f͚x뭷�?�Ȫ��ECC����~a�̙������ d���X��g?�����  �v�II��ιs�����q��$������}LȢtM���'�"��)r��~!�9͚5+�x�  �����������  @m���ǵ�^[>5	�ʥ������ ��v����z�S��ɲ��^�໵�5��!p�_���+p�;}�t�\�2��   j�T*	������ǩS����3  j��?�q �)-�CV���H�b=P?��K�Sg @����w�}w455  P)p���� �ri�q�ƍq�w @�=z4֬Y@}��Ui�}֬YQ$ܡ��ᗤՔ��T �l:r�H<��3q�w  PW_}u���Ļ� Tn``@� ��O���t@}��U3gΌ)S��������9��Q�߁�"��Uv�� @v��G?�O}�S�oB ��566��7�O<�D P�� ����P<��c�/�;Y5gΜ(��������� ����[�n�n�!  ��(�Jw�*�k�.ߋ  ���?'N��>���9a��*Z����@}�ï�5kVy�jtt4 ��z���  PC��v[ P���~�=� @5R8�bŊ ��v����+:;;�HZZZ�/w�5S�L�3fđ#G ȮM�6�Oe����  �޼y�b����� �rw �6l���3�sw��h��w�?wx�hP�; d�O~��˿��   j�T*���� Tnpp�|�l:M �R�$[��	�ɪ��ܡ	��}����_  ۞~����?�Ә={v   ��T�wމ�;w��>��  �D�,��/P�FFF�fʔ)1cƌ(q;�'�;������#CCC dW�h�bŊ�����  P�[n���8����\Zq� ���@���N����h^$w�Ow� �����_  �~����W����  Tg�ԩq��WǶm���Ľ��  �j������'p'�z{{�h�.P��қ�� ��̙3��#�ė���   �w�m�	���y��8{�l��� ���������^�^�dM:�1���w�Ow� )pOǭ��� �m?��O�{�)S|� �j�J����� �;w�\9rO \�#G��SO=@���N͜9�p��S(p��T�ߍ��7�iӦűc� ȶ�G��3�<����  ����_���q�ԩ �r���w �����?�BFx��Ei�hZ[[�Ow��M[� ���ĝw�Y~  �\SSS�t�M��� � ��u�ĉx����;YT���z;�/�;|��s�Ǝ; Ⱦ�{�ƦM�b���  T�T*	���k׮8r�H̚5+  >ʊ+�̙3d������鉶��(�"�3CV��CL�>��&v���  �/��� �z)p�:ccc�nݺ�����  �0CCC��C�w�&��w�_w���}�� �}[�n�W_}5���   *�dɒ�u�Ç �� �G��Ǐ�###Y���MSSSL�"��z��	A� ����8���/  T���?~�ӟ �(/�744 ��I��>@v��m��Y���S�N��imm�~	��#̙3�|a�O ȇg�}6��o��� �ʕJ%�;@��z�ؽ{��� ��jժx��7Ȏ��	Ȓ�s�F	ܡ�	��#477ǬY�����K�	?�я����v   �K�{ccc��� �� �+�i�l��5���QDw�ow��)5�; ��c�=�G3g�  �2ӦM����*v�� Tn`` ��O�$  ~]���o߾ �E�N����3fD�444DKKK �K�!�/��B  �0<<\^<�ַ�  @����� Uڸqc�;w΍u �7�i����%i�=��E���t:%P��p������3N�: @><����|��:	  T�T*�w�� �rgΜ)��,_�<  .x���=P%p'KR�^D����7�;\����ꫯ �CCC���ƽ��  @en����͠������_q����=ccc122�MMM1{��("��A���E�@�<��C�/})���  �t�F�M7�k׮ *�����}  ${��͛7�=��ɒ��Ƚ�����ow�H�f͊)S�� 
 9�� _�bE���o  �L���J/��R������  �����+�@�Xo'K��������9��&p������̙  ?|���W��_Eggg   ��T* ������]w� @��۷�CĐa�3Ɋ����{���P��p	z{{� �3�O���z(��կ  p鮼�ʘ9sf=z4 ������ �����Mw�"��E]1oii	��	���cY6o� @���'?�/~����  ��IkO��zk<���@�R� �k��k֬	 ��d�ܹs��,�C6���7�iӦ�;� @~�8q"y��җ�  ������T)� ���� (��~����!��dA���퍢�C6������ �?<�@������  ���v[�����X P���.p�b��ٗP�
Y0cƌ��onn���� ��.Q___�ر# �|9v�X<��cq��w  pifϞK�,�ݻw �K������: �������q��ɊԿ��v��;\�iӦE{{{�9s& �|�����s��\L��c2  \�R�$p�҆bddĚ �믿�W� ��dA:����7����-�lP�@�Sln�@�9r$��r�  \������w� T�ĉ��/���_ @qXo�|��iܵȑ�w��;T@� ��V�?���ZJ �Kt��7GKKK�;w. ������ 
$��?��sd_:�	��ܹs��R���@6ܡ�g�.�� �/����z*>��  p�����뮋�7 �K��_��_ P������CNXp'��[o�l�CbΜ9q���  ��{��^�y����  ��+�Jw�*���q�ԩ���  �<�<�L � p�����DGGG���E�����@N�����@��   .^��_�U P����ذaC|�  ���>���s���X@=+�z{"p�l�C��~Zr�� �)	��O|;  \��������� ��@��߿?�~�� ��z;Y�]�*u~w��;T���9f͚o��V  ��o߾x��g�L �K���[��� *788 @�����w�]���쌢jii)G�@vܡ
�6�; ������������  ��)�Jw�*�ݻ7<���  �x�x�g��;�����I[[[ �"p�*�7��> �|J7��x������   .N
�������{�	  ��	 ?�Ի�s�F�����-w�BGGGtww���� ȧt���;����   >ZZ^�`A�߿? ������ r(��?������z������Qdw��;T)��� ��z�x��G���  ���v�m���0 �\
�GGG���1 �����366�uM]K}[��1���� �E�UJ ^~��  �����~|����T7  \�R�$p�һ�;w}�c �Á��C�۩wE���l�C��O����q�̙  ��رc��Cŗ���   >��7�\^Er��:i�]� ��O��O�O������z5mڴ���"kkk {�Ps�΍={� �_?�я���|�� ��1u�Ը���^ *��?��?  �v��k֬	 �Գ���'w�&�;���y�� �sǏ�|0����  ��n��6�;@�6o�\>A6�$ d�w�� �Գ����)Sd��E^�P�gώ���8w�\  ����8����%  ��J�R����} P����زeK��!  ��m�V~O�I�N��6mZ�����%p�hhh��s��k�� @~�>}:x�����{  �p�]w]tvvƩS���� ����1���S���ޞ�!��P#����@�X�"���/����  �`����˗�3�< T.� @v�]�6v��@>������	��ew����ޘ2e��2 �Ξ=������y   �T*	����+�đ#Gb֬Y dK�^����?�N�z����ۣ�� Gsss �$p�ill,G�  �~���ŗ��%7� �#���ꌍ�źu����� ȖU�Vž}��/�;�j޼yQt��!��PC郁� �oxx8�������!  ��x��;wn:t( ������ 2&E���w_ �622Po���/�N��&p�J7���&>�@��\�2�򕯔�� ����>�` P��kז��S�  dC:�þ�ܩG�$����(:�;d��jhʔ)1gΜx�7 ȷ�@�w����˿��   >X�T�T��ѣ�{���+ �gϞ�������z4o޼(����hnn ��Pc��� �ᩧ��?��?�ŋ  ��҂{��4���w��u�wb�?�,Y�WI������- %��$�d�i'i;���i���s2�i����t�93g��¾�`a	K 4,���I�%[ 0а�l˶,����CE������{��z��[�Bb�����y?ߑ� �r}}}w ���w�ƍ�?�;�&��م��v�w8��!�ͭB�����7����o��  ��gώ�?>~�_ ����_�� @u۲eK�~��Կ��YD��;wnL�"�C��L�YKKKtwwǺu� �<�@<��Sq�	'  ����w�1z��c�Ν�} �z�v�m144@�3��j4��@��@�� O� P9�aٲeq����   o�����^ Tn�����c��{���  �ӆ�{�	��T��ܞ�Yˮ����p�w��͋G}�6D P9������v  ��:�S��IgP��� p��u�M7Ŏ;(�;�&�����(��S�P��0�f]ggg�_�> �r�i�g�q�  �91��SO��˗ �������C  �g͚5��}/���Sm�ϟ����O��$O� P�V���~�����?  �r�#�;���.r1{��  ��7�������<�$Ltuummm�>�;�����  ����f|������   �,w �fdd$V�X��� ��<�L��'?	�<���c�;U%[����(����"�j���I�m�q��  �!_�o������?  ��{�1gΜx����������\}��E�
����T�܉hmm�>�a-\�P� %��o;~���w  �_�	Rg�yf�{�@�/_ @���OO>�d �bz;�dt+mmm��;����? @y�ܹ3n�����>  ���������_�_|1-Z ��������|�T���w�wG�"l���100 @y|��ߏ���߉c�9&  �_y���_Lr߳gO P���>�; T���;֬Y@�ܩ&."������9�� p�qv�QG	��dFFF���F����M   ����U,}������������ 0y�l���rK ����R���}xx�b~&M_�6mZ`z;��;���O<�D J桇����gqꩧ  �+===w�1z����f��� `��|��E��S{{{q���}4v��صkW�1��l�x��ꋫ^0����b�̙�iӦ  ��k���.�(  x]ooo�t�M@�n�?�����O `���+q���������W���}4v�;~7,��jhh�y����N�w� y"!p����/?�я���  ��N?��b�;w ������$Y�lY����s���422�F��o /~�`tww�ԩS�8���]�0�,YO?���O (�뮻.>����   �ONRz�{�=�P P������?��  &�/~�b��X�.�y477�i�t�E��=�}4~�a��׵��P_�0�$t���e˖  �e���q��w�����  𺞞�;�=���188X�  &FF�W]u��v��ʩ�MMMű������=������i�GqD�� �A�d�ܹw (�[o�5>����̙3  �����.�, �\�,�X���p  �G?�Q<��30Y���������;���3o޼b�3���&Ȃ�瞳Z Jh�֭q�-��g>�   "N8ᄘ={v �������H����j��{KKKq�-[���G'��NϏ��Ԧl�x].��C����5kV�M�)� PN��sO|򓟌#�<2  ����g���������� 01���X�n] Ԛ���"��_ �����!�ի��-:;;���P�0A�$1O,� PNy!hٲe���  D������^�5k����� ?�6m��n�- �́���������w������p�׵��P�0��Ν/���� PR˗/��+W�i��  Pv�{����{����� ����bhh( ��@S߳{��G#�<�cM������e�/p��$p�	4s�̘6mZ PN_�����K/���   (�y���QG/��R P���>�; ��U�V�}�� �.��)S�ǾFFF�������1k֬�>}z��} w" ��&P�����@�e�s�=�ħ>��  ���)�w�����/"7�`|,[��4xg��$��<�6:�}��}���3������@}��jnn���.7� ��n���Ї>T�� �2���[o�5 �ܦM��駟�N8! ���g?�Y�X�" �w��~��=�x~%̟??��8�'�;L��"f�̙�y��  �)ws����㳟�l  @��y�ōM�T�M__�� �|��կ~5 _m瑃C�5����ڵ��;kq�o��_f�}#p��%p�	�/�w (���/>���q�  PVӦM�w�����c� ������� ��s�wƪU������T����9�=c�}������QG�����&X��Ξ=;^z饺>� �^�\u�U��/�ؒ  ʪ��W�0F�<�Hl۶-��� ��7ƭ�� T���z��=�ÎN|��>�g_��N������x�M�,���c֬Yśb ���z��?���ć>��  ����=P��6~��������  �nٲe144 Ԟ�����>k� z4v�����W����;�7�;L������!p �k����ۧ PZ'�tRL�>=�����	��0x��'��?�q Pf����߫i���_�2eJq ��#&Al3g�,^d�D (�����m������  �(o*�~���1�� ���⊪��{O}�W�6�Nz�w��D�={v̘1#��ۡ�	�ad��[����k�� @��q����1��  �2������s�=W�s�3gN  ����{㗿�e ���[ZZ�co�*����}��=?8���Vw�w���/'Sutt���"�׿���˿��  �2���	 �&�����G�� p�l�7�xc �����屯�3v�{���q���d`oPڛ�}���&I���IK��� �|��X�re�v�i  e�dɒ�Fݚ5k�����	��B�]w]��Xe��Gva��G���=�}�<����=e6u�����ow�$�oݺ���nݺ  ����K.��*  �wg�yf�y�@�2p�i�9� 8x�=�\�w�} ��@S���h����w�����v(�;L��Z�; 0��_�{�'>��O  �Moo��`�֯__z�{l  '���/�<FFF &K.T�2eJq�-w<\�vm1�<{�<���q�s[[[ �O��$����x����	ǎ; ছn�}�C1k֬  �2���)�� �MNq�����~O?�t @�ʉ�CCCű���ZZZ�����c=�����x3�;L�<�غuk1���W^	 ��������㳟�l  @��"�_��_���z* �\���_��  �Y���]w] @�ʡ�ylٲ�M����{��|��*�ۡ<�0�F���N�; ����/~��;�.]  P&���w�1Z�re�ܹ�� ��w�7�ƍ �́��744�����?����w(�;L���<Ahoo��62 @�����e�]�w^M�� �C���׿�� �r۷o�G}4�8�  ��_���; �L�������}��g׶������w(�;L�)S���ݻ�)�w `�3�<���w�I�  P��rJq�j۶m@����� �����b�- ���͛7���2p�{�����'J�MMM���&Yް۲eK̞=;V�^]�(  ��\�,;::  � o��z��� �[�|y|��� `����x�� 88�v�*����6:�}t��������� �C��l4pϛw3f�x��7 ��rw�k��&���O  e��<� c���O�ƍ-����k�W_}u  c����}����Ƣ��{��葿v����C��,_�s%[��wvv
��7����G��O  (������x衇�c�X  ov�7�k�� �����[�n-�}555�����GC�l���A��T7�;L�|����;w�Y�f/��� 0��.+�<g  �z�t�Ҙ3g��`����� ���>���  &�������3z��}t�{WWW �"p�*�+�2pϸ=�]�~}  �Z�fM�~�����  �.'4�y�q�� ��� ��4w�%�A P�v��Q[�ly�s�>�l1nڴi�1cƌ�9s�?�!�@}�Cȕf�6m*~���)p ��[n�}�C1o޼  �z���+p��_~9^x�X�xq  QLn�� �M�v튁����[�hoo/B��ӧ�����@m�C��=_h���S���*�
(�|�o޼��^)wv H�f��+�����  ��}�{��� �\�� �7n�n�! �����n�Z���&{���s�{��9�=��T/�;T��Y�Q���ۋ�;::�W^	�|r{��-��B[F� �V�\?��O��`  @=���K�.-��r}}}����� e�d��� (����b�d�ʡ��y�{b��T�;T�|��;;;�P2��4�Pڶm���䞫FF]u�Uq�i��� ����������ݻwǔ)n	P^=�P<�� ���r�����YP%��ڊ�5�4�����m
P�ӆ��588Xl��� it�?��?  �g���q�7 ��I�O<�D�r�) e��ڕW^  ������@�C�Ȩ�����%uttܡ�Zƪ������/9a)Cw�t�=��G>�8���  ��駟---�s�� �r���w J+��= ؟E�P��PEZ[[�i*)�իWǞ={�O�xݹ����@Nxϕ�� �\~��q���{^  �n嵲�O>9V�X T����Np ��/����w `_9dr���T/�;T�����<s��شiS �%��|l�>����p�wuuECCC <���$�O~�  ����G�0FO<�D���� �"�\r�%�=6 �}-X� ����^w�"mmmo����S�uf4Tߵk�!��ܒ}���1k֬ H�_}����/�  @=���K/�4 �\^���B��G ���{�_�� �?�-
��	ܡ���'9�}��������1P�2Pϸ='FTj�֭�sE{{{ �NW_}u����_  �ѻ�����舍7 �����P��!�  �ϴi��� p�*�Sܷl�R�������ׯ_@m�5wdسgϘ���{r�KKKK ��'?����ߌ����  �����8����� T���/ �,��կC�  �g���T?�;T���4g��;԰�3H���p��9y������p�Wƥ�^���  ����W�0F/��b�^�:,X P�z衸��� `r��QG@��C��0-_HG�<����۾}{ �exx��w��9.���-��9(�W^y��n�3��L  @�����{����� P�v��Q� 8�6�=P��Per�ԩS��wvvƚ5k��g�>222���͛7ǬY�஻�|���w�;  ��̛7/-ZTL�r}}}w ��M7�T� 8�ŋP�P����������oLu��֭[��|"���jnn��(�\z�q�E�  POr���`lr�{^?�A; Po�{��; �@�L�R� j���P�7n|���fΜ�6m
�zeО�ӡ��	���3O�[ZZ(�~n������?  PO2p���[���u�_��v����_\� p ���/��6x�B�H����Mo�s����W>^sa�Ν;'���a������x� ��[��V���K�  ԋ3�8����{�� �r}}}w ��-��RLp x;�/�vܡJ�����7>�5kV1�}׮]T�|\f`>�S!rk�컺����!����/��8,z �^L�6-~��=}�� �r����o�� �/��R�v�m �v��ۋ��w�R���Ξ=;^}�� �Ƕm�b``���>�rz|����@��򗿌;�#��?��  ����W�0F�<�H7������.���8 �-Z���H�1w�R���ŋ���l�"�C�ؼy��T��9��=�d;��n�����)ި @=��ۯ~��@�2 ���~�� j]zy�g ���o�G�U�����Ts"����֭[�<###�aÆ7=>�I�������@y��K/�4�>��hll  �u'�tRL�>���Ԛ��>�; 5oժUŠ �w2g��"�	ܡ��������w�D�fܞ[V���!�7vww�e��z��'��{�����	  �u����}o��G?
 *��� P�r��_\ܷ x'�/��ܡ������s��^��x�L�m۶���@�W��)�
���!����k���#�  �u���w�1z��gc�ڵ1w�� �Zt�]w^  �Isss̟??��#p�*��{cc�b��x֬Y�q�� &��͛kn��Z�A~GGG �}��b��Yg�e�  5���' �+V������+��7�  c��1e�Lj�G.T����غu�>���%p�	�L��cǎ�E9u>W�N�>=��z���?�A|��  �e��pޔ��\__������,_z���/ ���dɒ j������U[ZZb�Ν�����aÆ�Z���3r�:uj �u�UWũ��Z,� �Zv�gƷ��� �r���E$h�7 jɽ���<�H  ��3gFGGG �I�U.�����G�ǝ����k����oz�ղ�B?g��.A��e�]��  P�z{{� c�~��x����c� ��֭�k��6  ���P�TnP嚚��i�;v�x��3p_�vm�ķPMr����`ԓ���7"wS���|�������7~�7  jUNpoll,��P��˗��	yO��K/-T ��~x�QGP��Pr�����ԩSc���e˖ ��8����ۣ�ڵ����d�����㤓N�Y�f  Ԣ<�}׻�O>�d P�������? P�����ʕ+ �`-X��*�.�;Ԁ���x��s���ݻwǆ��Y��9�>� 唻T|�k_�����s  @������Q��9\'� @�Z�~},[�,  ��ŋ�mw������)�������V5eʔ�ra�e���Hʲ�yƭ�����@9��G?������?  P��|��k�	 *�q�c�=g�qF @����+c�֭ p��M�V�j��jDNq�wZ{CCCtvvƺu��L>�ʸB�y2��;PN�_~y�x����  PkN9�hkk�m۶ �����P�~������ �P�����ڦj��7���f�*p�C�gϞظqc1���rZ������I=�T�W\p��?����<  @�inn�SO=5x�� �r����� �����㪫�
 �C���-Z@��C���=_�3���ԩSc���188��ٽ{ww�e���3�ϝ �rZ�re|��ߍO|�  ����W�0FO?�tq��o T��'~�%��rf `l�Ν[tv@��C�ȸ���u��.wuu	�� ������b�9��{���3fPNW_}u��=����  Ԓ���N�bŊ����� �jq��w�C=  �j�����;Ԑ\]���='��Z�*���8�\�y����2pϭ�sP>���.�s�9'  j�ҥKcΜ9��k� �����P5����^  �*��y��P�PC���cÆo�|Nw���W_}5���ms�݌8ٿ�����)S�@=��S��o;~��~/  �V�5������{��-_�< ��@���??v��  �jѢE�5C�>�ؠ�dx�S�w����_�iUwx�ݻwC�G,�S>����t�7�駟K�,	  ����w�1Z�vm<���	 0�n���x�g ���C�5���m��{n��އ��x]Nw���###�;�E �����@���Ź�^xa��  jA�9�)nP���~�; ���g��[o�5  *�g̘@��C�Ɉ}������|�~���<�c��E[�lq�%��/�7�����?��  �Z����.]Z�0 T���/���  `2�����;/��� ��/��ܡ�������N����իW{�O��Ķ���ضm[P�ܧL�R��Ϸ���8����O  �9�]�06+V�(vx�� 0Ѯ��X�jU  T���%.\@}q�
jPF�[�n}��3|�={v�_�>��rqǆb׮]���"������@��"�/�0.���b�  �v��p�@円��'��SN9% `"=��#q�� @�-ZTts@}�C��l�{����SJ;w�,����n���I����)�@����+q��ƿ���>  ���D9�)� P���>�; *�y����/ P���>:��#p�����F?-���e188�7o����q�����
�|����_�$̌�  �������'�+V� *�����w�. `�\~����k� @�rp�����?w�A9M9o�m۶m���1���2�E�6m��>�v��Q,�9sf �ϱ99��.�3f  T�\�)p�'�xµ@ &�<?�� `,Lo��%p�����wvvƚ5k���P�F���~|�������y(�6ĕW^����  �j���%�\ Tndd$~����G> 0��ڳ�w `�r@�����Ow�Q�������	������(�����.L�����2eJ��t2��?  P�~��~-:::��� T���_����=t˖- 0�/���� ��jT��---�^=g��;uihh(6m�T\�b��w.*���.� �r饗��G  P���g���w_ P��˗ ��{�7V�\  c�a��%K�_w�a9��@�{n�2c�+ߩXg؞�;�cxx��ܻ������ٺuk�w�yq��g[� @�ʝ�� c��K/��իc�� ��+���^{m  ��ܹs�v�_w�a�"=00p�_�U�N=Ȱ:�?Ђ&N~6o��f�
�\�|�ɸ���_��  P����� c������� p8�޽;���/Ƕm� `��>�� ��jXKKKL�2���?Ť�]�vԪ�3n�ȝꐓ������������N*  �69�i�����/ ��0��o�3�<  c���V\��j\�9M�@:;;c�ڵ�hhh(6m�{��	�K~]r�M.��cdd$���%�\3f�  �6���w�1��=�466 +W��;�3  ������@}�C��io�ϙ3'֭['�������`P��9%'��sLSSS ���k������=  ��d�~�-� ��k�O=�T����z �X�\P,� �\���8�O�5.�|�>����<s��b�2Ԃ�^�pzǎAu.�V]]]V�B�<���w�w�O|"  ������-v۽{w P���>�; c��.���~ ��p�GFkkk �O�u #��[���s²��Z�k׮ذaCNSv��YLt�5kV ��}���}�QG  T�iӦŉ'��<�H P������?�� ����;bŊ p�}������@{{���9�}�ԩ&bSնm�VlQ���-�����\<���sN���Ŏ1  P-zzz� c�裏��Аk~ T��g��믿>  �n���@9ܡ����������b͚5�('��+w��-�E�P.�?�|\{����  բ��7��կ ���6W�\��� p�r�չ��w� ���c�)9��P�����Pp ����˦cSUFFFb�ƍv��ܒ_�9s�DSSS �q�]wũ��g�qF  @58餓�sA= �����P��/�<V�^  �K�q�-
�<�P'r�з�s�rGGGlذ!����~�C~-3r�5V�By��.� .������  �ly����O����@���� �~��� �a�p��hii	�<�P'2p�X��&��de�;� c�Q��ܹ36m��g��<r2fn7{�Yg1  L���Q�=��s�v�ژ;wn ���ů���  8܎9� �E�u����X��cǎ��iӦE[[��Nz�����`P��������x������;�#��?�g  ����7 �|0>��O ��ݻw��g��^4 p�uttP.w�#��]�������_�h###�q��w��>�B���m�r���ǉ'��z׻  &ӢE�b���z�� �r���w �׿��b� ��m�ҥ����H{{{lذ�mO�f[�fM��&ʮ]����������S|�sQM�0�C>ϟw�yq���%  0�zzz�]� �\�y����! �@~����w�  ��ԩS�A@�ܡ�L�2����s���������ꊵk�L��۷���&�S�3r�3g�`P"���J���_�E  �d��������g���;. `�>��^�^  0.�>��w�G�ufڴio���M׭[�"�n���188�WN�(v� ���������я~4  `�d��7�r6 �[�|�����s�|�+E� p�嵽܁r�C�ioo�9�}֬YEt
�!O��aNo�m۶�;� (��.���ذt��  ��0s��8���?�y P������?�� �}�~����#� �x�7o^���PNw�3���EH�NSܻ��ݻwǆ�aԦM�bʔ)1u�� �!wp8��s����/� �d�������?;v�pm�7y��'�n ��r�1�P^w�C��S�>}��b��	�N���'l����T�\\���@9�Z�*.��������  �����˖- *��}��8��3 R�<�sbxx8  �C��8gΜ �K�u(���Ξ��K/�p8��͛$>�t�|���@9���q�]w�'?��  ��v��'�ʆ�������	�(���ܹs��� 0^�.]@�	ܡ���Dsss�ڵ�m_ggg�Y���z�dϞ=�dn�p0�y)�_��(����:�=��8�  &R^#;��S�?�i P��?��� �t�M�r��  /yMo�����TN�ڴi�������"2}��W*�{��b"w�+C����ӧP��.����⋋��  `"���
���駟.�\Pn�>�h�z� 0��,YS�H[��<@�:��=q���k�S��P�ر��ĝ�¡ڼys�f���5�r��ܶ������Ev  0Q2p`l�+���x PNy�7��7 �����8��@�uj�ԩE<�N��[ZZbƌEl
+�o��a�bΜ9V�B�<��Cq�m����  L��K��ܹsc�ڵ@����� %��t~��_v wyoڴi�(�:�S��"Cww����ғQ�m��*'|����+p�r�����㏏SO=5  `��q�q��w ����rZ�lY<�� 0ގ9� Hw�c�Ϝ93Z[[c�����2F޵kW�ᒻLlܸ1:;;(�\�r����E]� �������Q�����ǒ%K������;��N  ���ӧ�G I�u,�����"L~'s�̉U�V��Ν;��=�D8�rq͖-[bƌ�C.l9��s�_�bq�  㭧���=,w��r9�]�Pk֬��/�8  &BNo�kx I�unڴi5�='��
3�<��!�ܛ����9@9<���q�7���  �����8��c�������e�����@�۱cG�u�Y144  �-��E��(�;Թ������szjNq_�n]@ʉf�6mrъ	�����c��'P��ַ��㏏���}  㭷�W�0F=�P�޽�5<���+�^ ���q{F� �\}�:�Ӑ3^~�ߛa髯�j�f��6Į]�&J>���].�ill�������.���>:�<��  �����_ T.��l��zj P�����.���� �Dhhh��K����PӦM;�)�---1k֬�k�ΝEd<220�r�SNrϭ�r�/��q�9�X� ��:��b�ԩ�cǎ �r}}}w�:�����UW]  e���E��7�;�@{{�A��#���XN�ٴi�)�L��l�3f���y晸�������  �K��'�|r<���@�2p��>�³�>�� 0QLo�G�%���S�L)&#��\�A|^��<2hϰ�םj��{Nr��/���8����p  �x���������b��̙3����/���X�jU  L�������
�}	ܡ$u�{n=G9�ƍMb����ewww�@(�K.�$�:�(+� 7�_|��@�FFF����|�#@����;c��� 0��D1%���6p�={v����K ��g��&'��_�����;v�/~�q�ƬY�  ��?��
��C �\__����<��cq�� �Djmm���ܡ$�N�ZLA޽{�;�ކ���3gN�Y�&�_CCC�iӦ""�j5�À�<^}��8�s�_�B455  N����3ό�~��@�L���֭+��� L���n�!p w(���A����}�ڵ.dԩ�>غuk@-ȉι�̙3(��t�5��g>�  �í��W�0F�V��իW��P�r��/}�K} �p�agK�,	��C�J��'�]�k��ԏ���bv�PK���9���(���?�g}���я~4  �p����������� j�E]�>�l  L�E�EKKK ��J$O
�L��w�>���G����cϞ=A�۵kWlذ�T~j���@���;P�]vYqa���  8\�Ν[L�z��������	�j���?�� `2,]�4 ގ�J�P��O�:5fΜiK�:�m۶"�X�Z�߿�H���;��8�o��o�.�ٳg  .9�]�069�=wu���<��#q�u� �d�3f���#p��9��=�w�{mۼysԃ܁`�ƍ���@9����/}�8r  82p�����mٲ%�|��8���ڱv����\,R ��w\ ���LKKK477Q���ӣ���� NmɋR�ر#����t.��&�rț��\sM���i  ��p��(w�� T.���jG�����?_�g ��ztww�;�C	��������9���^jG.`ذaC1��Q�J�!B{{{ ���|'�,Y��[�  0Vy},��Gy$ �\___�ɟ�I P����]t��� ��:��c�`ܡ�5p���5k���w&WN^ȯo^��z�iӦbG�<�r��+�����  ���^�;�=��c144d@������� ��2u��8ꨣ�`ܡ�2mii��;w��ohh(���ȝ��	�dk(�\đ;̙3'�������_�B1e���3  `,2p���+���{��~8>�� �k�ʕq�7 �d:�c���1 ��J*��l��2 ]�vm�gdd$6n�;v�(�|N������b1P��1�9�ė��%�[  �O<1fΜY �r���w�*�C��j�O �,��n� K�%��{b+�H׭[T����S�->��r�N��f�
�~���UW]��  P���v����� �r}}}@uڶm[�u�Y�u��  �L�-���� 8Xw(�)S�'۷o?�?s�Gī��{��	�C^��5����lsss���P��sO����?��  �J���
�������[� ;w�� �z���/�0^x�  �Lq�����C���C	�3���(��3�m�{ٴiS�x���%�r����㨣��w���  ��������O}�S@���7�?��O `�͛7/f̘ �B�%���3V?���9�]�>��������vx�|.۸qc̙3�x� �oxx8�>��8����>  �\0�`��X�zu P9�;@u���o�9  ��q� �J�%�hkkkl۶��L[[[̜9S\=I��u�1�?��������ܻ���� @�˅w_���s�)^' �P����w� T.C�@���{���+_�J��� �d�~���3 ��Jn�������.p�x���裏�������/����ܹ36m��g���{�"p�����7^' �`���
��(�����}����ٲeK1dhh(  ����@��Pr���Ev(+�g̘Q�9F&�ܹsc޼yo�~�t��x饗L_�������6mZ �bŊ��7���_��  �Cq�g��1 �j�����I�{���җ�/��r  T����@%�PrL����֭[�����>_MMM�hѢ�N�ί[Nq�m��ʝ&2roii	����oőG���'  V���w�;�x� �r���������۳gO\|����� @�8���4��P܁b���\g4�s��`|L�:5�>��"d?�c�=6V�Ze��G^�ͭ������"@9\q�1��x�{�  p�zzz� c�r��رcGqm��u뭷�����;  �Ekkk1��Rw ��ۋ�sxx���L���ht����ᗓÖ,Y�Qn��,��^z)�����ϙ3Ǫ`(�<��ۿ����W�R��  p0z{{cٲe@�r �#�<R,`����?�o�1  ��ҥK���1 *%p
�oٲ��L�k׮�ݻw��ܹsc޼y��v>���wؿ]�v���@tttPyN���>�;８>}z  �;�������P P���>�;�z���.p� �*9г��9^y���)S�?� C��M�vȁ{�����*"w�.O�rk�ٳgҟ3��ٶmۢ���x��aժUq�Yg�����	  ����v�i����� T���? ���m^�ܾ}{  T���r�g���{�����=�� ��@������u{www�[�.���T.��ܚ'��8��c����lӦM���ԩS(��<.������>  �Nz{{� c���O�eggg 0~v��_����^ �j�=فd۔}Z9�po9lu�i��S�~�a<P.w�9�8�C�'y�z���AefΜK�,�*��B{����;ظqc�Fʪ_(���//^����  ����; c��>���'��122�{n<��3 Pm�#�0�y��s���؛��PNw�ӧO?��=y��D��ݜ9s�0�p�2<��b����������|�Y��lٲ�|���'  �@�9昘;wn�]�6 �\__��`]w�u�s- @5:�#���vS߳���s�������s"<P���F_��]�N��̚5+���'W�-:�۴������/����ڵ���n�d(�\�r�y�S�r�  8�3�<3�� �r�K��ػ ��;��iz_�}�i�}_T�[MY�$S��8��TRIj��1�$�1"P\�ȠY�4f�h2�hH$�����,���@��;����_�{��Uu�D�M�{��|����U�V��'�  �����R,Y��l�����-��z�`���
�C���ڍ{�ZQ	�w��(Y#XFFF�?�E]����GKK�����5@0�I������{�U^^�   ����?� <���ڽ{�*** ����~[K�.  �WE��=���k|7VLj���޻��xw ���隍�t[O��;;���� |2�ڢ~�N�����ڻw� ��]���Ijj� �m�/\�Pw�q���   >����ӵ1 ��Y�;w ��C���M�R  �EV�����D`k��� |�^�>����x[7;�|��BKKK;���)))!�~���.|mC�q-�v
��ف��d�۶ms-�g�f   SPP��V�o�. @�,���/~Q ���DZ�N���(   ��ܘ�:uJmmm��Q���`���9���, c-�����ĉ��Yxn����Ϗ��gm����X �foLjjjTTTD���k׺Cg����.   ࣪���@�^y��2�5 �Z�~���
  ��,�ԧO��ݛ�-Sgy������{W �����;����1��j�Ϟ*--ջ�+��nVl��ci���ڷo-�@7��)kr��! ���㏻	���    ���N���{L ��ن��o��	& �|P�7o  ��Y^,ȥ��O����w��Yн+����@8p~�|��pX ;�1w999JOO��o�9�p{<nH�d�^�]�v	������k^vv� �ҥK]��5t   ]&N���VZ[[ ݆�@���O��   ����yyy��Y��eR��A]��z�=k[��a��U�wSRR�={�(Ȭ�_�~q=����n�� �Ϯy��!--M ����n�v�m6l�    c�r�ƍ�ƍ �ܯ��: zn���Z�|�   ����8����j}oooWAA� |w geO;!J8:777�-Wv�ֿO�x�f����s�N���Z���`�������{�Q߾}   ��C� ³e���׻&: @�m޼Y�/v�'   /�lE�찤��+))I >���O�����������t����$v�6h� �~����ݻם�p~�X\SS�0���K ����A��z���A=   `�ԩ ��&���꫺�+ �+�Z�`� @B�A��|��#��YP;�����y�L�:##C�5�K���]���;�{l�خ}���v�bM��~��d  �`���t��4  t6l � �dk�?�����,   ���q�#tv8���w ���ѩ��jmm���Z����:tH~g�������Dkq߳g�hq����E��������ؾ}���N�r�-��  8[ۚ2e�V�\) @�^|�E ���$�͛���Z  $���B�T�d��	���8'{!%�n�F�ȑ#����FYY�JJJ�e�{�v!�m۶	@��b���pZ��_~Y=����?�S   ���*� &+�9x���� 8���6-X�@  @"����b!<�����8���L7�����=�X;��r��VTT$̍�}����a �����4��b�I4�^{�   \p �oÆ���?/ �ǝ:uJw�}��l�"  �DQPP@�"L)))���q�pNv�.##C'N����ޱc�|��nm�ֈ�H7v�ࢋ.��o�- �g�{�?v=�����f���*   �l]k����4  :� �ɖ-[����   ���>+�pn������p��z�������i��	t����{�n�<yR �����ֺk��.K�,Q~~�&L�    ���p����K��� �!������SO	   �Xv"���\p�����s#�༬���Cma�jq��De7eee*))Q��?Ð!C��o@ϴ�����A999v�h�"�q�<x�   <p���- @��e��5J �����z��  �H,{���)�HKKsY< �F�@�ة�����>699ٝ�;z������8���l%���r�ڵ�m( 虦�&w=KOO��hnnּy�t��2j   �&N��ֆ::: ݆�����o���sS$  Inn�RSS����tw �N�ݔ����D[�� kEE�on��$�СC�ꫯ
@���չ`��Gmm��Ν�����   �}���=z�^{�5 Bg������۳g�.\���v  $
��׫W/edd��p�-洐wkkkHo�Pkq��{����Ӏ܍���a;QiA] =c�tjjjTTT�k�sۿ��/Z�H�   KUUw ��͛u��	wp �����nZ�]  MNN�����VP
����6kq5�nJJJ"�n7eee������JmܸQ z���ӵ9ۡ ��}�v��'?��ٳ9�   p衇 ]GG�6mڤK/�T DMMM�3g��  ���P����!�����5[�q(RRR\ ��	�*))It�����������OCC�� >nݺu����/]����  ��#G�O�>���  t6l � ���ڴ`��۷O   �(;;��\���̴p���6k*��k���'$Mv1h� ���)��Bz Bc��޽{3��?��������   ��&6q�D=��� ��� 46vѢEz��  ��ho��ہ�!��G�6�������幐��XsEE�۰���\����ȑ#k��� ,O?��{-���k   ����"� aڽ{�[��ui +�Z�d�^~�e  $*ˊ��M��� z��ͭ����#��a�׵���iq�������HMee������F} �ώ�)**
� ��կ~��>���	   �fw @�6nܨ�~��� X�l�V�Z%  �Df�*��+s�����cv*���.䏷�>}���9"!))Ip�A�����}�����/j!����@����v�if̘!   �W�~�T^^�
 �iÆ��c�=�+V   �Y�8�����w =f������Z�KKK���HMMՠA�\�>������өS� 4mmmjhhp�w ��~�{�JOO��ɓ   ���'�|R ��Y���K3��=�����o+  �DG{{d�{����� z̚�-�����X�Z�srr4p�@����ߋ/�P�w��Н8qB��ɼ)�&9,Z�H���רQ�   "� �=�;v�� ��^?���  �謽�JP>ko����g�����p7���{II�;]�MÇ2DP{{� ��&S���[))),6���t<x�   �?S�LqmKL���X�;w ~d׷ŋ�m�5  @$Y��a9; =G�@H��8�=k�6���E���0@�����Y���A��m�6�-Z��֪���)@ �<yR���ӝwީ�}�
   �b�U#F��[o�% @�6nܨ/�� ?y�7ܺ�M{  Ht��L�g��$�!� $րn����[�z�����p�z|2{����v3?t�xm!����E d?�7�|���.   �RUUE� ´i�&�����{ ���۷k�LJ  �ay.D��f w !�D��N����G����;M8p�@������!C�h������6w]cjLǎ�-�������   �����e� ������k�
 �n�޽�;w.R  �7ho�+E�����p��*�;���{QQ����iP�~��i׮]jjj��<yR��ɼY�СC���[u�wp   �1cƸ��'N ��7p���b޼yjll  �_���
�a눽z���p�r���>Gzz�k9������d��(??_�{��W^yE �gS.,�n�� ��ݻ�h����k   _�޽5a��Y�F ��mذA7�p�  Qپ�Mq<z��   ��2\}��"#++K BG�@X�YMM�N�>�������iEE���Д�����}���ϒM�HJJ��y��7�h�"��G?�:   �S�N%� aھ}�+�)(( $��:w�\8p@   ~B{{�XZZZ� ���;����755��y�N ���nm�tMZ���õn�:ߩS�\Ƚ���MI </���/^��3gr   ��iӦ	 +�����\s�  �����p���+   ?��Vnn����#
 l,7�n���Bnq�v���rBcb7�v*�������vw}�� \�?��RSSu�u�q�  ��lz�M�;r�  �۸q#w 	���C��~��n�*   ���=rl?��;>� �fa��������yl,KO[��`�����"kذan�6� >�F��*�z ����?�I3���7  ��6u�T=��S �nÆ�Da�Z��mڴI   ~c���Bd�󙔔$ �!� "��YMMM؟�Nv���B�֘���!D��p���}��	@d���­v0@0=����:�}M   H\� |���ڵk�$ ���N�}��Z�v�   ���ZL���ہ� � "셹��6�o;�����>��~���6dDϐ!Ct��A�p 2��VTT�i] ����?�_	�  $�iӦ�W�^�� :kq'����~����'�  |+--����,e�@dp��g/�'N��s٩����O��_�~�����ͅ;v@d�b�M��k�1 �,�n�����M   H<V�`� ۶m  t7n�1 ϲ��|P�W�  �_��ۗ�Begg@dp1���������n7S���WAA�;��������" �����q���\˗/W�޽�/��/  @⩪�"� az�W��֦����X�����ʕ+  �WVfJ{{deff
@dp1LONNv��p���}���>�5�3�%�lt�СC�y�f�;4��Ԥ��,��{�����g   �L�:U���/ ]ss��z�-M�0A ��?�ӟ�T�>���6M�JЎ=*  9��B��o˸�� "ʂ�m^Ejj����TSS�N�Y��N���Ӟ={���  �c?S��Ʈy ��BQ�A���^   Hƴ�s��� �nÆ�xʣ�>�g�yF�+�6m���k�j�޽  �<VNN�9�EZ@D�����QZZ�,����~E���?b���  ��PPaa!�x���M3�Ts�5�   �!%%E�Ǐg� �d��뮻N ��<�|�I�l�r��骨�p���K.q�r  |}��"'))�����T "����ĉa.k�0`��6����X���9�N�r�*���8��|����&�  �8�N�J� ´e���׫O�>�x�կ~E��C>n��g_|��[ٿ�  @h���i�0{>�| �E�@��MP$���Ç��ѣi��w��=??_ ��+�ޫW/��?��   �}UUUZ�x�  ����+���+��R /�?��~���`k���~�24�w�^z�֬YC� ����
�Ł ������4%''���]����$�����Ң��FwH@pY�}�ҥJII��_.   x�СC�Ի�Ǐ :��A�@���������G��� {������r ��rrrcGXzz����,� ��n����c�t�� "�����
.k��������3f   �ec��L��?�� �n����xX�b��-[&xCw���o	� �3eeeBdQdDw Qa���:�B
�F���k۶myv8���H�{s������^��[UU%   x�ԩS	�@�:��_�~�XY�r%�v�I���C� �����UFF�9VZ�s
D�) Q���}��	��}�����Y "���Ԩ���-����N�q����]+(   ��� 6l���@,<��sz��)��P���XB�  �_ii�Y���C�@��8w�����J����yn
F~~� �]-Z���G�4i�   �=��Ū����ݻ w ��j�*-Y��MQD�پ�3�A� ������t!r.��eee	@tp5iiiJIIQ[[��?���ڳg������566r����۵p�B�t�M��  x�ݧp�����n��M��h�p�<@��#"n���"� ��Y���L�,;0л7\ Z��U�<~���OÇ���� :,�no�8E���o��v͜9S�_~�   �-p��� ���9�]G�a� ���+W��$�����sr �����\Q)"��B ������L��ֲP�S�����{�' �aS���9���O�w�}:}�����
  �;&M��$C �&�:u��3���@����C=Ğ�GD#����M� ����ĥ��BdQVDI) Qer�b����WWW�ѱ "ς�555*,,t�T �fp����6\y�  �7�f֨Q��i�& >,##C'N�e�]��p�XZ�b��-[���6�����|= � ��Yyejj�Y���G�@��:w��܊�
�ܹS �����M�((( t��[ZZ��OZ   ����*� ����C�=��n�v���'�|R�<����w!�  ���b�kVV� D�I ���3�I���V��.��"<xP���vmhh`d3 �ڦ~�ӟ�	*���g  ������>( "*vڧM��F? Ox�'�裏
��p{B� ��+**r�-D�M*�{ �E�@LX�;w������J����=MMMJNNv� �B���/ܯ����  ��1b������z�����iҤI.�>}�tx������`�<.��2������&� *�򔔔�g98 �G�@Ldff���ֵ��maϞ=����豟1[��; t��[ZZt��
   �c�{��/ ��Mi7nܙ��aÆ��� �E��կ����F��x�ۻr Qqq�{FdYV#--M ��+����nIJ���YSً/�( �ca֚�7J�d�ئ]ss���   �SUUE��oX����g̘�o���u�~�l�2�X�B�/�ۻt��_x�8p@  ���[� �G{;;�Č��744��%�����M��
@��4��QPP  ���O�_	�  �ϴi� ��֚&L��B�\r�k��D�5�𩧞���u��ԧTZZ*�����"� �;{�MJJ"�
^333 6��[İ-�.
��Ѵ�v\ �������� �X��ԩS��W�*   �^߾}կ_?�2 ��׏;���ak��Y ����?��O��3����p{B�  ���[���B�Y���@�pS��N���lSd���ھ}� DWSS�[$��� t������}�[�"�   UUUg�� ��X�����L�}���.�  ���x��Z�J�/�ۻr �YYY{�Qb�7 �C�@LY�5:::�4h�����a ��땜�� ���g�u�{�]w�۬  @�p�%���g�S�LQ�>} ~a�_�/�_���!�ޅ�; ����ӕ��'D^jj�{ �� b�N����
�e�xl��k��& �e�WkjjTTTD����\���J�   �&O���,p �f%3�G�v�v�Y	 �Qgg����Y�F��D
�w!� ��ۣ'''G b��;�����R]]�e¿���={�p��[ȷ�{AAoV|���[ZZ4s�Lw    �g�#F��[o�% �6�UVV�ii�8q���٤��K/�����n�B� ����L��g�� b�. 1g/�vS���$�ۨQ��v�Z3 1��֦��ް������:q�~��*%%E   ��iӦp5���g�v��R ���V-Z�H�����n�B� �VD��B���#� .llw���s����o�>�>�&''sr�Ǽ��˚3g��Ν�5   ����_�B 	����<y��O�>=�� [���-[��`���/�\%%%Jt�� ���9~��[�@�p�����Z�oÆ��Ç]�4�諯�wʴ4����~[7�x��ϟ���|   zƌ�&Z z��uƏ�����҅�  �jkk]yî]�o�+��BEEE�B� �DE{{�XyXRR� �w qc��=*��-n:���@��>}Z555nA�7Y >jϞ=.�p�B�   ��ޏM�0Ak֬ tGyy��@����! �����u�-��СC�7��ߕW^���B�!w @����Szz����C�@����0;;;0`�[ �����;u�k�)((p� ��l�ʬY��`�8P   ����*� >����A�_r�%*.. ����߯9s��رc�7�9�ޅ�;  ����	�a���� >��+;�F���,`;b����mmm���Wnn� ����C͛7ύ�  @�M�6M ��6�ǎ{��}ذa �y�رCs��UCC��A�w!� H�����*D��@|pWv#`�ӧO�f#�l���� 6N�<��i�l]��=F�-   D�M�)))ё#G x,g����Ǐw�o ��y�7�p�B577��p{B�  /��)�ۣǞ߬�,�� �*))I:q��Çw���lc��l�8;s뭷j֬Y�>}�   Yj}ꩧ ,�g?���2e����# @Ͻ��KZ�h����ob��!w �WY�B���?����L^�+�����!�6iȐ!ںu� ĆMȨ��QQQ�;T e�w�q����z]}��  @�TUUp|��[l"VWK�|  ³z�j�������!���.]!����oL� x��-�������"� �,�l���V��***\�Acc� �ƩS�\���9a�l�:���C���O�$   D��-c�[ ��<WVV�	�O�8��< ���������s�<���W]u�


tvp�e�r xBYYwQd��>@|������`�p�#�q�F�kh���S^^� �ll�òe�ܵ�+_��   ���\:T�� $����3�v;�B� D�O<�G}T���G� �iii�>G��o ��233U[[˸������R>|X b���Y)))� ��6�z�o|�m�    <�%�$;�2y�d��;m�4׊ ���҅+V�a{	W^y%ṳ�5�3f�^ � �;�����C~����x��xeee���^kq?z�(���묍�NMM |�g�yF'O��w��]�  �����_
�7�{��`A5{TVVr� b����,Y�U�V	�A�������;  �Y<''G���� ��3�����55��������}�v�-��QTTDh�9�^�Z'N���ٳ9  ���ǻ����V�k���v{L�>�iw mmmZ�h�^~�e�;,�~�UW)??_87B� �x`�Xtفw+h��x�5
gdd� ��������S�N���F����.pN/���n��f͝;�6  �YHh	Z�~� ć��&N���_|�JJJ ����&-X�@o����v(���yyyB�r Ē�Fs@;�,��T7�;��Nv�)5j�6n�( ���ޮ��:��׶m����}O?��]�!   z�B�܁�IKK�رcϴ�6�C� �Ǐwe
{����p{�� b������W�{�)����; O��F6�5H����{O b���Y��Ɍ�p^��~��z�>|�   �3UUU=V�QYYy&�>~�x7= �-j�7o��;&x����+	����;  ڊ��x�e����ݛ8-�%�D�;w��Q!8F���[.�n�� �\5g�͞=[�'O   �oȐ!*((p�� "Ê3,�~饗�G�>} �͛7k�:y����#��;  Z�5���D�.���!��s233U[[K�9@,Xk�[�n�سk�m
s�����h���ַ��k��F   �ql���>�� �ƚ�ƌs����R �8V�^�ŋ���1��#��;  JKK�ˏ2kǷ{# ��'egg��%�����-�X�4��:u�jjj�X3] ���5c�ҥ:r䈾��/s�   �&�@����K���g�&LpS�  �eŊz��ݚ��\W]u�rss�Ȳ��M���_��Ç �pX����]L����; O��{]]�N�>-���F�����@�Ys�,��� t�O<���p�n�   �VUU��?X�>Yyy��@����:1  1Y��g?���y��[�G���~�S�"� [߾})��2����� �!������6/h�����O��kiiQSS���� ����ϻ���7���  �yXۖM�۵k� ��ҦL�r&�n� ����ޮ{�Wk׮��p{�r �+==��������Q�x��i�
��Ç���Zmmm{v��]m� ����_׬Y�4�|   ����d֊6t��3-�&Mb" ����-X�@[�l��p{�r �æ���.{~) ���; �JNNv�O�<)GJJ���z뭷 >���TXX�^�;��ݫٳgk޼yn   ���˗/$�!�h�>}�233 �'�Ν;W���\���J��q@� 
k�bPD���9xx�% �f7l܃g��:p�����S�N���ƅ�{��% �ۜ��~�9s�h�ȑ  ��Y[��gr�,??_'Nt���/�X%%% �ߞ={\����シX�ݚ����#�!w @OX��G�Y.�wp�i6*�M�౛�Q�Fiݺu:}�� �^GG�;db�� �]MMM��[���_�\r�   �a.=z�^}�U~����q�Ɲii6l#� `^{�5-Z���*�����W_M�r tWQQ��K!�l�.99Y ���; ϳ�rǎ��Z$��}�޽---jlld�@������;�ԑ#G���^   ����*�Hx�Ҍ3\�}��� L�V�Ғ%K���)xKff�kng��;� �'))�Ih1B{;�}�x�-���ֲ0@��d�8���۩eN��	����#����^_��WԫW/  �}^�t��DRPP�	&����^z�k� `���z��Ǚ��A�۽��; �\����k���[�; o�j��l��-����	�b7�#F�ЦM� ~쐑m\�F@O����סC�����E"  ����:lr�����ǌ���>|�  �b�Tv`�����=�۽��; �l�t���}�H)Hvca�~4@��N-..Vuu� ć]{kjjTXXH3�۰a�f͚��s�(  ����U�'O֪U�x������<h��v�� �G555���o��͛�!ܞ8� >���\����$eee	��p��n.��5j������F ������m$9 �Ԟ={���}Os���СC  tUUU�w�q�h�GNN�  8�Λ7O��p{��
��^�ZG�  ������a��\  �G�@°9��d#�-�u�V����V544��@H���ٳu�7�M  � ��;k�8q�.��2h� �[�l�m���&.�{�'.�_~��� �,l�{�ذ��% qp�0l$�m<yR���
<xЅkď����<��joo׽�ޫC��_�"�   �������k����ŦbZiDWC���-@ @O=��sZ�t���	�p��W_�a#1r�`�)��ǆ�/�z	���J&��b��܃�p�G�֋/��ӧO@���չ�V�@O������]�k�̙JII  @Y�;wD�5�uڧM�F� [�y����Z��p�r�`��uYY�L�w 	%--M���jmm�'77W�޽{ ~lS���FEEE�ի�  k֬�ѣGu�-���x  ������~�;����ӤI�\�}���*--  �����&�_�^�&���C� ����3m-6222(�WG 	�O�>�������f�6�-�����w������u��  T��~��hΜ9���  $J��.{t���7�LK�����C  "�
N�ϟ��;w
�d������p�r��)�V*�ؠ�H<�$;Qgo�;::�س3kY����y�ܾ�#F�ЦM� �l�FCCo���',�~�7j���  ���l����o
8���rf�1c�k��p  �e׮].�~��1����!w �~��qh=F�0��<$� ����?.�V�^������t��-�n��X+++SII	:�455��V;| �jnnւ���]���g  ӦM#����ii&Lp��K.�D���  ֭[����'���d�$���j����; ��T��b��HL�$$�ѫ��c�s%''��4����n�G�[��ȑ#�!�������w׆^ ��N�:�����ڷo����o)))I   ~gm�v�`����cǺ@�=�F�  �V�X��~ح�������� � �d��6��Aa���HHv�grG�ٍ^aa�kp��x��[���!C�u�V��ӧO����Mx8�u zb�ʕ����M7��b  �ѣG+33S'N����;WVV�	��?^)))  ��۵d�=����544��s-�]��o���lr{`�C{;���HXp��`V"z�F///��}<[�+**t��!�� @|�D���Z���� l�6mҬY�4g����
  ��lj�ĉ��/�f�l]��)S���
 �+����(J0�܃��; �����;�|gee	@b"� au݄466
�gMR��ޝS��jq��1c�v�Z: �����٤	{���̙35{�l�7N   ~UUUE�݇lM��-�>c�4H  x���,X� .�;!��!� �`����d!6�<��> qp��rrr���D�9��f�����7��lq���A���
@��8q�];� � �ܹs�կ~U����  �GpGⳲ����3-���o!$  �襗^�=�ܣ�'O
���{�r�Ė�����"!6,�nw ���U 	�B��`�\���i7Զ)��jq7C�q��k�_}}�[dMII ����S���/�}�v}�;�q�   ~2p�@��E{j�)//?h�6m#� �g�QO>��{�1�:uJH|�܃��; $�~���&CnOJJ��E�@³o�ѧO������lq�R��a��?�$���Uaa!oD����78p@7�|�JJJ  �'�^�b��mV�0y�d���>}�;�  @�hnn���߯u��	�B�=x�@�5�7!6ho���;��g�jk�lmmBcm�D�����ĳŽ��@о}� ��q�B����)t ����j�̙�馛4f�  �EUUw��d�Ǐ?��^YY�㩇  x�{ｧ�n�M{����B���_t�UW��S�!w H�_޷o_!v,����, ���; _�����j��l��ZP#qc�w3|�p�� ^�?�kkkS}}�;� �b�us��ї��%}�_  �XxڂӧN�⫼��L��Z�333 @"{��Wu��w���I𷺺:�Z���{�r��`�+�D�Ж�w �`'�Q��>[�***RRRR�>g<[�mg�ȑn��7�<y��!  �lJģ�>��{����w��   ���S��w�yG�-�<6a�h��KT\\,  �����z��'��c�q�.@,�nM�W^y%!�� � �f{XpG��=
  ��7��ݱcǄ����vx�����R��W���Y۲��	��4۴ٷo�n��wh   �UUUp�[�;v왖�aÆ�Q�  �Iss���~�[�N���ZB�C� ��&���>�N�>}���k�V����ن]aaaT۔���nF���Ǐ���] �Ϛ�jjj">1 ̻ﾫ�~���馛4z�h  $*�۔D�m"WVV�	��?��  _�����w.B��C� �'++��g;�擞�. �@��oXp�Z�-D���`��Y��(�x��۟o���ڼy� x�������@���׻�/}�K���   �D4nܸ��������0��34e���  ��i�&�u�]jjj@�=x��w؞x�~���b�� |�N?Z����S�0[��e{r�[����C��رc�6U�&m���	 "�������?���o��  �DbS�.�~�z�g222�4���v+>   hV�X��~ؕ� ]�OW����Wuu�  �a���c�^333�?���+6r8;;�(�w�l��������f���Y�2j�(�Y�����5�B��-+W�t#�o��f�  ��SUUE��l����L�}�ĉp ��,Y�ąY��!�<vo|�Wr�8��pii�[���Ê/ ߱0wCCz��-�*�g���C��֭[�;l҆��OMM D����p��я~�O   ���8����3�v{��� ���ۅj�Ν΅�{�r���۷�����ر�;++K ���; ߱'�i��{���[qqq\���l#�O�<�����BG�QMM� x�-��X6���{�馛�����k  �.��"��Z����j���.�>m�4���	  ��믿�;�S�������-�l!w
h���; Ğ1Z%b��P���p�K6v��N�>� �E)�{!8��������3Fk֬Qgg� x�Mٰ�7x�	 ZlD�ҥK�e�}��ߦ�
  x��?�2e��}�Y��c�$�3f��M�"  �a���?�A�>�(ӌ�c�.���N�=�@l��׏����#&��D��/ن���ljjR�؟�K����d��~�ĉ�}��2D�� x�O����A ��իWkǎ��}���  �2k,J������y�1}�t��  >�M�}���v�Z�"�<�� 6


\>�e��$ �D��oY�������n�v�ln����]���4h�>�´ ��&<�A���,@48p@�f����_�A  �ʂ޶���5-�=q�Dh���URR"  �=���-Z��:�prB� ]�.++b���ho���; ߲�dzz�V��5�)--M^�^mll���`7�cǎ՚5k�	xLCC��N�� ��P�]wݥ͛7������  �k����bKt�Ve�1]-�Æc� �9�.]�T���"��{�r���۷���FlY��2S ���| �fm�~���������-�^455ŵ}�B�C�Ѷm��[jkkUXX(¦ ba�ʕڹs�n��&���
  �k,��wk+���<h?~�[�  �ikk��~�3��O�܃��; D��nĖ�(X	�� �k�c7�---���Lw���W�Xb''��9���w����w�d[H�i�� ,����|G3g�Դi�  �%UUUZ�|���MY���K/u6 ��hѢEڻw��h"�<�o��O}ʅ܏;& @�lo{���qǁ�\���w �g�j~�ۍq^^�rrr�H�{����w{�ƌ�u�ֹ@- ����pM�����X�I?��~�>���k_��`  �3&M��ϭ��k�����JWK����  "��_������)��B��c�7���	�@�lo��)[���@���٦�-Ĵ���lԳ5۟+�Xh�B��nO�����w��! �b�����ik �;x��SOi��ݺ���!B  �x���"�W���������3��	&(99Y   ������#���
 �,��׿�U�_~�?���@x,ӷo_!�222�D ��O9�@�S{���Jt��P\\��7i.��x��2DG�QCC� x��\�u� +o������z͚5Kcǎ  @�Y�<^����3����*egg  D�ѣGu�wh۶m����^���{�r����IoB�q���+ ��@ ��=��u�.�3�֬D���^WWׯ��Yںu�\s+ o���u�*X Kvr뭷��k�տ��&�}  Hl,_�tiL~/+��2eʙ@;�c  ���/�����'� �7B��C� z.33S���B�Y~��@0��Qg2�Ⱦ���<�EW�{ggg\�{^��;w
�����ꇃ= �ݟ,_�\;v�����}eee	   ��ڨ�Q`C�=��>i�$��  @l�:�o~���׿���[���B�z&@�����P����WĞe} w �a�'mC���]��B��`���.?�?��ܭ�9ކ���j544��ttt��6'�ă5�]������_   �f�'�'O�s�=��gc���ӧOwke   ~l�����o�!��,�nagB��A� �Ǐ9�D������T� �N�%ʛq[(*..�킑�-T�w�,;v�֭[G;
�A---n�Cvv�  �lo�����W������  Ĝ��C��a�'��q�����D  �,�~�=�x�8B��C� έw��*++�æ� %++�5bX+��edd���Ѕ���bv�y���x).l�Ei����=p��s;� �f�~������_�7���   beڴi��o��jܸqgZڇ�=  <Ɗv~���j���� aX�}��պ���	�!w �d����u���l�� ,����{!T�I�����SX#�W����������#GT__/ �cMF6��N�@<lܸQ����5s�LM�0A   �`�`�����������3f�@����]  x��q�w�}ڴi��DS]]M�=`���Y�fP�<^D{;<$� ���-��w;�i����$vj�b�f�f�r�v�Zuvv
���>}Z555��n��l#z�ܹ��g>��}�kJJJ  @�Y�{W�������@���^�  �۰a�/^�J�DE�=x���Y��J�����. �B�@ ��丠�WX#qIII �,�oc�Z[[����ӶC��֭[�{�`��K-� �bn�z�)���;���UZZ*  �h���?���
j8p�  @�hoo�#�<���~ڭ) ���{�r��Y�'--M���`"� ��Zܽ��m'�m+ȍ�v#z��ay�m9r�S  ���ihhp�  ��o߮�|�;������.�L   �2z�h�   ��&��u�]ڽ{� ?!�<���]-�����.� �FY8Қ��ɂ�4˝r������x)���رc�f���{���ܢ9ob��ɓ'u��w��W_�u�]Gs     p,�t�ROL����{�rd���tie����
@0pXp��x��[�ڂ�YYY�����u��!O�����Pee��~�m𦺺:��ݛ�s �`�:;w�ԍ7ި�
     Scc�x��_�^��rB���ػ �����/�]��w9wa9E�[4��11f4j��I�1G�ɴ�N:�iڙN3���*i�5���$A�{�A#�D\�c��ҟ1V�cw����|��f�ic�?�w|>���D��E���B|�{�5< ���@dYdn�-��I�{�V߾}���,��-|������>�8��Ο?/ ���0���*,,�< /�:uJ���������ԧ>�>k    ��8|���魼�\@T�G�;�(�}h�ގ�az;m� "-6Ž���G��RRR\�i�;�/�`�����w3a�m޼Y����������݈ >���/�k���o}�[�0%     7[�|�g���O��~�"��!r`xe1� �;�H�Ӗ���w��0/-11��s�C>�	�_��� ����ٽf�k9 �b�Νz衇�D�)S�     ���kS�<( �b��E϶߇�#rv����۷�?Lo�7 ���S�{��������egg���ޛ)'����:Q[��'{ͰsNo���0��@w�q����/s�     !�m�6=��n}�#w���ܣ��@XY�c���� �* D^wNq���Ntre��f=5U�rM�8Q�7ov�������]}��� |��٩�+W�رc��w�����     [SS��x�	�Y�F ��E�6mҼy��#��@(==]��	 |�  u�w��-ngZ畳�uuujoo�laf���ڳg� ��"���J��K ���������~��     �[o�����ɓ'���9s��=bb���u�TQQ! 2{�8p�?6Ԏ �& @]?�=33Syyy��"\9�疓���H�~��To��� ���TUU)??_ ���/jѢEڽ{����     ���/詧�Rkk� \�{�X�`�"w �g]��=4 1|� ���S�ca6W�\;;$`χO�cƌq2������f����:�[;w�ԛo���~X�f�     ��ٳg����D���� \�X�~��7s�uD�:�}����� ދ� ��������ȫa3���JII�Fnn�Ν;'_؄�I�&i������ ?544�/�iii �����ќ9s\螑�!     ������g?��������}�ƍD�B� ��}���H�/�x/w x��^WWw�S��z߾}�b��Y�j��������Ǐ��,��d{} _����ȑ#��������     ����J�=��v��! ׆�=z��р�5ď��3
�{Qb�{آʕNq�W����ի���,(��/�\w�u�p��UO����ۄ*((`���춚���wܡ/~�,�    g[�nuq{mm� t"��!r$���n_񕓓# x/w x�˝�nA�}��z���L444���O�4�M]moo ?��E�B�;;��r�J8p@���w4|�p    ����ب_��Z�z� t="��!r��\\\�~r�� (��x?w x�˙�n�?���JII��Mq��e��|a�m�����_---n��� �[o���{�G��{�     ������������
��X�i�&͛7��="����ڟ��T!���������w�޷o_%&��S쟵='�:tC���������;񝖖& ��>�l�2�ݻW�w��
     t�a��W�X�7��eeeD�C��W��Կ!��yHOO �u& |���n�


��(l�r}}���|2a�m޼Y����/{=��2�� �������7��/|��ԧ>��O     �ؑ#G���X�O���E�=D� |T\\����������x�w�sss��HHHp�Aee�|����q����W_ uvv���b�E
 A��ܬŋ�i���ַ���'     pml����?���zʻ�:@��G�; �X�c]�������!p���n��Mm�U���6-}���:{��[��/;�TUU���|&!�}�����C=�9s�     \��'O���'N���#r�"w >���A�	���v �B� �`AuFF����?�)�s���7�Ǐw��ŋ�_---����F �S[[�������]�n�u     ��W�\�%K�x7D�:"��!ro���_rr2�F\�; \�-�����p������&�$11Q�'O�����B9 �A[<MOO ��ݻ]��7�7�?�     ��Y<�ӟ�To�� ��~O7oެ�n���و r/������|w @����3g��7��5b�=zT �VSS��ةp ���:�����le�{AA�     �����К5k���ܻ�9 ��w�y��=b,r��[�~�z"w ="!!A�����SSS �B� ��k��䛑#G���� ���iaa!� kϞ=z衇��/}I���ԫW/     ��ɓz��Gu��"��}_��m�{ee� �;0��A�� I �(� �@��������O,,�4i��l٢��6�Mp��R�|L
 ���ТE��q�F}��t��     DU{{���y-]�T���<�oݺUs��q�v~�/X���@�JKKs��6�=%%E �Q� �������,����7��hܸqڿ� ��6����9! �~�������?�y�u�]l�    "�ĉ��O��Ǐ@��:uJ���D�B��;ٰ���3�������A� ,��[__�&��fРA:w�����o/^TRR�222 A��ܬ%K�h׮]z�GTTT$     ®��E˖-ӊ+ܭ� �=z��t�������?���� ���Ŭ��UTT�G�Ǐw���o���.r��S ��������c�;     ��;�>�ӧO@��G�;��f1u�~�?X� ��� h������sZ|����I�&i������ �UUU������@��g#��n�C���o��7    ���W��Sہ r���F�cƌq����@��ի��������4��"�; �����Syy�|����#F��ѣ�7��E�,r �Ç����>����     ���ݫE������oݺU�g�&r� o�����+���;v�&O���'r�Faa����?0���bg xv��})ihh��F��.�p��Z[[�����hoo�s�=�={�������.     ��� �|�I����ܚ
D�[o��~�G��/\�0�����v�!�����0@��5=}�� \	w @(ؤ���F/�m�-DlٲEmmm෦�&���+##C &'O��w���}�ݺ�{XH    �Mn����O� G�=a��'L���G�\����^�	kf���j� B!11QYYY����������ľ}������u�N Ll��3�<�M�6��_���N�*     |eA��?���R�!r���F�'N����?��N�\�����yĞ���$��"p �Fvv���lᖏ�����b�����?[$��� l������@7�t�|�Aw     ���Z׬Y�%K����N �^D��������"w��YH=h� �6��Z ��: �а,��.\� _�;�M����:::TYY�"w����͛�g������;x�    ��ɓ'��c��СC�C�=a��/7n�!r�LQQ����d���ƫ  T�j#�����,���[S�L�֭[��4�O����"i^^�  ��x�b�_�^?��F�)     z���/_�\����ݺ |"��	z�n���q��?g�܁K���999�콙�� ��;  t,D=s�|e'T���z ��hjjrg�w �������w��O�Ӻ�����,     z;��������+A�=A�ܯ6n�ް�|0�n��Ꮼ�,7 ��;  t,�JOOWCC�|5d�UVV���L �g��-����
 ��n��iy7n�W��U�x�    ��TTT�[�JKK W��=z��_k��޿�!r����b��?X�n�; \^� �dS����)_�"�-���' ���kRR# "����G�>}���o�V    ����U�V闿��.^�( �VD���Ƚ�������;�'999�����1�kE� %;�����b����'Oֶmۼ�������y�e@T�޽[_���t��ꮻ���    p�<��{�� �J�ueΜ9�ի�~�G�ӦM��ѣ���K���'�����='�kE� -�����$_٩�Q�F����࿶�6UUU)??_ MMMZ�d��l�⦹�g     �T}}��-[�&�wtt ��{���wW�C���������`x�xu ��}`���������Ç���B.\ �577��3����(9~������^���'��(--M     |�qÆ��/~�j�o]��mϳf�"���"���c��u���.��?�����v ]�� j���.D�ɣ���5[|����🽮$%%�S ��g�ʕڶm�|�A͞=[     |�S�N�g?��^�u@O:q��I��D�ӧO�u�]�c�}D�*۫-**� ]�� z���*++sSb|�����'j���^�}����*�� ��y�_��_5~�x}�k_Ӑ!C    @LKK��{�9=��jmm ăE��Ϝ9��="���t�C�(��=1���'ֽp�/��ī<  �,>���Tmm�|VXX�aÆ�����?;��� Qd�y�}�������%    �ry���U^^. ��ؾ�{t�+r�1c�F��x!rG����1)�C�����D� ��r��Р��v��N�[0[YY) �kkks��vS D�}�z���~�z�{ｺ�;8�    d7�.^��� �"�����=�q{�;������v�%55ս�@W"p D�EVvZ��-�M�<Y[�lqW��_ss��!"++K euuu.dذa�������*^    @�kjjҊ+��Ϫ��U �#"����ݗ�=��aW\\�޽{~az;��@� ����^Y��3[l��}׮]��� ���׻iiii��;v옾���j����җ��5�    R�~m���|�Iw�! ���=zb��ڵkUSSӥm�3d��.��#�����s�Pzz����# �j� �H���י3g��

�b�b ��F���� ��>k�_�^;w��}�ݧO~�LT   �9z���x�	:tH $�[�|�7�G�E��zk�F�>��1D�6VTT$��^9t ��� "�N��&��ή����.\�  ������R���JHH @jhh��ŋ����N_��W�-5    ��I�K�.՚5k���! �؀)"�����=q{�;�dȐ!��Pff&� tw @������F����g�8b�[�lQss� ��^W,r��"X�?9}�����IӧO�C=�    ��ֽV�Z��v[_��#r�������ʬY�4l�0�;���^�����з��l@w!p D���Ƚ��B�KNNv�Nw���C�_KK�jkk�2 `�����׾��~�����>�T    �����'�ЩS� aB�=��1n�!rG��> A���~8S�t'w @$�5Iuuu.D���F�+�b�l �����[��� �sv3Ͳe˴i�&=����6m�     �y�w�x�b�ٳG V����3g
�p5�{���"w������=d�	S�t7w @d��婼�\A0j�(UWW��(����>}� �Y(�����nc�+_��JJJ    ����&�X�B�>��Z[[ aG�=W�[�~�7j�С
:"wMAA��rss��@�#p D�-\����I˾�/��e�7���:;;UUU�^�*  ή��Gt��7�_��[    �<[�ڰa��|�I�� QB�=���)n�!rGP$''k����l�[FF� ��� "ͦ�_�xQ�}��<y�v���6 �����m���s� .�>��_�^۷o��w߭�|�3܀    =��7��O<�#G� ��"w[˿��h�T䞐��9s�h���
"w��^���1O1�@O!p D�}!���Qee���"ّ#G�� HKK�jkk���- ����ç�zJ���o���^��v��H    t�s��闿�����` ��=�~�G�E�&9w�\+���᳾}�*==]�Ojj�{ @O p D^VV����]�#F�p�ϟ?/ ���Р��$���	 ��***�h�"�^�Z_��5~�x    �N]]��/_�_|Q��� �	�{��7r��Ȱ��1D�����c�����'� �?NF///Ą��`����n�)�`������ӧ�  �Ǯ��������tW�    �^[[�~��hٲen( \ۛ���p�oTX�n7AO�6M���.\��8PQak�:x�x�����������u�I�  ���ɁZ��/S�L����݂ �����J�Eq ��ۿ�y�7E�PNN�     ��֑�mۦ'�|RgϞ \.�m������~�z]�pAQ��o��D��a���5C���Ç���. ��p�6��� {3 z�;  �ˮRjll�w��0f����6m���� �2�m�������[w�y����    �4;4la���� Wj���1b��׷�r�;2v��^��#�l �
������m� Гx� �%$$��=H�rC�Quu�N�>- �����9� W���^K�,�o~���_���ϟϡ!    � o����.]�
�՘1c�F����܁���W^yE/^Ov������ɞ���,@O#p �=�T�ESMMM
�q�Ʃ���= ��aS���� �:�ϟ׏�c�Z�J_��W��6     ���B��կ�f�w�  \����1D�D��v����Ƚ��O6��F@O#p �}���UVV���N����2e������& �`�R,rg� �͑#G���}Os��q�(    �"��|�r���jnn \���c�܉�l������yyy��ݠH �w  �ǂ����@MD�)Г&MҞ={ �Mee�
�A �ճ��-[�h۶m�7o���~���O    ���Z�v��.]���*�����=&ʑ{�^�4u�TAD��X<m���/;|`�{ �  | ;%����6��"�aÆ�ĉvE�E�, @��n���y�f-\�Ѕ�   ��ڿ�~����ɓ�ku�q{LT#�C���D��v����� ��������& �w  >@BB����u��9��ѣU]]�Y �����~o	0�봵�i���.t�뮻t�w*55U    ��������M��p�q{�;�;�������_�_�7w  >��D�*H_�m��)STZZ���&{��� t���F���ʕ+�ݙ    Ȏ9��v�� ]�j��"w"w���������������@<� p	vj��w�Qgg��¾N�4I;w���7u���.���a @ײ��%K�hժU���{u뭷�w��   ��8y�~�imݺ�u_ ]�Z��"w"w���F����W\\����9bz; � p	������Vuu�����믿^�ਪ�Raa!: �MlsuѢEn��<�Y�f��Z    ���ӧ��T�� �CW��1D�D�����k׮%n�W�����L�_��X+ ��+  �>�744���UA2t�P旕�	@0ttt���R� ЍN�:���Gn�_����    |r��y=��3.Jkoo t����c��ۺ��)S���>JKKӀ� 6kd ��  |[�������
�	&����-` ;Lc����� �^G�����}�3F�W��c�
    �Ɇ����z��7t@ptW���=v�2�;⍸>JHHPII	C�<����s��  \���wMV]]���N�N�6M���jii�`hjjr�S222 �~�����}�Mr���n�   ��dk�˗/�ʕ+Y�Э�;n�!r'rG|X���+���;EEEJNN�e���O�	�;  ��N�666�:���Tk�޽[���� ����B ����������͛�{��-�   @wjhhЊ+\�N����T�C�N䎞��mO�INN�����q�8 �� p���,�@��yMaa�[�<|�� GUU�


����v �)ڰa�6mڤo�Q<� �;   �.g7��Z�J�=���� �[O��1Q��{��ɓ'�	����*..��������O(e  ����&�qa`Ĉna�̙3YVVV����  z�����j۶m.t����Y�   p����\|�t�R7�  zB�����F�o��z��	&�Nuuu����)))a����y��� ��w  ��Mq��b;;;4��fL��6=���� �佡�ܹsu�=�h���   �+��ҢիWk��媨� ��x��1Q��_{�5������}׭[G�/���W�߲��8� �K�2 p��}NNN ������i�\�e�,�`�+��pJff�  �a���M��e�M�:U<���.    �[�y��]�n7�@O�%n��r�n�qǏ/�+���6���f�QZZ� ��n��� ��� ��`�m����Mzz�&M��={�@pX������� ��B�ݻwk�޽��    >�MQ]�v��{�@K|���1Q��8�~����^�}� n��TRR���o6�ў/ ��;  W)??_������T����O#F�бc� 8l3����+� �����9��    �)x饗�r�J�3 q�k�C�N�kC��)99Y�s�8 �Q�  p���}د��U��fMM�Ο?/ �`j�*낂N��'쵙�   �����7��/�ষ@����������w6܆�yyy �� p�˙mV���)h�:�ɓ'k�֭n!@0��Mrga ��������w7�    7[�y�������f@<%n�!r'rǕ!n��T\\,�/--M))) �� pl��E�gϞU�̩S�j۶m��􁨲�R��+� �?��gΜ�{�   ![~����+����U oA��c�܉�qy���;�7d�%&�#�Ξ���\��xG �����ӭA�v��I�&i�޽.����� �c���o��cƌ��w��6�   [yy�V�\����w�� �Ը=&ʑ�E��ƍp)����}�2�+ ����0D ��;  ]���755���CAԯ_?�9RG��ਮ�v�; ස�?����O�Ӻ���M@    ��ԩSnb��M����. �E�����F����w?���a,n�c���38`� ��{�Vvv�  � ��%��p���PPY�n�Ϝ9# �`Ӂ���TPP@(	 p��	���?֯�k�u�]nӖ�Z   �?~�}��ۙ�:�@x�%n�!r'rǟ�����Z���w#�g]�� ��]T  ��]���ب�/*�&L��Jjkk ���\�n7I  �����z��G��SO������N���   �?�&�g�}V{��qC �7a��c�܉��G�����"%''���)##C �  t!L���;��&�N�6M���jii�`hnnvS��� ;��l�2���Z�p�>��Ϲ�)    ⣽��Mj_�|��=* �UX��"w"��#nGP�zv^^��?���s h� �B���䨲�RA�����S�j�Ν��] 8��땔��~� �b� �\�R����4w�\�{�8p�    ��L�v�Z=���
)S���"w"��"nGP�4���b!lr;���;  ]�&(�MT*;�{����7��ਮ�vm,t Okk�۴ݸq�;px���kĈ   �=�V%;hjNmx  �n�ĉ���c��'$$h̘1B��#(lxII�z��-���SlP# �;  ݠ��@eee���TP����Z������c7H��
 @0�-:�w�v�ȼ��4i�$   �o���^z�%�[��4��8v옆���tEET#�}�����R!:����l�@�H��҄`����0�@"p ������l7M9�Ə�&X0 ��������| ����������B����]C�!&   ��8p@+V�p�`��� �.۳Y�f�n��Vedd(*���ݻ׭��7N��_��o��~��E>�?�}�����C333 AD� @7�+���Ң���S�LQii���� ���USS��  �`��=����o�]���#5�   �ZvCҞ={���O�ȑ#�����n���۔�����j��~���=:log�D���<x�yyy��"p ������@OJNNִiӴ}�v7%@0�&�-2q=  ��}�\�d��y�7���;�T�~�   ��Y�i�&7����L &uuun�;�{4X䞘��ѣG�@��p����z�`�!9)))��� �ndq�]�T[[� �E��'��{�Mq��� �p����+WjժU�5k��ǌ#    ꪪ���K/鷿����� ae��ڵk]��x-����Fb�ܣ�����E322�`�	���� #p ��ٗ[thmmU�0@#G��ѣG �����J�w�� �OGG��n��Ç��?�q-X���M   ��cǎi���Z�n]��b�rـ%�_-�%r?"��������yss��x����D��^?�� �x �������|���+�F����������M.��!{= ����ǵh�"-]�ԅ���'���%    ���ڴc����:t�  ���������f� r'r�
���N�x�H����}� ���w :w  z�M����t�E݄	����LCKK����B D�lZ�l��}�Y͝;W���g5d�   aa�y-�|饗TQQ! ������F�~�[hz�u�	�@�x<x07�L^^ ��;  =�,�i�AֻwoM�6M���jjj�`��l�)--M �hhmmu��3f���nM�>��m   ֱcǴr�Jmڴ)�� ��*++�q�F|G)D�j�{�n���=:��}��e�V����� 4� �!			*((�ٳgt6��"��۷��HMM����� �r��A���?�����O|B��~{�&�   ����Ν;�������� |����kÆ�?>�{�G�;z�EҶ����66� � �d�e322T__�����&LЫ��* ��������  �SVV�ŋk�ҥ�馛t�whȐ!   |ck�W�֪U�T[[+ ��9w���ovO��ȝ�=*���l�����@&+++R� �_t��  �	;1��Ԥ��6��ضX��ѣ���R~~>�R a���.z��5i�$��_��f̘�(   ��k����^z�Mm�u ��+//7r��w�(G��?j�(!,r_�`���[ZZt���bn ;�fC
 L� �a			*((p��a`�e��9sF ��;kjj���# @���v#�=bc���'�m   @OimmՖ-[�b�
�<yR �kg�6�ϛ7��=v���~�G�U�Mr'rGW���֊,��`-
 �	�;  q������L���)&N���/���Z ��&��u��� ���=����y͜9Ӆ��Ǐ��   t�ӧO���֮]��� �VYY�JKK5w��HEoD�D�QA䎮������"!XRSS�s aC� @�ةg�����t6�c�ԩںu���� jkk�uu\1 x���v����m�ݦ�}�c�&   p�lZ�Ν;]�~��w� ������.r�3g�{�G�;�������0�$`���� #w  ���z���r��M��6m��o��( ��d��[XX�+j ��&�-Y�DK�.�7ܠO}�S3f�   �+e��-��i�555 ��S�N���g�&r� "��!rGW<x0C�(;;��� aD� @Yn�0�����i���ڻw/�������Pee�;p�D ���)�6��#F���߮�o��}�   >���o���t2k֬H���G�E����w��3p%����!X,l�F � �8�ņ�/���MaЯ_?�=Z��`�����j���
 ��r��1-Z�H���/t�M7�;�А!C   �Ħ����ˡ� ap��	�Ϝ9��=�ܣ�n��Y'r��JKK�����֤� ��;  qf_8lrryy��bذajllt�@ ���S� �r��=��i��T�y��)55U   ���Nk߿�  ~:~����{�D9r��{�ȑB4�"�u�օf�����1t�P"� JOOg-@�� ����eff�j��رc]�t��y���Z�''' �+�ީ�An�h'Ndc   N�:�bA��@p�����DM�6MQ����"���}��D�$[�-))q�����7� �  O���	�aYd�/�S�LѶm��������*a�  \);�h���(**��f�}�  @x������Lk��z��7�O"�h��m"�.DCl���Yo#r��۷���������v�� �V  ��-*YTZ^^���@v���ںu������F�L� \�ӧOkɒ%zꩧ4c��v�m� $�   �u���Y�F�6mr�:  �f���O�:UQ�Ƚ��S;v�p���=:,`&r����Ѐ���0� 
� �HJJ�;%][[��HMMu��������. �kmmu�;W� ��}�ς��I�s����>�12D   �_EE�JKK��+����  �r��!ˍ?^QB�N�D�x���$���0�*�ؿ%�  xƢ�~d�iX�	�'j߾}MMM���w  �*v�j�ʕ�1b��~��7o�;	   ���h׮]Z�n�[�cp �ہ\�8n�8E	�;�{T�#�^�m��E�۷��� �  xƾT����-2��]qv�u�����v�Dbb"% �nq��1-Z�HO<�f̘�bw;��   �����Лo��§M�6�! ��ؿ��I�~����`�&D�;���gff
������%@�� ���deee���FabS:mc�ԩS����Ѝ��  t�ZZZ�EEE���[�Tw{�  @���:�6n��� ��,r���6�(J��o߾��k"�� r�6��� ����޽{ ��J  O���-�	��cǪ��Ql��`��*++UXX�D] @�;}���|�I����F��ٳgk���n�   ]����0������  f���n-xԨQ�"w"�������6l�@�!vxiȐ!����G1y@� �1J����SX��YS�Nնm�TWW' ��Ϊ�*���	 ��`�,��ǒ%K4}�t��6m�4�  �+��ڪ]�v�poϞ=joo  ��/,�9r���ȝ�=*���G�!�zn����L��q�)���  �Y�������0�/�3f�p��M�࿦�&w(��  ��f!�}n�GZZ�fΜ�9s���O  �Ҏ;�B�M�6���F  \��{�����=Z�w�Y�~�M7i���D�!WTT��UL�7k�M E�  x.;;�E���IJJ���i��&@0X�no�� �xhllt����5���sӦJJJ  �?9}���l٢�7�w�  W*=��ءC�*J��G�������������ಃf6 ��� � �/�eee���P��i�)S�h���n����F���B�1 ĝm0/_��=즺��s���  E�Νsa�֭[u��A p�l��Y����Q����6D�������v!<RSSU\\,W~~>���4�  �B���\UTT(l,�?~�^{�5�-pWVV��7,�  |q��)-[�LO?��F��ٳg��ov�!  ��w���СC�  t�X�l{UEEE������&���`ۛD4X�n7%���M�6l{y���� e�  �M;ojjRCC���N�766�رc�?������]k �O��#�Vj�%K�hڴi.t�����  ;x�e��8|���� �;oo޼���R������a>�Qlx q{���G�����dlz; D�;  b1�E�a\T������ӧO��������� �G���n�=l3g�ĉ�;w�fΜ��  8�|���.j߷o���  =�"w_����v�)%jƎ�ɓ'�D����SVV�\v�Ȧ�@��  �%�N�;wNa4a��Fq�"�\�kiSSS ��lcڂ0{$%%iҤI��  �{���ڵkQ; �����ݖֿ�Q��vۧ����=�l0UX_���n"e� ��;  cNFF���
�.m�ԩn�fmm� ����څ�� 6ٝ�  ����A;w�t�૯����6 �{oڸq��ϟ������֭SEE���n�?~� C�Lv�eII��sG0�sg D� @ ���I�a��Hvڴiڶm����o������TAA� @�|P�>g��p��P)  @O�A�y$��g  |f�S6l�-�ܢ�}�*�ۉ���܃���C�2�*ಲ��A �� @ YDj1�ٳg]\6����>}����Ɣ*�{�{ZUU�D @��7v��ۣG���ٳ�F^NN�   �҅�g�7��I� � �E�,p{VAF�N܎f��M7ݤ͛7�{�����)�'� �� ��JIIq'xkjjF���&��ڵK���f��ֺ�]  ��><x�=�������6�rss  p5���]оu�V:t(��+  �b��-_�pa`�D9n���ƍ'�RD��9;d�������s�� B� @�Y\������0�/�&L�����v�zRR��� ��x�nS�fΜ�3f�_�~  �0��;v�p� ��F����_����������R�yƦ�	�����~ � �  ���>s�Lhl��m� �UWW�+�,t  l�3������W���]�>g�7�=!!A   �,�{�7ܭ�[�lQUU�  ���[o�U999
�(��S�N���_/�J<ح����w��*))a�w�ٚr��@O!p  �,"�I�a^�6l�[h<q� �ͮW���Taa!�  �l
�ʕ+�#++KӦMs���)S�� @���չp�o߾]/^  Qc�8���ܳ���3�{� �ֲ���.�>p5���aQ������B�Y�a�  ��;  !������&544(�l��M 9}�� �����M����  QQ[[�&�٣O�>�8q�n����M
  .gϞՎ;��&��   �W��n{W>"n'nǵ��}���ںu+���h��n���(��~	 > p  $��*[8��4�&L��ϟ?/ ~��՚��'�  ��`��ݻ����ȑ#]�>}�tw;  �w�|�M�ٳ�=�i ������$��������ﭺ�ZQck�]w���0d����=>rrrԯ_?!�l
AA�  �� ���k���M�
+��7e�wճM��7�U"))Iiii  �:;;u���xꩧTXX��S�jƌ�<y�{�  ~��ۯ���v�������	  |4[^�v�W�;q;q;��{|����)�>��0 \�;  !����"s�����_n۶�-��� �8�  d��^��=��഍f�����  ��nF�)�{��u��n��  ���=�u����ns��)�q��5j���@�޳l���i?l}���l ��  �Lnn�[�kiiQX�>��,r��N ,���t7L�� ���x�� ���߿�&M��6�=�   Q`����{7�����  ]�n?Y�fM\#w�v�vt/"��a7����(99Y6{.mЉ� \�;  !c_�
UVV�	S���.r߱c����_�;ZUU�b  �������v�s̘1��Ç�} �.`эMf��ǏS� �>��]�V��zk�G�Q��m�`�̙n-�	D��o���&w_ff& �2� BIII���SEE��,''GS�Lў={؈<g�-���r�  ���;�����nj;v���f=m#  \;t�ꫯ���~644  �[^�n�.\������$n'nGϲ���k�n"��e{�����/11�=� ��C� @HY�r��E566*���������^ �Y@`p���  ���y�����#Fh�ԩ���]7޻wo �?�������ؾ}�t��I ����<�w��Z�v�v�GII��i��N�5��؄|��vmk� ��C� @�����f���+̊����ڪC�	��jjj�t�>}�  \��u����կ~�ߍ=�Mv��l&: ��־���?�{��o��֊  �_��E�,��=�q��Y�4l�0�d��}>߱c��5��C�%�	Ph  ��� ��/�:{�����ZZZt��q�-f�&��61i ��a����o���4h���h	�gnn�  f>��_]pC� ���JmܸQ��r���+���k׺A+QB���n r�z�{m���}�z�퉲F W�� ���S�YYY���U���J���~�m���-�@  ��;���W�v�����4i�ƌ�w;h @���%'N�p��-f߷o�  �����ڰa��ϟ�e�{���o��My|B�~ml�EFF��'�$~ �r�  D@^^�����#�lBe[[�Μ9# ���(�ѐ��#  н���]�N� {���PbS����  ��ܹs.r�Iז����OD�W����pHOOWZZ�  W�� ���/�eeen�U��b��:v-���_6mϦ���  �9�  ł�������B   �,rߴi�n��f������Q��m�9s4x�`>#r�2v;{qq��Zm  W�� ����v��]�v�Eq�ԩn�$j�@���ֺȽO�>  ������2�݌4n�8�3++K  t���v?~\�r�7�xCUUU  �c7�nܸ�"�(��s��%�E`X�nq�Ν;��/���쟕��#,n��\  w  "Ŧ$_�xQ���
;�g̘�m۶���A �d����;���L�F�H �@=(�s�VkWcomݵu?��;�����U�UVI�U�eH�{	ι&g!`��d�����7�+�~�s>�����s�)x `������������������]��s�=Wu|�'���F�=ڿ��*� 	����Uh{��N�v�v:ˎ;�[!��entt�
��ҍŊ��p���.቉�r�ƍ�����W_-�|�I��ӭ[�����ի�< �}����?V��������ʕ+���Ν;˿���W�i, �+�x	�7��V�~  s���*�������!��|��}�v�0��{�ps�͛7Cw��_��� �F� j&Sk׮-Ǐ�����~�嗫�{B�Щ��L1bxx�  �����eϞ=��������{np ���͛���/_�u9p�@u��
 �'u�ȑ�������'ܞ��.]*u��㭷ުB��Ʉ�)�hiE�H����07�I��2�,U�U�W^�J���
О�]�V�?-_��  �#��o���:�������]ޟ��*��n�F,t�\�}���uh���,  �!�zzz�믿����u���H�v�v�����ҵ�T��t��*� ��	�@M��ׯWE�:HW����we�޽FbCK�t4�� й�����ܟ{������244T ho����U�����
����O��
 ,��$���k������p��˗K�$ܞ��6m*�Mr�u�����RW���e�֭���C��c�?��p������ǫ��u�f͚��_��|��g
������5� @wH@��/����F���s���VSX�zw�ر��?T��F��ƍ ��rN���5ܞf0	�oܸ�@7ʚP�CҠ�nR۶m[�:�{dm�K���S jlѢEU���ɓ�	|oذ�Z(��?�Q���)�Ν�ޟt� ���`��x0���;@s� � �(��:���~��U7�Y��Ǯ]�ʑ#GʩS�J]��=::Z���
�#,�c�/w ��e˖UZ.\(u�y��k��
О�H�mժU ��w���M�G��/̞crr�  ��\n߾������e||��A���W�^-~�ay饗�����/���n�Le,t�lZH�. 旀; P�ʺ~�zu�Evŧ���d@{�{ҕ+Wʊ+
 P_Ӆ�S�Nؽ|O��9@�6�'�~�Сj�#G����(  �$��w�y�jԔ��w߭E�=�������e�;��<�����?����C�d��o�)u222R֮][�.��Z�dI`~	� ��(�FT�ų�>[�<X��t�ҥjA(c�  N�8Q�����u����3�T�[�l�:b����nt���r�ȑ*�~������봶 t�L������*�ސI^�rn�n�l�r�nu��9��O?]�.�a���� @%�f	�g��۷K]<��s�"Y��@{J�ּ?�}
 �a��O>����nߴiSzo)$�6��:��k����ǫ�����n���ŋ ��LnoH�=?� t�M��{����ޫ&��KȽ{}����o�-u���[5d��]�x��	@sH�  w���U���V }��E����s�֭r�ܹ�f� �I�A�����_uwO�}���U�����2<<\ J޳N�>}_��ѕ�N� ��J���w�y�Dϕ+W����-!������?�u�֕�I�=����!��S�p{0l۶M#�.�ϤL��9|r ��EX�_�^�"��_����"Y:��'��trO� `��9��|�����R#���7o~d��I��&'\?v�X�������:!w �:��������B�	F&�_����7�w�:��S���R��]2i$�hw ��%9���TT���o�۲gϞr�����l��|�r(  �p�̙�طo�}�_�bE��=G��9�~���X�hQ�N�:	�7:�7��駟� ; ��R�J������n��9�~�ҥ����r�l�H��'�����ٰaC*t�d�1��p ~!cҲ�x���Z�������^*����ŋ�~pϢ�"  �JB�_}�Uuܫq����xw��7nTMҍ=�F�=����  ��v��*ܞu�'�����{err�t�������;S������eݺu��ϟ�|n�d��i%<���.\(u�x����+�T!�i�����,���
 ��ҁ�h�������t}߸qcټysu��M�6UǓt%^�4i� ��cǪ�9�����  �3�p{ý��;%�^�p{L屚�fP!��R�p{-t��( �' <Tv�g�c�:�%l�ꫯV.W�^-@{�u�V9w�\���hѢ Ў����o���%�~o��22�8_' ���W���f�ӧOW�9WǩS���  ��|��V�Z�1!���o�5`��5�� ��n��_�ZM����ηm�V�z�Bw�cZ��o��"� <R��P�bo�,]�����kU��IG$͗�trO� ��$�����W�tx��>���s�O�`OP=��s��Fx=�vv �֙�p{C'���`)��G���r��(�ɴ�:��Ә)�vk7�)�5[��p �����Y��*�f1�N2^�r�[{�ׯ_/�/_. ���?�:����i>�C�ٜ�"[���!�n��K�.���bo�  �cÆ���.��\%�C����]v��]nܸQ�I��	�ױi�|��r������L�����=::Z����'�5I��p +k	H�[r�����W_}�
�OLL��$��BH^�  u����7�5+V��xo	ƧS`���̜M�Ю�y����ٳg�����Kgv�� :C3�������|�6!�LN�=�du����ۛUcro/	���/)�.u�iӦ��N���|� �Z� ��W�Ou,/_��
���ok۱�Pg�|�q��,�  t�+W�TǑ#G�knϵ^B������n�	�g�3̇���Q5Ǚ3g��7��y��6�	 ��mܸ�
��b�m6�6:�' ��r-��;��7��{{�{�=���Н�F�	�z�y�˅�������T���k��ء�d�4�,.Z��  03���yT��Ɇ��sm��ln|}o��{.�y�g�-����"a��W�V_7��M��\�Np=��  �G+��Y/N�|!C����l:���ºu�V����ɾ��͛7�S�Hg���p f,�Y<y�d-��Y�x�W��������/�,���(  �/}s��c�nO0G��_7:§@�0|�����w����c�#ڮ_�^N>�m~��'���s\�v�n��K�.U�6�9� �'�iӦ��[o�4������������w�}���[7���
�7�/���?��r���RGY�-O=�T��dm+M X� �ɂ\�$��M�O���O?r�6���l� `��}���ꘋ�ܗ.]z7 ���P|#$�.�)(�Ǒ��5��%s4B���������͸��Y��y��:���I�&O�<��|?����ސz���3���9  h���7�]���!����ӹ=Ӟ��{k�=ܞ5�m۶-�{͕�Z_��#� <�����H�(��MFI��w�+{��n����Ot �;��3G�7Z眲�E��m� �[mٲ�����&Ӆ�ʐ{�#�y��������c�8��<u��m�֭����Н� ��D��!� �J��?^�b|��/��Rٻw��;��.T�7�8 `6�� �'�N���V��nO��4���ӧOW�m&K���;v��-��$u��3�<#����� ��XX� ��dQ2��ccc���ۥ�֬YS~�ߔ�����>�v��c:��5�N    �n׎���Ե���?�?�p�C�	�&�>00P����B�͑p�����r�رRW�6m�&~ӽ��̩~ ̌�; 0k����,\����뫐�g�}&�mdjj��?^w    �i�p{úu��[o�Ut�+�^�p��S�������p{��N�,C��&r ����9ɢ������˗K]mذ�
����B��F�z�b�"]�    ����7n����p{������G}��G���u��3����ŋ���p�=� s�jժ211Q&''K]e1�������D�^�     4�����k���Q뱍������*�;���nor���F�!䧟~*u�lٲ�u��B��gؚ5k��Y �C� ��\�e���ج�A:���;,��%؞�;     �Չ������~��Y��n������bŊR7'O�,~�aǄ���g'�s^#��U�zo۶�����W�K�.- �w `^��>�A��P�pwB�Y��?�Y�ܡ��Q!%z{{     ͵cǎ�ꫯ�N��9��{B���.��y�ܟL�?���ĉ�����p��swKmqxx� �^��y���W�l�p�B��͛7W��/��B�Z$O+W��=    ��!���$!�����s{��?~������p{������	����V�^y�׬YS h?� ����扉�2>>^��駟�n�ܡ���&�=�PH    hw;w����d&!w����7�?Z�t�O��:������/��,YR h?� ���B���X�,r͖�;4���`-��    ,�g�}����+�%���[oUA�C�u�Ϥ�}�r��p�yN�]���ݖ-[V�hO� ������xed]݃�	��>H��?�-�:*,]��     �|�v�*/��R�f�6m*�����G}TnݺU}/�Ǆ�3M�n�5�� �~?��;�����͛�-�F�{��&� 4EB��V�*gϞ-u��3�T�B�0?2&0�/�L    @�=��s�w��]��4/J���?�&��5���O?M�;���!�~G�4������z���Rk\�Xt��y� �&�'&&ʕ+WJ�%�N(�쥈0<<la    ���L]���.###eٲe�n�=z_�n���|P�}��*�Z7��'�~�ԩRg���e���Ugo����˫L ��z]�  -���,�$�^w��B�0;k�	    ��2�6����ߖ�شiS��#G�T���no���,��^�:�7:��=ܞM<;v�(:zw�L���F�N�S h�tY^�vm9~�x׏0���ܳ���/�,�o�.���}d�ʕ��    �.���*���_��Н~������v���4�ڽ{wmB�	��s��3gJ��v�m۶�t��BwK�q͚5U���'� 4].r?q�Pw�3�2��v���GK�$]t�   �����W��� ����gU�x��ݥ����F���w߭&Uw+��;�~�e˖�|��B�˴h� :�� ����ٳg�<���խ�;<\������   @�(�ׯ��$�6�`����@g��?�Q�
�w���%�����wm�]��g�6m�jQt���^�5@�p Z&����r�ʕ�{��ۉ�;�oŊU   �s<h����ůIw̫W� :��{�8|�p��_�*���n����q�J�KM>�un�� @Ke(B	�S��͛��ԟ���;�;L+W�4pvW  ܭIDAT   :@�	��ظqc^��kזC� :_B�Y�}�
�I��Ѻ-�.���Ԣ6l�P��L�_�dI��� -��=66V���
�*���;u�x��j�)�   @��M��A�֭p�"�m��{���q��jS��-!���w��]Ξ=[�.S��l�R��L��u �Gr h��WS;y�E��_
�	���g�ji�ҥU��L4    �C___�q}���U�˄��*� t!����?����ojR3��!�L�N�v��;�۶m��t����2�� �J� X˖-�¬�Ν+���'�Nݤ8>88X   ��Ռ@�������g||� �=��;���_�����E=�N���lɒ%U�=�g�_c����s	� &�֌ûr�J�s���~�t�<ׇ����6   �z����uz+����� �EȽ�	��M��ܯ_�^�{/\�P�.�w��Qz{{��,B��й���ş��spG
�/��Rٷo_�u�V�n�n	�V���e    ��P��	�t���/^\v��Uh/���SB���?Kåtnv��ldX�k 揀; ���������X���*ܑ��rw��m���p{�e    ͓Ϻu�0{֛r=��o�{�ݻ��ro�}�]ng~�{�]��g�E�������B=�1��On�l� ��K'�\d�<yR׈{�>y�Wʞ={�͛7t����244dQ	   ��]�Z�reY�ti���( t��ܳ�o��o����ߖO?��0��5�.�~�M�6��]3&Htw �-����ͳg�~����W_��P�*���p   �GB�	��^��lܸ�m��ɿ�رc��>!�p���Uӂi���v��]�y睶���oÆ�9'��:�n� �C� h�؜��,�/_.�,]r��H!w:QOOOՙ����    ��I�	��_����J�yw�{�<�쳅��ꫯ����͕�fB��侐�f	����{��ŋ�r����H=r���) 0w� @[��OB�Y��g�|��o����oF7�Qj��zѢE   x2ڳ�<!�n�nݺ@=dJm���p{k%���rn�_ꪛ7o.�G��ҭ?!w ���; �V�ccc��͛���X�����kU'w ��E�n)�  @�us��A����k���[�����>+��B����ǫ�W����S�n�ZԦ�epp�,[�� �]������Q����۷?ˢL����k�
��ۗ/_^   ���7О��|]�)h�6] P	�'t�s��Bs�/�V��nO��K�.Jp޶m�p{�,]���<@�p �RoooU�:u�T�~}}}w;�_�z�@;Iq:�HYL   �W�@�t֭['�P3	��o������_��?����ZrO#���/_�\�rޱcG�H��hl��;	� m�����.�������;�bɒ%�b��C   ��hO�=����hP� �%�{S�!��#��^r߽{wroFg���n�#��y?I��z� ��wx ��%�~��!�id��믿^ur���B˦��^�}  �������]�m���s�ݼy� P��{֓�m�V�����/�(���������3�.�~��k'�n�p���˗ ���; ����:!�t;�~Y�I�=#=u�g��+V ��ֶl�RN�:U6d@=	��M��g���ɓ�zI���O>��r�=���6�!w���e����h5�z���� �n� @�K�+�����255U�_����ke�޽�̙3Z%��,��@m޼��ܹ�:b||�
��>}��=�|U� �K��3�lÆ��$���;@=	�ύp{g����p����4a�^��g���� �O� �醕���~)�ԗ_~�|��g�ĉ�-+�A��Z�n�}?���:��L ���F�=�6k@�ho�ܧ �W#䞠�֭[3��矗/�����rO�����+W�\)ܱq���<��I}2uJ ���; �1�-[V]��={��K)������5�?^�Y�ˢ�� �U
(�+���$�#n޼YΝ;W��|��̈́����`�=�x���}���֭[�zJ����k������с
�e�!w��_jl<�~�/_^
 �`E �(�`M�ҥK�_J��7��M���-�.0���p@ݥ�������k�R��x�b��=G�)X �uo�=��	[g]���yR�Zd  �%�>3{��-_�u�3=i�=���z����^��nC	�%�###��p :N
^�y�ڵ������@{����!!�,�f� ��|t��gk�t9v��Y}����w���� < 0�׷�0{�1�oݺu� ����ztt�p?���0Ӑ{�}�ש��,5�͛7�'���O ԇ�; Б�;�ĉerr�0��{�*�Z�d��Ԍd�;�j�Ƥ�m۶U?/�Ν���ccc����U� �9��ΐ���� !�������O�n�.�������Py�g�x�"�!���K� �EB �Hٝ��W�>SSS��m߾�
%�@(�l�c{:��  w46~�B___ٴiSu��7�)7nܨ:�6:��ֹ0 �/�����j�h����!���� ���+ �֭[壏>*����)���ٳgO��o
��a!w��_Z�bEٺu�p{Me�4�x ԏ�; б.J���ɓ�_��e˖���?��O�O$�� �~�$�P��,YRu��)�_�p�n�=�?M8�nڻC��'ؕ�5 B�w|����o�-t���w��]�y��\(����{�������մC��zJ�;� ԓ�; ���]zdd��d��m޼�
D�߿�Z�Gi�o�� �_�s�"A�t�ϱk׮j3�ŋ��{�l�z�j�n300p7�.��=r�%���R�����[o�UM7��\����/��}��]�~�
����Ն����sw�U'�L��^�fw��p :^�L߸q�
��p�֭+���Jٻwo�y�f��d2BBr� ~���J�gxx�:v��Y}/E�tx?q�Du��Nto�=�6dw��g}��� �555U���?U!�4�={���HB�y��lbM�]������\�Ԝ�  �+��tB�:T>Z�ݧDF'''�+��y-�, �K��촑��t�e˖�LϞ=[����=��L���4��֗����B�k獄 ,�\����.o��v�wrO��O>��<x�@]%Ԟp{�SSO	��� �&� t�����]p�Ѳ���s�}�/_^uB  .盝�5*š���l=w���.�	���@�	�9O�ڄ�3 L'!�t��搻p;����Sv��Q5e���ȵ! tvE �O=�T5�������JnŊ�7ިB�/_.�W^7) ��uca%��tK���/T��.�������D��488X��4�L����	�d�+WL�h�F'���z��B�	����-�*PW������+uˬ��< ���������ƪ�@.]���}Ϟ=�������eժUF<��<�ۥ����v���	�'��{\ �$ҡ=!�7n����t����oK�����'5�d�`�W���W��� �/�>�裪���J7n�;��[��V��L"O B� �:���U�)!�GK���W_��p�����NR�M� x��ҝ��J̱s�������w;���ܹs �	�& ��Y&��L�ۆ���ph��7o�?��O]rO�/�K9|�p��ʺ���h5���ud�N@��; Е�����.-E��^z�|���U�{�_���C `fV�\Ym�N�i˖-������ٳw���9s�@}�3_�f��u� �hϦ�<�jX��A�ui"��u!�������A:�p;����OW�����y8 �K� �ZY��+W
���o~󛪣��#G
�)���S, �LBKL/���]�r�����ɓ'ˍ7
 ���@{��a��ժ�{#H��Ξ�g3�.kj���s Z'ן��;2�MQ�����iӦ222R���/��t&K�w ���(555U�����Ń_|�
?��ׅ�E!�g`�֭[W���kl
H�>��xO��tz���( t�{�	�H3���?4�Ϟ�@�t��	��^'��s���G��G����7j*AU�\�ti�	� ]/�ׄh&''��}��*��W_U�1�|	�gqH� ���S2;	���i�]�vU�KWք�s$�~���@�X�lY��+�	��=Ze>CN�����H�<4C�����z�rn�;rΧ�i�688X `:� @�K�&�$cccU7wott�����CȽ�eahhh�i�[ ��|�&�����m۶U?�z�j9y�d��O�, �v�I��/_^�<�t~��8��f���7�	.�z�r�gğ���r�رu�k�M�6ꭱ F� ��\ �P������da)E�}��U�t�t<X�bE �F7��K�-4�� ��`X��v���L�ٜ��q;<��,"��3g
 �r����v����p��Ȉp;�&�lt�Q xw �6z{{��S�N	��P��o��F���O�����!�A	�%�  �]V4_��h�v:M��>������U?׮��pXX	���mr�t�>�H���˹��O?] υ���Q��ZI,��s��f&c�_��*�>��дV�[XOOO �G�S4��;��i�z_�~}h�ZH:�A�h�5�y.'�><<\�Y��( ,�F'�w�y�:'Z�˟���j�0�Y��y��%T�S��p jgpp�ZP�t�Raf����N�{��-�ϟ/��}�@hq �O�-)��|�O�. �N&y%Ȟpm����ty�?���SV�XQ:I��y=޺u� ��nܸQv�޽�!�F��ĉ�,�v[�n-�F]### fB� ��t����k�
3�1q���Jٿ��Q�ƍN+�@'н�5._���`f����OӼ�*��Α�		�X;hrn�;R�-���LeʆP �	w ��r��������I���_._|�E9z�ha�e(��.]Z ��'���N�* ����T�M�v`ae���;@�X��{��~�a9y�d�:ˆ�tn7]��F�4T��p j+�))8%��Ff&�ۯ~���lٲ��w�N��e�} �<�!0w	P	����z�_~Y h�����[,�I��X�|yٶm�n�T�I� <)w ��n��oݺU��g�}��e��W_�۷oZ�����z M���_h>����^
�!S#���
 ���������܅�Ꭼ�m߾]�&*�B��] ����K�t�̂�����%>��sZ( �\�I�]�~�\�|� 07gΜ�BU�+��B�k0��S�N �K3C�9�����S{	��رC��J�� �a �a� ���lٲ�z��,��d6l�Pur߷o_�8L�d�g�ʕ�� h�l�����G6��=u�ƍXX�(��=���{��*�>_�'''�p{jLPgi����6��k���� �l� ��-_���q���I���_��ٳ�����_��n ZG��5�� �O��	���K���/�( ���!�4���%�w��;w�&gCW�`��c  �144T���ʥK�
Of``����U���7�ұ=�����ɞ}��211Q��;aC\�r)��|� �'w`�Y�����T� ���Q����s
������c��v������ 0�  H����^�Zx2	b��������ӧs�bŊ288X ��e�֯���	�'Ԝ�ܞ;w����[#��/\�P �gϞ��V��\`a$ܞ��6�����܅��F��5��z�� s%� 0�\t'�~���Y�xqy��ˁʏ?�X�����M ���	��"WF�nٲ�:"E�����.t�K���c}�֭���}�v�Y�y����sĄ��X�~��;@H�}����wޙq�=��=Yˀ:k��3	"�YW]�hQ��p �F��{ll��*ɓ����/��˗���_U��&�L�- t�ǅ�S۰aCu�͛7���	�ZnS<n�u���O�`��8qB���Ҽ��ɓ��"��	 =��s��a�s��2��tr�&�GI >�ۅ۩�t�޹s����'M��� �� 1 ��Y�NK	�'dœۺukՁ���?יs���"]bt6 ��<�H�l�J �
�f��/Vݾs$�u����,��W�f~�̿|NR_	�%p��جie����po�5k�T��:C>C���G�����L���V�� `�� <BOOOս3A��I'�,p�۷O7�������+͵{e���32G�g1>>^�x��᭹0F�5r~=�� w�?�
_e�9�/k-�x��Y�����Iz	���s~Ese]qddĦ�򨐻p;ܑp{��a44x�|p x�,�$��( ��R�{���˞={�0�KQyhh�
�@�Iמft����+[�l����[iB��zjjjV�\��L#M�#k��H�K>;s�3�@��������|�)��YA�����������p;u���L˽��3�6�0�� f 5�W��:b	�����@y�7����K�
wd�gժUբ  t�5kִ����ڦM��#�Jx+����%X4�i2�!��<�ݣhoL��1�)�	�����J��to'�t%n�v��P{�S���&� 0C�<��b:c1;Y�J'����W�ٺ�����-* Э*Գx����n��٤x��Ż���^�:���j� ͓ 3���Mzy�y9۩4�����|	������Γi��w���5���:ؾ}�p;��r�J� �F� �	de��3g/�`/��r9p�@���K]���W�'�� �v����8�����;wV�K���m�	��8�|�p ��<Y��v�Zu�I{K7�t�=~�x��jt����rg*�M' �)�SPw��s{___�{�zspp� @�� <�t�N�q����Lf/��B����_V����=�v! � ��(oW)�mٲ�:"#�'&&
͗ ���d�yҥ{�֭���5�LL��̙3��t�ƍ���M��ٳm��ۭ[�N� �H��<L�Tg#' 4��; �,�=������{�g�E�����bTs��fT_} �֮]�Q�J2N�H��H�X �K��=$О)1�̞�s���O'���H� ��$ܞ)���xP��Z�D( �M� `�ʅ{
�:O�M���_��ٳ��ڭjO�=!w ��)F���`fa\�|�Z3�166֖kG��e�͗F	�ա� �R�ھ}�p;�Ш�gr' 4��; �,eWzc�p;t��d�����7�,{��u�t��� 0����.� 4WB�W�\)+V�(4׽���ݝ9s�LMMو�����  ��r~�cǎ���_�A�w��	 � � 0Y�i��ua��t�H'��>��k��%О����� �MΓFFF
<(!�k׮ �/����/�e٬�������ի��d��ٳ6$�H���v��3	�03��;���
 ���; �e��Q��u�Va�����~W����C��N��\+W�,K�.- PG	���tN�:U h�l�߾}{an��ǫϯܟ�h�N6@��F� ڙp;����[V�^] ��� ���%K��`
��o�.�^������{�a��/����3χU�V	�Pkk֬)0�t��5����hOC�+W��n��ߋ/�Xh�l�Lh�H ��<e�ΝմexPꝩ��� �$� 0O�� W;�����g���D�߿����7[����y�l
�5Ծt�R,<���׫ϧ��$�~�ܹRgΜ��\h��2�/���0 �NҴ)S��ۙN�9�u� �B�� 0������L)2wY0y����޽{��|�K` ���bd-�J�������I�n������ٳU�=���455U�a�_���|�֭p �JoooٱcGY�ti��\��� ��; �<K�9�����.E�7�|��۷�m��t���@ �chhH�i%H@k�3���>[��ƍU�;a����`��y~���� h'	��ܹ�����m�4 I� �	�u�V�x�ba����_|Q�;V�IF7�Z����� ���k����;@�%�\77o�,�O���M�=�4�R�%�GYGʆ �����.���乑�� ��� �$����ʕ+��K��������|��7m�i-�i�8?��S �ٚ5k
LG����_�^u,��k�j�s�&�@��$���o�b%�f��VΓ�?^  ���<N�z�[�N��g�
 ��V�^]������c����8����W؅b, <��L'�J/\�P h�t�{���LIP�ѥ=�/<�ܗ��q��B�%($� ,�LLN�=Se`:	�gS��� �w �&K�+��tLc~da�7�({��i��,�$��� �/���U��A	��0�.�k׮ҩڛ+���X�~} X�k�رC��GZ�j�( mC� ���N�=������(o��fٷo_5j�2�;;�v������$���Ț��۷;n�|���>Cr�[�K���ȺRBe�l �*���Dj�9 �]H�  ���E���)�*`͟�R|���?�����O?5��J��<� ��e�
LGx`�d-"����$��>66Vh�s��UMz{{��h���u, ��L[L�]�&%� :�z���� �Ezzz�1�)��:68���]u��o��t�mŊepp�  ���;�I@1�9 N�#:-���s����͓�7]�7m�Th�4�p Z����l߾]��G��#�^�6���� ��rotr���*̟,�%���g����,�W�- ��˘�L<��={�&O��I�?�|�$9�H(�̙3���Z��{k� @�%ܞ��M��dCq�x� Ў� Z,��F'w��W`^���o߾r�ڵ9�YY�I=� 03�W���i%T	��:u�T�� C'I� ���Y�:����[&'' @3d2�mۄ�y���f=7� Ў� @B�)Цx(�>�˛o�Y���_u
��,�$��iE Xh�l�9}�t`ae�F��3z��d������:�|���(K�.-4W�D9o>v�X �o���T�X��? �+w ���a�Y	�߾}�0P��W�7�|S~��'��Y��} f��s�F�u��É':��:k'ـ�A@s5>�7o�\h�l�p �[�@%ܮ���,_����@;p X@˖-�
�) 
�ϯ,��ڵ�Z����/[ϯ�B�N 0;	�e�-<�err� ��p��K'Y�xq�Y���po�� ��ʕ+���h��I6� tw ��@uΜ9#��O?�t5�q߾}ը��dL�U�ʒ%K
 0;�,M t�ԩ@{�����Tu�Ipo�L�5@K��akU  O"uF��\fJ�.� tUG �6�.��0~�����K�����}ٻwo�x��}?���[��u ��L��������_�~}�$	`�|�ϟ/ׯ_�&�\	�y}��� 0	���<N���6<P_�  mb``�*4_�p�0�R�}�7�_|Q�;V}/�󇆆t) �y x����^ҥ��	ad݄��ƴg�y��|�L � �E�'6n�X`&�"S� �S� �����r���_tg~�K����+V�'NTw `~���t�\�R�]�V X8��zÆ�`{'~f/^������
�� !��	� �V��f"ׄ�( �D� �ͬ\��
�_�t�0�n޼Yݿ�� 0�i)�� h�L)��B/�|�@{ooo�t	�7_�y������D x�6m2M�K�=w �4�  mhժUU���˅��*��� �?
j<��ӧ ���7��	�wC��A	������T�������Wh�<��9R  f"��O?�t5�f"׆�W�. Љ� �TcqJ�}~�;w�=z�ܺu�  �+a:��N� �.�������S���
͕	,�������X� ��\�M'nf*�O9��s :��; @K�=��W�f'����ƪ�, �:�3��ׯ�K�. �&a������v���ձt��R7	gd����po�tp x�\lݺ���<gr�x�h  �˧ @�K�����]�Vx27o�,�� �hٲee``���fG���r_�|i�'NZ#�r>���  �Y�hQٶm��7���ի]G��� :@B�)����f&�������d �G�IF `�Vi����Ԙ�H��4Z���/4_Χ��� �L1ھ}{Y�|y�����+� t���������Ο?_�9RnݺU ��J7 ���;���hO�5�y�4 X�xq5�����֭[͗5?w �AK�,���}}}f*����� t���S�r�۷o�����> Z#!���Sp��ƍ��;���s�3�줃��Ȉ��po� �����;v�����E3 ���; @itr?q�D���,�ljj��vu��� ��ѣG�#pϹJ#��[P}�>}�4��ڛ���������s�l�� ��$ܞ�0S�t�u�Ԓ�[� t�E��-�
��111Q<� l||��p�#����r�jժB=$�P7�7o.����5��&ͣ�uk\�r�:V�XQh�<��� @}ec���۫�2�T�v��W �M� t�,Pd�"ݴnܸQ��ҥK�СC:�@z0�1�	�gTn�M�.PG###U���ʹD?7o�,4W>��[C� ���[�
)�Dӿu��	� t�,pe����Xm��)������ ��L]9v�XuD�i��{�˻"^����s�����&�_|��\���6S5_��t��L& �z[�r�Ͳ�J���-[V �	� t��6l�P�����T9r�H�p�B :W�_�	��Z��
�g#_�C+���ٳ妮�@�9s��^�Y��r� ��|���*}}}�$ �^��a����T�!M\��� t�F'���$J��C�)�@ʹ̩S�����U�����jC_��{ooo��������r׉���ǭq���r���200Ph�<�>\ �����ƍ<��˗W����	� t�t6�C��ҥKU�/� ��ݺu��;w�:xꩧ���`vϹO��F�w����Z�����2k!7o��lyN����; �K����<�4 �5 t;w �.��!�T�����۷ PO9�x�bu|��w����9P
�	�{������rM��_���\������\yN�ر��|6� @=��Ö-[t�fVR�yc�G ��� �H7��d;r�Hչ �A�/_��{�	���y����u���299Y ��̙3��x��i��:ܛ/h�L*���/׮]+ @w�Fͭ[�V������uPOOO�:��
 �e;�r���*�,�C�)� 3��<x��q:��]������M�6�K�v��nݺU�nذ��\�]����x5=ghh��|9o=|�p �OB�۷o7}�YI��4�X�dI��p �BY�htr�Ԑ��+W�p{�t� �իW�s�+V���.� ��:uJ��FFF�M���/���<w �>��%����W`6V�Z��@�� t�N�'p���r��� 0���;s�L�;�}ZcѢE�����X���~��g�g2 t��K�V����ld����@��p �b�rO���ѣ��ٳ `�4p4W&�c>@�e�O����8͕0��{�e]��Hpi���Ω �K���W�v��V�W�\Y ���A t�N	�߸q�<x�\�v�  ̧�rNDs�Xpǭ[���d7n,4W�;h����r��y��Y�vm9t�P :[6�mݺ������e˖�իW �+w �h��{�R�p��; �|KH��;}�t��l�po�U�VUk��/�i�����; t���nٲ��l�:'k�O=�T��p ��,�dtw
��r���cǎ�۷o �fpo�t+�S-ZcѢEe͚5������sz׮]���� йr~�y������9'�� ԙ�; @�����M'����'�>��Ka��~�z�t�R��s�Ε����:��J�C���p�Z��ͷbŊ�|��j�! �9r��`��ի�VB��Y�X� | �L:�/t���͛ը�+W� �f*˖-+4��� ��u�V5�l�ƍ���͗.\(+W�,4_BM, @gH�}tt���<��A�Fi �C� ��2�>>>^�R h���h>w�_�5��{�Z��Z�q�F���pow �===e۶m���\���� �w ��Z������ˑ#G�Nv  ��f͚B�>}� p��'O�/]׮][~��Bs�9��s���d ���m߾������t�( ��� j,o6l�B�7o�l��s���266�� �\o4W:�f## �;w�\5��x��K�k��˺N�x����Z�|y��ʕ+ hO˖-���������%� �O� ��/^|��{3B��3>\._�\  Z)���h�to7���>u�Tټys��t�n�lj�ƍ���B�eㆀ; �����*ܞ�E6J�^��  ��L �������ˡC����D h5��[#w �����ͷr��jJ]�4W֎�[#�?��C �K:moٲ�,Z���\����LH��	� Pi��S|�������ˑ#Gt� ��{k�;1 ��56͗@H�];v��\yN?����3�  �O:mg�@2s���S�]�( '� �]���'''g�猍�U�  Қ5k
͕͌gϞ- L/������݉sWי'���.��lgH���*�������񶉝�;�66�����ܼ�d�¢s�[>�*ʮLWeZ}�=����>����y��p��{yy�-���8����p��� p���lff&�M�Z:/��, �ü) �;���*�r?>>�o��&��� �<������hPV�ۏ����wzz+++177������������=:w 8_��>??o*������� ��p ���N���� ���몙 �	��#[\�q�m-�^���xu�-�'(+�i�z���ݻw 8y^v���	8SSS&|�Kp �{�J�=��ݻW�� hBW�p�iKKKAy/�<x�����[���\������ׯ_�������S  x9�  ����AZ���-��?~\�] hp����� ��mnnV�δ������[]]����j߈�2P7<<;;; �'��nϐ;����Q�  �	� �:::��/���������߯� I>���emll�� �*'^���e�����ښ�5��	w �O���^��2g&[��U��p �'e�=-�@>C���~�޽�� 4�\�\�p!(K{;����g��eh������qv�p�G���� P���T\�ržg&�LOO ��� x)���jw�܉/���jp hD���6 ^���RP�lqωs����/�ˠ�lp ��w���L�Y�˷.���p �}��W������i  4*G�X]] ^���V���G___PV����u���Qtu9j,-[?GFFb{{; ���O�4 8+��ݦL��� �O:99��?�8<x  ����3&''���>}����������lp����!w���ȟ��; �������CCCg%�'�$�	 �>w  ~���^|�����  �.����[^^ ^��{=�y3��1���p�G�޹s' �����ׯ_��	g����
��t o�� ��M\�o�v( 4���pxuKKKA=r=���ee��z�H  gkpp0�]�&�̙�p�Bu1���' �7g� ���w�^|��'qzz  �bzz:(O���mooǳg�b`` (+C%��e1��ё`Xr*���hlmm �f�����իU�J>O�/��6 �l�q ��ğ��'� @������t�i���zqq1(�D�z�R^z�|�rP^>�� �fr�hvvV��3711�23 �1w  �K�������� �f3>>���AY+++��p�G�rfsb�sPV>���Ȁ��;w x=���199p�rOrxx8 ��%� @e}}�
� @3�x�bP^� x=~��'���ӕ癮�� �z:;;�ڵk144p�FFFbtt4 ��'� @ܻw/��?��- Ь�����������ne	��#���'(+��t����  ^Nooon��(������� �w �6����?��xc �%LOOe=�<666�ח����,m��Ƚ���6;;��ϵ�; ��ll_\\��.�(�^LMM P�U @��v�>� VWW ���(`m\�e����7#�^�\d�doo/(kiiI��&p���/ �q���1??PBNȢ�. P��; @ʦ��?{�,  Z���zd��7�w�q������o��<���g:�T��� |�K�.���L@	===�>dGGG  e	� ����.>���8>> �V��I���� ���O�V�����2�$�^���FTM����r:A�W  ���3�w%����%� 5p h����g�ŝ;w ��d�%e������Z ���Z��<^�{Ny	nnn.(//n������k׮���@@	y�"�a�O ��  m���0n߾�q hI��p���Q ��2�~��������*���ٳ��|���7���  �*�{nϐ;��"ܞ� @}�y Z���v�������  �H{{=\�8;��N��o������z�3}��9 ����X,,,DGGG@	�l�C( �~�  -nccCS ���뱲� ����������AYٴ(�^���f���G___PVooo��=? hg�Λ��	(%/�cOOO  �p hq�\144~�au� �j��!�p���]���l[�9�e~~>(/�kw �U��s�111PJ>g���.p�9p h���������_5j ��<d	�� ���A pv����ƍAYy�`pp�jͧ���!�^�l���/ �MWWW,..V�NPJ�ۧ��b``  ��#� �&���㷿�m|��G��ѣ  hZY롽��e�z䴗{��e���t�NOO �E�s]�v-zzzJ�.� �K� ��d��o~�s�N|��g� �����)oyy9 8[{{{���mI��Z���������ee�/�W��� � ��W�^���΀�r�� ��; @�y�f�9�?�!�?  �J�{=4���-���e�5��g:�g���`w �A��fff��%PR~���� �� �T����w����?vww ��tww���XP�ӧO�
YZZ�����AY���188�}V������ Ъ��}~~�������  ��; @�&�w�}7>���X]] �f�m�ڻ�[^^ ��00���ϯ��:(+/mP����j-|zz �jzzzbqq1J��ljj* ��"� ��r�������㫯�
 �f���p(g?���btt4(K��;;;���3a��^����� ��l��p{W�H�����c�e5 @tttį~��jd�'�|��	 h
T�<w����]���K�.���k׮��zX��V�-�sssu���3! ��;  �%1FFF�>����  hT��599�������@9p�y�fP���`����Ӡ�|�����>�, ��e�xvvV�6����n�'� ��ɠ�{���~lnn @#�5KN������ ��l��p//��#CY�&>99	 hVYb�Ly����S}�[��&� �?���������GţG� ��d���� ��	j1>>��뇯��*(+/�!�򺻻cbb"VWW �Q�G��C���y� �1�7��Mܹs�u|zz  �B������˻t�RP�|���-w ����X,,,S���k����  ��;  ?��͛122������ p���sjj*(���j������AY���1<<;;;AY�L_�~=(/CZ�~�i @3�����L\�p!�Y�^���y� �r���ދ��?��� �<MLLT�K����'''@y��i>�e�J���|�����tuԺ�f���������"� �I� ���-g�����q<|�0  �K�x(oyy9 ����alnn���xP�ŋ��ݻAY����E�ļ���999Y]N�F���׮]������d�=/�f� h.��  ���������݋O>��j� �[JQ��;@�����k033�#[���7�hd###q��U��*��ln7	 ���;  �lqq�:�������   �455�urrkkk@}2��;�e���W{�.NYyi�ƍAyy��O? hD���K�.\�KGGG��	�@�p �d���ދ>� 666 �cccFY�`}}=�����d�='�	���A������!��� �"۳��竽�Ӌp{OOO  �K� �ז�g�����O�S|�� PZ�w(O �~ϟ?�.�OLLee���ݻAY{{{������AY]]]U���r @#���k׮))�vya8�� ���;  o$[��_�%����O>���  Jp����J P���%�\�t)�G^�p�G���h��_XX�ܡNn�ˬ.V @kp �L,..���H|�ᇱ��  %LOO�	�������ʉt���������͛7��2���?�9 �d�xff�z'A�^4��@�p ��LNN�{���~5V �,���`PV����e��䤚�FY��.�^^N%�y4�r��� ����W�^��n�nnϵP^d Z��;  g*�~����'�|�|�M  ������p~���b}}=��������Ν;AYyi./ύ��ee�0�'��� ꔡ�����P������  Z��;  g.��������eݳ} �Mq]�(�����e�;��������� u������9�8�� ��� (&�Q���Ň~��� �&4��C�;���0�[���r���Hlooe�3���o�e��?��? J�`��̌2�M>�y1X� Z��;  Ee����ދ�?�8=z  �#�]g���>}�b"�9ˋF9	Mfy��.�^^�OOO�e�����8>> (���+chh(�<�� к� (���;~��ė_~��yu�	 �*.^����� �����X[[3���8z�Ν�������؈������ONNZ�PL�3ܞ�>p���}� P���z�:d�}�v��� ��p�G�p���Z����S���%���dw J�P�+WLe���@{p �V����{�Ň~X5� ��zd���a�[�ne������hlmme����EP�� ���277����E� ڏ�;  �������W|���F� ?)�^���e儝��� ��������q&��l�p//�OOO5�� �_]]]qtt ��<��ի���p^r������� p.:::����V���裏���� �}��]����� �1d05���`R^�]��AY�ﳾ�^�(+/����d �T��ds{���yyn
 ��� p�fff��wߍ>�@c( ���ͪ 4��z���"]��S��Ғ�{Mr2��; �+�F�/_��!�E�v hO�  ��ܘʐ�'�|�~�m  �-��ph,��/���������������Gy9�  ^GOOO,..���@�y�ˑ��� �'w  B�O��������?��q||  ]]]�>kptt@�X]]����{����Z����LwrrAYSSS�::�x �FFF��ի֟4�v @� ��277WmX}�ᇱ�� @{��,!��VVV�� �#����9�ה�m�_|�EPV����֪r���s��s ��.T�\w��yn ��;  gll,�}�����P�� �W�R^6��x�X����/Va���Ӡ�|��둿;��)9�cqq1����p; ���;  ���'����q������O5�@�����;@cr�����e������\ߺu+(//n ����W�V�1p���i��]�  ^p ��ݸq��к}�v��� �>:::�k�	����Ƴ��GGGU�&e�����>>>���Π�����wG����+W�T�b8o�� ���#
 @��w�}7>��#����LLL��`}}]�	�A�%�������	�ʀ�_|��k���ϛ�^\}��q �y�l~~��^� ��y�"'
  �-'�  4���o��oq������O�C~ ��]�x1(�ɓ'@������e�:�5���AY�L��#�� �000W�^���ހF��０��& �?p ��ܸq�Sx������ �u	��#��h\."�#/����lBY9��W��UP�� ��S����	�����"� @�����������Ç hMy�Ey� �mmm-�?���AYp//�飣���rLYZ�D��9� �����*؞�*�(����a� ����s������ݻ�駟���I  �cll���lnn���A и�{7/#]�|9(�ҥK���e���j��l�ͩH�=
 �O���I5�(2ܞ����  �1�  4�7nTmT�oߎ���  ZC6�R���r ���<y"�^�l������iPV>���phO�������6�(�y�=����  �)�  4����{�����x��a  �/b)O��9d���tbb"��ւ�<��q� ���􎅅�j24��e����%� @K���_���q�޽�����j�; м4��cee% h|���qxxX�)+� �孮����Qtu9�,-/m�������688X��{{{I��s��� ^�]#  Z���b�������n  �gxx8�����r�d���w^J�������g�}���tN��|�rP֋�TSZ[N»r�J@�n ^��;  -'Go������?��� 4��Pޓ'O�摿����uH�pL�+/�i�z��������###�F� x�  �������<�?��O��k �9��#��h.&գ��;&&&buu5(�3]�K�. �ghh(�^�Z�_��tvvV�����  x�  ������۷o���f  �O��Be �e}}=Dj�A��<���K~|��y �����ʕ+�(��y��� �M� ����������O?��w� и���cxx8(k?�����qzz��˂L5Ȁ{�!P���I5Qfvv6(��%҇ �-��NhX9a9���� ��p �-ttt�/��jS��C �x���#�d 4���%�d#j�#d ���p�G�	�4��g�]p�F��f�92� �(  h+�������\� �E��� @����̙�����ՠ�'O���t�R м��x�ɩЈzzz�p{ggg  �w  �Nooo�ۿ�[ܽ{�9�� ��{=4�4������ߏ����������tN�˽���g���@��w���b���4*�v �w  �֍7brr2n߾��� ��<�:::���� �����V����悲2����)+��L��./�~��A �r�̕+W��ihy�6+::: �,	� �ֲ�����}|��'q���  �O��]^#M�h^O�<�����wfy����s-���r2??_�_@#���� �R� h{]]]����q�ҥ���ϟ? �~���Ayp�y---��^���T�.NY����� �m`` �^�����,����n Jp �����lՈr���X__ �^?��ς�%�浹���������m���y��366V&�ƒ!����H�4���AE @q�  �7�qⷿ�m|��gq���8== ��lI����:99���� ��e�z~~>(+Cf�������BPV&��ƃ�����S��gh���pLNN @i�  �:::�֭[�A�G}{{{ �555U��)+�� �-����e+eggge	��'���GN��u]�9�э��(�  j#�  ? �����?��'����� ('�$)/h~KKKAy9a&�)�?��L�'� ����?33c?��1::��� Pw  �y������q�ҥ���ϟ? ��9Э��@k��ڪ�����ee������m�tM2��������W�V�����!�  up ��0;;[m�}��G��� ���ֲ�������� �5<y�
FQV���?�3(�3]�|�M+�߅���ܞ��.�Ӊ�� ��	� �K�V�����q������O���$ �7799YMM����MM� -$[Ņ�˛������8>>�p���;@�zzzbaa!����A�۳�bpp0  ΃�C  xE7nܨZVn߾]�� �L�(/�� ���������e<���<���}- �366���պ���i��� p^� �5����{���㫯�
 ��e�$�	����p��ٳj�e]�t�{�;;;�隌��G___��� �ttt���\LLL4�|ns����7  Γ�;  �����կ~Utg����a  ��Ÿc�[YY	 Z˓'Obqq1(�e��d���kׂ�����o�2���caa!����EN�5BOOO  �7w  x���qrro��Vܿ?��� xy9�[#Ty���� Z��{=�2^WWWe�3-�^w�2�"���L\�x��wh���B��' @#�* ��tppP�(ϐ{n�����z|��w� ��<�\� �z2Ly�d999��]?���L p��������'4�llϵA�{ ��;  �����*�~zz�w����DVXZR�	��C��5�i~{�w(ee���uyO�>��e���V̽�� ��MOO����v�N___�?���  �D�  ^A�3؞!����?��ϫ��Ǐ ����!�к��3'�Q�����3-�^�\�gI �/����ݻ�f400P]�p1 hD�  𒎏��p����O���f`��eVj��6<<llwr�� �&�zLMMEWWWe---���׃��ↀ;���������h69*��  �J�  ^���~���T!�W�����z�jr�p|6� ����  �-������Q������3��� �'�sss1>>ЌFFFbbb"  ��;  �����X__�`X��_�|����_� ځ�{=2�@���ݍ�O����PPV������)x���~(+������A���暈�����hF��w9 h�  �2о��V�B�{�6�G����j @�p�GN���=y�D��ڮ�ϴ�{=���o���\fgg��.Ќ��)[ۭ� �f!�  ����
��u���ѥcccq���8<< hG��@��\��$ Z[���_����������JYٔ�ƍ�<w����5�����Ќ2ܞk�|� ���;  �����*�~||\�#}��N<|�P�; mI{{=rMsrr ���S^6�NOO��Ǐ��2�N=L& �a
�����0�ߡ�6�ι�  h&�  �7vvv��������]���m����j�����#� ������{�t��r#�^^�lmmU{&�522��ٳ ���ߍ��.L3˩¹~���	 �f#�  �W������ӧ��w�Ab��?x� 677 �A��R�F_�������sI�>�L��#��{�� ��/_��̺���g���;  ���;  m/�ӗ��������������U�����q|| Ъ�5jll,(��䤺�@{XZZ�7neMNNV�𦰕���7o�	��U��_�z5����Yooo\�x�jp hV�  �����XYY�`� �~���U�}{{; ��ۅ����ׅ� ڈ������2�=
��K9qϺ�<�	�v��|����x����ɉ�e ��	� ж������<,m$9.���뱺�Z�ks���1�� �G^�΋�###AY��888��m��ǃ�������� h7��>??_�������T  �w  �N�����5��]nB���ƃ�0> �
�z� �K����w�ҥ��L��#[ܿ��� h�n�{𳳳��i	y�d� �w  ����ϫ����a4�ls�v�Z�Xv��}m� 4�����������~�����?�yPV�e�{=�(+�o��vP��;�Nz{{���l��f�4r}�Y  Z��;  m#ǵg�=ܛ���X5*��ﾫ�� Ь����#(+�@{�00��Z&'�<|�0(+/m���j֭A�����v{��\#MOO���@  �w  ����V��C�f��p������^ݵ�Ќgꑗ� h?���շo^��,�zdK��Ɔ	@5������� hE��>77�嚖���e___  �"w  ZZ�����ƳgϢU�5���f��R����}-//���ҥKA=��]���pZQ��_�|9:;;ZA>˹�b$ �V%� @�ʖ�<����m�p��A 4�l��Ce���о��͛7��2p��歸��h���/~��Ӗ���� h===���PM��V��u��]�  Z��;  -)۳�=�[Y����|�ܵ���&''���vTi���� �S�]���ƅ�r��m�>�ʀ{���eI�2� h��~����A+���֠�k �8Q ��lll���V��
f�{��Aw�q 4�<����о�����AYٜ)�^^N�˽��,IY���1<<;;;Ь2 <??_�N�V��t^�p� h�  ��l�ZYY����hG���U���G���z h4��X^^ �[^vp/O�u}?~,�^�\���*/���� �rFFFbbb"  ډ�;  -���
se�W;��쌹��*�~��}m� 4�<\����p �o��vPV^"����$(+��[�n�e8����
�f����?���~Z�s�
 @�p �����V�姧��_e��;��}�]��� �����* FY��� ���7��Ҳ��m���MY9�/'�utte�L 4�|/dc{^������=55 Ў� hj�����ls�֚�m�x��M�����.���⛛�U�8e�G����ط��f"P2D�-�;;;��c~~>���ZM���:SY ��� hJ���Uk���^�ㆆ�����෴� p���w H��'�^����來5e=2P'�4�l���oNQ��N+�P{>�]]"] @{� ��d]�������bT���X����ٳ �:��孬� ����;AY�����kjZ��ƭ[���2�~��� h4Y播���V���_]��3 �v'� @S��ݭ��OOO�W���7oެ.�����I @i����;�������z @ʀ{~;k6-+�y����AYy�/'�uvve�L 4���?;;����*/pLMM  %� @���؈�������{6qe�\�9@i�ޡ���� /<��������ʵ��{yn����eyy95/��3���H�����Ъ�&�  ��� ��^`���g'Ǹ޸q#677���l}�r�2�� �[9�K��<����d?�zd���;p�2�~���_ZZek���`  ��� hh���UXK���< ���G����z �YB���; �(�����/����ǫK�AYyi�W��UP^����@�2�;99�/_���΀V���/^����  ��	� а�>}kkkqzz��m8ա|���� 8144�urrRM�����|Gdx��2|�����\�d	BW�#��\R�C���W{	��r-���<� ���� ��d�}cc#����z����;�S5�e�� ��l�����b� �(������
�p�G^�XYY��������>��9�/��/]�T5�C+��?���P  ��� h(���U��X��	9�utt�:���� x]���� |���,�^�5O}r2��{=2h*��6<<sssU�Z]N'���v� �%� �02H�-\r��Vm��{��qՒ �Jث����a�[�ne���G__�K�5�g�z�d�;w�@	�^�E+.��.r2���D  �r� h;;;�����Ӡ�d01�ܿ��;�] ������By��!y	*/,�.��0��~����ϟ?���|�J�Zۻ�DVh}�֞���V  ���  ���@{�3�N���ׯ_����x��Au� ?%1F.���� ����
OOOe	��#/l�ōl����J�Vs?�,�>�+W�&khy�4K��
 ��p ��Wm�Y�#5�e�ѣG����q�%HW�x��y���r2�D=�p�ǥK�܁7��ߧ����ݦ��.r�L�M� x=�  �����*��!w�K@d�N�Լ�~��� |!�zd� ~���Rܺu+(kll,���}'����>�����/�u���|���v���y����3  x=�  �ngg'��׵7�<�x뭷�Q���� �����Ey��)9�+��l��0��~��{������������j^����\w�����h9wrr2  x3�  �&�� ��ӧAkx1Zvtt�
��� Hy�m�xyϞ=���� �sttT}���R^�����=���7;;����ﳹ� /+/������"�Kr�O�7 xs�&  �E�///W�Z�����XXX����x����; @W�'O� ��|gx?��w건�$�^�l`p^Fooo���U��N��!ˀr�-  gC� ������V��Nk�w�y�
N���W6�S^�� �ed����ePV6v������^P��~���1_|�E �����-��N:;;�K�=== ��p ��l�>99	�Cf���Tm���ߏ��� ���h��<�. ^���ju�<8���o��&(kcc�*U�����g:���'��.�K;ʩy�� ��	� P\npwwwW����#������Z<~�8���������.�N����v ���p{~�g�*e	��#���Lg���2�766V]* x!7\�r����v488X큙Z  P��F  j�㹳�{yy9�?������lsϐ{6j�h}���Ay��^�U����2�N=�p�G>����ݟ��Z�iW���չ  �� P�lq�M�c����#:��gbb"������ ZW�f��t����G6�ĳgς�����zd���/���W��9��ыR�lo �,w  j����_�O[[[A{���7o���z<|�0����֒}�둗�U�T����r<TZ^���o��677c_в���k}��=ey��˗�hWY�k����  �<;�  ������S�;k?y�#<?~� h1/���ļ0 ���䤺 ���(�ҥK�5��AY��ϵ�5(���ؒ�ggg]����{0���  ��� �s�#s3pyy9������m'9�6��<0��E�a���)���0��{y�vM=��k}wh9�snn��'��<˚���.|  Pw  �U�r�Ѧr?88�O����[��Ç�FZ ����tP^�� �ud�򆇇�0���nP���RP��L��_�ڲ�&/j���@/�,�����j-  �p ��e�w�����ӧO���M�Q���㪕���4 h>��!����o��ϟGwwwPV���ݻ����{{{������t����@kʿ��R��4�,���  Ώ�;  ���yOOOlll8(kSy��ʕ+199<�t�dFFF�jprrR]�ב��*�FYy�_��9���իAY�o7>>^M�Z���P���E___@�ˋ�y�˅P ��%� @C�`\n�a{�Ӟ2y�������Çqtt 4>������w# o"������g?�!�^�|�ܡu�^|�	r�&�׳���iS  ��;  '7gffbyy��N�ʃ����x��Q���i�hpy Hy�F�7�a`��6�����Ӡ�����9����?���Dռ���y᯲��e ��!� @C���g����^о:;;����6���� �1i)�G�� �Md����a���eexP��������ݍ�����|�3k�"4��^�r%z{{�녏��)� �#� @��ò�mnnVho}}}q�����ڪ��@��J)O��7���|����e���_���	�]�������դ=��d�=��p�*v��  �G� ��766V�ʭ��j�"FGGcxx�
c�����q p��0������~ ��ZZZp���K��z��'/n�C��"��f�wR6U������!w  ��;  M![agffbyy9�?������ѣX__ Η�{=r- g!���788XM�y��iPV^ڠ����h|��>77W� �O�Ѧ��\�  h`�  4���!�l�����gbaa!&''��Ç��ٳ �|��C���������o5�������V?�P@Y���U��I�и����ʕ+~'�?�@{��X  ��;  M�Es���Vlnn���i@�ܼy�
hd����ze0ntt4(O�������^��e�>�W_}���	�9������X�����N^D�L���������  4>w  �R��2L�m�ڢH/�W��ȐFj� P�<<wp^^N*�fR 8+KKK�5�t�RP�|��_���� ��X2�{���$�{y����  ��� ���cVgff��{�U��-,�\d���ﾋ��� ��<D���� gɻ�1<<;;;AYp�p���O8###177Wx���]&''�3  4w  �Z�D�&���5������ު�->���� ���P^^���������������%����?�y����7[�MV�������*���S_�  ���;  M/Ӳ96j�p���4��ܼ~뭷�P`6� g'G;����i����s~+e�+ee���ݻAy�fd+/���%L�_���	����׼��E8  4'w  Z���hrσ5�Q��<����<�Ƀ���e! �H^2��f�upp��� g-������s�#/�߸q#(//n�C�����˾��G�t����!w  ���;  -������� ���a����|>2���ѣ���7��(/�C.gPB��)/�+�U|gg'(�3]�P�����BZ� ?,�[�� @�p ��Ѻ��O�>�G9�tqq�z>������ ^�PK=�] Jȋ����U�%ee���{y�<ommU��(+��L���8�2��<;;[܁�S\3�>44  �w  ZRnfNMMU�6O�^����[oU�>����2̒�[��w (%/R-,,ee�/�KP^>���e�D�	s�"p�����~����������_r�e� @kp ��e�Mnjf(L��'���ƪg%��P���$ �ifɐ;e���z @)���w���͛7��2�+�g'�*3���|o�O�)y�� ��#� @���˗/���j���|�������������bmmM�?�O�D��5��W ��a`����.Woooe�w}~�k=./�������������jbb"  hM�  ��l��֛������
�!���177W�6>|(x �#��Jy9� J����l��wߙ����f���ee�=��LN��788����?���e5YT300  �.w  �Jlf�&T~J6�_�~=vvv�������m�y�HyZu�C�o�^���a�;w���3-�^^��'''cyy9�W���9Q2�ہ��5��� ��� h;�ꑣ^�5�����o�]]�x��q �4������� �	��#ܩG>��=Oy9�I�^^WWW��&'H��q��䔃�T��  �>w  �R"���Ɔ�༔l)�0g�����i ��lˢ�\��\@�����wtt4�������=�݅G�8<<��G�眓��[:�����wyN:�5  �C� �����U���ښ�2?)���?ە2��ڙ�{=20 u��ىgϞUS�(+/�����,�{?���ϟW��r?$�"��!��>tg���V�+��{q1���7  h/��  h{CCCU�=[�4��2���cnn�
�?~�8677����#�C P��X������/��2(/���g��؟�e����\�W7<<\����x59�&��3� @�p ��+��̝w���/#7�3���̣G���ӧ�FFF�߁�'����ޝ��q��>⾯�)�
<�d�d.揙?v��v��'20`L��w6w��ޓ_�mE�D��T�� MRJ,�]�Uu��~p��B�=����υh���QlO�
pw���u�  Ɨ�;  �?�$[]���.�o�ۺ��_���r~~^ F������J�F �/	�{Y(���f7�>�{���>���r����,�L�}ww� �/E*Yȴ��Y<xP��I[�Ç�z  ��;  �-��������u���V��W�^�m�///�(p�� ������UY�Ko=~�X�����jp;A�qwzzZ�/ڡ7�͹=*���i2/�gNSS�L  � �;�Mmgg�N�iN�2q���Q�?	��-`�����p`r��7�z+�����{yO�c��	���?���ͮ��ON��4)Z__�@ �7� �=�֝4�e��������V�q&�3���Q����յO��|���^��r��{/^�(����˨h������mm���=��=k �m�  ����j�{ڸ����E&��@&��={fp���6J�u:�rrrR �����fgg���j]TOo�yNvVK�n����<o8>>.@�yq���\|������)�  �6w  �	�g��իW��jff�|��W5����S�@k�m��K�( BX�~eii��[ͮq����Uy��uy��Qi��@{�+X	����R������=��  ��#�  irr���2��m�m#Χȃ�����50�ah#���� JZ	��^�1|��w����m�'��׿���/_�T� ���P���K��p<xP666���r �_"�  w�-h������u�O�	�����	k�@d�����B�%� ��0�7�|S�,L����KH��Ci����_�U���3�����<�|���u�Yv; �p �O�ɍlG���+�d>K�j~����]�����yV���#��\ �AI�����������[警� ����Ǐ0	�f����ͺ	�|��4����D ��!�  �(����H m_��,ei��H��ٳg��� ��H �u ���t�nSY�Ko��J���nOIA��E��9s,�155U�����˱�}+++  �B�  >���jm]k���slll���_��ۑ_^^�aѦ@P��|�� ����]�������w�z/��]���!���"���sD�vz�a7==]=zTwE  ��p �{077Wvvvj���i�ϑV�L�%螅	:Z<Z����'��0Ȃ����7��jZ����{yO���ki��m���?�7&&&j�V�����R-s�q  �B�  �I&A2rppP���MN���J[[&��4�����M���LJ����U���- 0h����h���>�{/�����Ͷ�3��ea���f���n�9� �W�mVVV
  |wk  p�VWW���l#k��>$���V�(�~�".z/�+�� ٝ,�s�Ko�:K���r��g5	��Ev�1�c�|M�=�G���p�r\��� �� �  =�	��RK( �C���D\�V���t�&��^BW 0,��V�����ӟ�T��LЦ�{��+����ÇuAQv� ����R}n��$  p� �GҺ�I���CAd�Uv�ꫯj"��ׯ_{=�ϴLR�{	]�����������z��Q����6^k���w�}W��˹5�R��i������ό  �'w  豕����F�����%s��կj"��R ���ʄ�魛���� �^�Eڄ766��ez+�y63==]�"w �nۡ?r�g�m�\ �=� ��7*	 ���SP��=�ނ�@/|��������� ��8;;+���emm��[��p�����s���Li}}������R6�����蝥��Z��%  ��  �'yЛF��e�:-�p���{��/_�t{h�`��I���?~\����p?&&&��v{{����z��;%�/��lyy��
�;��M�}qq�  @/	� @���oB�^��mxp��P�ݟ?^>Uh=|���{?��c�a�ų����
��v��,��4�fM�yh��gZ�GE�����?��	�C�d^c�>c ^�: ` � 8��	h٦'t���K�өA��� �*A����B�	�0�r/�{�������[��ay?���ԅ�y��`�(_�������r��C�5��yF  �"�  �����j�����@/d��׿�u9==���Y�4�^!���at~~^�!�zokkK����9a�f�Ev\d����P4�C���';�e  �I�  ,�3)����ڴ��4��w!���J �/^��A��~�m�o�@��G��븇Y�w���q&����-���"  �&�  C`rr�������n��z�	����Ԡ���ax��Hp �U>������[	r'@vssS�Q�Us� wB������d�����&;`漐s�<��WVV
  ��;  �4��=�\z)a�o��F�;�^�ȴuh�`�%����	;�;���esssl������eii��~Y 155U���
��|��9i�ۡ�fff�gN�K  `�� `���q&o��Fw赦����W����" Ti���:�N9>>. 0�� ;b��Io��kT�5̞�\�������� ��?��&؞]4�C��� �{5 0� `�r&-3�����r}}]������W_�@��;	�{BJ �Av}p��GE��>|XC�	�
���]�vd�Y���j-����_Q�3��  ���;  �l����W�^�������3q������a<ip�Qmi`�$T�O��O��J�}bb���ܔ�����#_�߅����Q��/9o�(�	��3;!w  &�  0��`9�GGGewwWИ����'Oj0��˗u7�6�,�O���X��s, ��s?��]z�	���� �S��O©yv!��[yo�����@�	��`�nmm��   �H�  Zbyy�6k�����@����Ԡ{�
	Y��]�F_��{������ ��������777���{�������~�Ү��� �O�>-�F	��s$�<oczz�.Ps 0�� �E��ygg�����0�6w�)�/���NBf�E��0���#�S�� �������`X��D]__������C���i�,�Ic{޿y����R���+  �N�  Z(�iisO��m��l���|��E���.�h�B��/��� �'�[��/�R���}Vv�K;{F��ڇO��@[��Ç�� C �`��  �@�  Z*����~������L��y+�i ΰ�F���lY]]-���; m�ŭ��ibb��;	�&�֏��@{�����,<���(0��M�=�2�0x������&  ���;  �X&��춸�X��4�~��H����+ϟ?/���h���^��� h��+)z+�c��'О�_~���z��A}����_�a�`{s��{�����eee�  @�� �Ȅt��r?;;+0�0I�\&Mkн���}F��,N��r�/��{	0������4��E9��������R���6͹&τ�a8dw�\�MOO  h#w  ��<�	�E����� d"suu�������ŋ���C�{��� �&�����������Ok�]����k�<�����Za��^gXdWɼ�ͳY�   ���;  ��l7�֤��...
R�3�����0����=z��˗ �&��فdbb��;���ess�.(�%igM�=���-�j1�r���v�cP��1�BdWI`x�N�fff
  ���;  ��<��$S�Ě����ꫯ�v�	t���`8e"Ԗ�`�w �(��_����VZ�����=a�4�'О��k����?�P����&�,� �K��.  `�� ��ʃ�L:%X��ի;ok���t����I�Y�B�e��f �*�k��K��	��-����|"��釜s��D�CZ�a�4���Q �Q#�  #.�JiuK�����0Ȅ�'O�|�3���0x���E> �Vϟ?/���������h睲�z�Y`��5�>	�'ܞ�;  �w�  0�����]��a�	Ҵ�'��6�>///0M��'�@�5���T����2�]VVV���b999)p�R��P{���`8�y���zY^^.  0�� `�����6���]��cr����//^�(�N� �����s ����U�k����1�����Y0��2�����0Ĳ%�+�Y �Q�  �L��iaʤU���3l����8>>�A�����Z���� m��H\;�`	��dO��Ǐ�B`x�x�3�,B �q �  cjaa����֐��l����R����8�՛���N@�{��ϟ?/��
08	%çHPv}}����|n9N��>==]  `\� �K�{�NS����0C)8O�<���	��z��\]]�~MLL��Iv� ��k�˧�L5���q;��GGG>F��	������_�����)  0nܵ  �%{nn����
�L�nooנ���^�z����d�&�����(�������a���������9#����733S�ټ �8p  ���LȤh��ooo�4mll�0���a��̇ϗ=�N�SwN�Q�E��0X	�����o�wI���VWW��`�5��kkk�[  ƚ�;  �3��z~~^�;C/<���899)/_�,g�'p�`T�\���Ng�-�K�}��Q��  ~"�  ����}_`�VȄ��_]���k���ׯ���M>^��^�Q 0*�0����C�177W~���mrr��x���±�.Z� ��y�  �W�'8��B��0�fgg˓'Oj�]޷�e	�$C�e�	 YT�϶����&Y�-<ƨ��y}}]�}�e'�,XN�ݹ�'���  ���;  �����kX8�it��N��lkk�����䣣��[�z/��� 5m�����?�����ӧO˿�ۿ�����@[��6��f(%?	�/--�`{,��lq
  ���;  �Q2Y���P^�~]���
�A&����H�%���i���{�d� ��ŋe�tڟ={V������3��&�4��?��	�k{����  &�  |���?~��N�&$,�G�d��_��WuG�,�H����e��e� �rm����/Jw�=��1%��Yh�}k^;�Na���Ζ����M�h�쾐�����  ���;  pg�:5a�4�js�mҐ���U�	�$ srrR`\ebuqq��{	(����H�������?3��Y8�n�� �.k(>��0h��9��ӧ�Qy#�jy~���K�^y&��*�?  ���  �$�6����j�6�����Zi�K����ڞ޻���� 0�6�e�=��|�&���ٳ{�nϟ���
�@;�$�+���k�]FC
cr\km ��'�  |m�����W_�����^Nx&aT�р�˹�b0 FU������~v>��ڳ�����^�	���/�1 ��=}||\�m���ur�S,�_������  ܍;c  �isgT�����ɼ��
�PM�0�4��G�9`T�����^O�~�ߖ�@;w���T��VWWk{;�~9�sloll8� �	�  ��isO��P0m��Ӯ���tj05�5���5DA�%� �*��s���_~���nI��	��u;���������������/���,���5خ�FK�e'�<s  >��;  p��澵��͝����P�����޴���FA���^��Q�`���	��Z�; <����|������쬼x�^���lA4+��_��>!w`t��}ee����im �{ �  �6wF���t����1A�,�6����˂�� `�%��Hx}�<}��MK���u6	&��1h��g�={&�Ν$��d���+0z�ڞ�+y  ;  �3M�{�ө��h�������j������Vw�o�H��?��Q�]����]��m��K�ޥihov888(pWY(���!�
#Lk;  �;  �senn�4^3J�����N]ȑ�w��v,�-�X__/���; �������,m���,��=+������%̞�����=�"�G��p;0��\0X�|  ��  @_LLL����:ɗ6�����brr�Nhe4;dD0���.�?��c �SZ������xh��@����|FW����=�;  �#�  �U&����˲��_M 3r��#����eww�[��a��_z��ࠜ�� `8	���,�ϽY�yM������ʎ�Y<�p{B��h�1���  �{�  @ߥ�&M����E�Q������"N�5���c�:���� �[&О����:ڹ/٥0��ik_\\,���q������  �w  ``fgg���N���]�Q�l[��&���'�na��f�4��{	S ���訜�����@;���捍�z/55e��EJZr�ۥ  �˝7  0p���u� ���������=m�	�g��������p���_��ׅ�H�=�r�����l���.p߲h=ϭ�֮��KS���  @�	�  C�	�&��IjMk��L�gb<C�;���-���t�� 0��pnyF��ߞ>}*�N_4m�	�[�%�햖����z���(  �`�  C%����5�m�a�iugԠ���@;����"�� hkfffjk���l  K�  :i�z��QY\\,�_�6��X��N?���g}��\ی�����p�v8::��s�`t�s�E�/�~��4\2�5  0x�  ��ZXX���{{{��Z�5�B�;�� W���_���y�%��l�mR���@{$P��_�����ɽ�@;���h�yHZۧ��g  `��B  ����D�`�d�6k�Mw�{��9��.�A/����~�����n�ݡwm�����.L �A����@{ ���5�AH�B�3eA��oy�s�E.  0�� �V���);;;���n[���a�4�����Vw����<��������Z}&�����l��r�:>�=�r�r�����s=���3���b�=L����Ɔ�.  0�� �VYYY�i�>99)0n�[ݯ��kb��i߆^�¢�{3�����^�9�ix��ڪ�g�&-� @{�{L�3�.��I�v-�+KKK5Ԟ�� ��겋��.  0�� ��I�NM�=-�0�r,d�>#���_�~혠/�VΌ?����g� N������<=�A��� �`�7�|S�8݁������677W[�3���@4�yN��  ��'�  ����BS6˄-a\�X���ޮ�C��	�8.�,���ꈄK�E	��u&���$�  �.فE����@{����Y����ZC�	�t˳���[�  �"�  �Z�wҼ��{�w�1�qyyYw9pl0(ggg�/�K���:I�{�򞟍�W�^���� �K��D��a�{�<j��'42o�y!��VVV
  �>�7�  ������\}||\������u�q�f����ڜ}rrR���o�4��|���o����dsޣ	����f��K h�\3�rii����s��������&��	���yvv� �K>�����  @;	�  #%����5ț`�f�;;;o��+Z[佘��w�՟-//װ{����&~ ����>.����zݒvv�v�Y�06�����x����\1
�� `�	�  #'�<>����_�.��������H��	�;Ni�������Y��4��5l�h����� -���7�|SFQw��ٳg�3�rͿ��X��WWW�0�(猜+2X  #A�  Yi�I[���A	?Ip8c{{��5&�q}}]`X$���?�SSSu�Fw�}��.9����
 �N	����@{^s_�.�r�������!u1̤�0  0R� ���ƞL���+-ՙ�~.�Iv<�x��I�d���h[°Ix<!��H�=�&��� �0���q���i6ϵqۜ���k�v�&��yv�ݚ�x���sG��)o   F��;  0������V�t:5�]ޭY�qyy���=���������o�{xee�M�{��Y��/?��c �-!�6�l�@{�?r-�{]h�\�����Ūy�X9,//�E1�  M�  �Xɖ�i�I�]�vjx�,IH8#�$��L��0�r^o������r�������5����p �n	���7e�$О��r����3�vZ'A�<�I�=�����psss��=Ϭ  ��&�  ����:��	$����3������q=v������M�a���?�PGdB��Çu$��׉�����$T�� �n	��,,}��Uy���@;����<�I�}vv� �U�daLvX  ;  0������U:�N
\]]��5�@g<y��s�������H�/�K155U�6iwoZ����� �~��=::�׼��v�=;(�Ʀ��k�,���s�,�����  @{�  c/�cg�5ͻ�qҞ�m�3�I '����M����˗u|��u�<��iwO�=���:�!�� �!-���3jr����Z��WVVj0�Se�;?  ��p  (k����bm�>==-��ˎ	g\\\�pN��4eC������o�w�}W��[�������]� FG���o���3���K�yM�=��fY�k�,|N�]��\Y,������n  `|�  tIH7M��N�@ �fff�GY,�V���������Q��}�>;4�yM����q FCB蟫	�g4���3
b��PjO�s5疔�d�  0��  �aaa���M<|�G�?.'''5�qyyY�Ͳx�~�#��<f�Q���,nK��c%О��	�7-����FA��yV����Ɔ�_�^��Q�-)  O   �#����]\\�!��O��)[Kg|��5�V��F�? `��x���ic��ͧO�
�3�jOS{��)p߲X&���k   �	�  |@&p������Y�_\\��u�ݟ<yR�4�'$  � �����7o�hg\��������eff� ܷ<ZYY)���ebb�   �M�  �#e�wgg�MW>_&43����{t�q  ����/_���_�~m�FVjO����l蕴��\��v  ��q�   pGiZ\\,��������MNNֆ��4a����s� 0����?��?
����#����K�%3�����  �!�   � A�L�dxww������4�X��;  ��h������� �ֽ{_�  ��   �aff�<~��t:�t�]=�?aw  �O'����B}�35%�  ܍�  �{�ɚl���m��-�;  ��5���;����~J)H�?�   �J�  ��d��L/--����r||\��v  ��P;0hyV�����r  ��   �,[�>|���www���Ez�;�~ssS�d
�  #)�k�4czz� B�G	��\411Q   >��;  @��9mgg��I'h��i��2������ixO�  �͚���P;0p�LJ?   �;  ���s&z�=>>�&}�l���c����M����e  vYě]����k�=�9 �633S��)�   �o�   }�����Ͳ��R��	����
����/���imu�1yvvV   �E���!�u���aД	��  �W�  �([�?z��N �����_�!�Y!c{{���k��  `fggk�=-�Y�+�����L3���,  �K�   ��{wvv���q���+�������:������'�c����   �B�$,�P{����666��   ���  `��ȶ��X[�3ia�fff�_|Q���U���<::r�  ��i@N�=�vaQ`��I��Y�  �O��   X&�3��	�i5F��H���Çu���Ԑ{��iw���,   299YVVVj�=��`��<�<�  w  �!�������꾷�W���
0<&&&j %#NOOk�=�����  И��}j�}~������8y  0(�   C&���?.�N�ݵD�p����ckk�\]]�	�������   �#�Ѕ��7�b���
@[4������  ���3  R�T�HXv_`�X&766긹����	��صH  FS�������3@�d�~��333  `X�  �L�/..ְl�ooo0���w�ی'O�����7��	�  픆�As��`���Rh��l�y  `��  �@��p�����^�t:h�Lglmm����v���i{  �W�Ǜ�������r[[[�H  j��   ����t��/���y�����=Ҏ����:�����{�� �����{j FE����H  0��  Zhvv�<~���wwwk+4�.�L^^^�#.//k���࠾^__  ���\\\��ϴga*����,���mrr�   ���;  @��Ungg��@��] �+;4lllԑv�4�'잆�N�S  ����������	~j3F���BY__��   �D�  `d2>ms	�&{ssS��J�&��������.d��a1  ����T�wN�=-��`Te���S�  �F��   ��bWWW�d}���h���I'#����I9::��z�� ���=r�+++�>9�� �.M�	�g�<  @�	�  �����:��	�����FG���nwO�=[...
  ��4�^����`�|�E�9�  �w  ����G��ɭ��]-�0���������xO�����  �(ʵp~6����I�.r�ˮ��  `T�  ��lM���U���j�]�3���z��%����.nIؽ	��g  �F	o...�	������ �M��[�ۭ  E�   cbnn����Ԁ���~���*�h˄���BY�rssSNNN��;�N �a��ل؛@{��8l  ƅ�;  ���$X���u�C�uyF\^^�	��� ��ˎD�5���J�����y	�g�F  �Q'�  0���Դ�%�zppP����I�L�g���i]��;=  �k݁�ܣNM��薝,������L  �  ���WWWk� ΂�0�2i���ѣ����Y=7� p_�Ȳ	�gh"x�, J�}nn�   �w   ��	�7�����o�D�h����5�ބ�� ��4��^3a���ź�����
  ��p  �����:���A��`ti��x��a=7������M�����  0�r�� {F�-�= ��rkkk��	  0��  �;i����,+++e�X�=x�of4����Ӻ0&a��7� F_�foZ�s?	��K�=;+��{m   �  ���ѣG�=J��%�����_|����3|���(  �W����ބ��*��i&&&j�DF�  �'�8  �AM�=n{{{5�
�K�nx����vO�{��%  í���nhO�0 �.a��O��.�  �n�   |�4�=~���Rwww�1w��2�"#x�t:o��u�� ������j��	��܏,j��έ   �L�  �;K�agg��Q���݁O��{&�3����M�=-�y��  荩������֞ & �G�  ���  �du��![�'X����U��{�H�;  w��e�ߚ0{^p�7r���6��	�  ܍�V   |6Aw�W��h$�޴�ׯooo  ?��r�Ȟ{�f�vv��˹6��	�[H  �i�M  po���{{{���{��V�uψ�ۛ���w `\%L977�fq`��333��iv�H�=��   |:w   ;�/M3޻Z޻��777 `T����J�=�B��l  ��   �;0�jy?==-���oB� �&''k�=�V�k� ^l�k  ����  ��k��	������/M�^F#��o��[� Z�[fgg߄�3������=fU�  �;   }���T��;0ho�I�ܛ�{3�� �^J{�G�څ��S������  �@�  ��t����tm��h\\\�v�&�~zzZ��� �]$�0d��LFB�������4�'؞�F   zO�  ��i�
t?88t�N�h��������r~~�&�����Y���)  � ����ς��� ��y�[e�`;  @	�  0P�,\^^�#aѽ��ryyY �Q�Ysssulllԟ%����ݛ�{�E; 0����	�7�����@;	�  ��;   C�	�$���_� î	�e$ ��b���|o��y �+�ܺ��	@�Z ��l  �   �����A9??/ m�@D�ݡ����rzzZ�oy�H�=-� �𘙙�a�ٛ��l�� ��	������)
  �a��  ��������tZorr�,--��H��;�ތ��� ����D��f�g6 �-��ܛ%��  0\�  z	�looנ���a����-0����e=�%�>�� �y�ʛ�݁��je/��   �O�  ��H�$#�σ���U���u,//��Y��v�y0�}�u^�ϯ ?��w��G1��|>��jee�g  ��p  �u�����E�����q�������F��M�{w�{ ���ggg�|66#?�F>/�`{B�   ?w   Zkff�<z�����֠{Z�5�(������������	�gd� �Ev4i��M{�Ԕi. �/�yf���T�   hO�   h�&� ���a9::t(t��0�[���v�=��� � �a�	�'�ބ�p���ύ���}  @{�  02���ب�\	�'�.�	�������{�ݛ��&������ |����^oF�ƞ�p�O�����  @�	�  0r�Y[[���������@0�#$���vyy�����a� ���$!��{�u~ �)�3y���P   �   ���C6[R���Ԡ{� ����t9��-����� |�z�k�������ҷ[�`�׹�^J�=���k�.   �&�  ��K�d���H����a^p?plγ����x�kw< íibo�ػ[�3���|6%؞���   ��$�  �Xi��N�6�X�N�'M�mM��{4A�;n ����ԛ���a����`��y���X��  F��;   c)m_iN����� �?�~�� |w|󳫫�������y�. 0��9���\��,  ��!�  �X����#a����rrrRC� Vw >a��]__�]�=_��=C i`O�mw{���u-� �M>�VVV꽀�1  ��#�   ���>|X���j����H�`���q~~��wi���{w��	�'$0̚��&��4����{m� ��|�����]�   _�   �%ᡍ��t?>>.� -�� �>777o��M�i�o���= ��`zT��nb�~�Q�k�,\Mc{v�   w   x����7[a����V�9��R|$�ބ���ς�6�w� �Kx�i^�n`׼ ?�g���bml��  �n�   �2ٺ��T���Y�w:��xH�CM�� |���kԛ��&��vp=a��7 ���ge��$�n�   �"�   )�dg$�xttT������m���Gw������ﻛ���荷�ֻC��a��g�� ����i�[��U   ~��;   �QBP���emm���Ʞ" |����n���k4�ބ��Gݡ􌷿o~�`����s����   C�   >Q�R	�g�6m�	�'` �%�&�{�a�w����i�ς-�x�iSoF��+����z 0\��>??_��d7<   �w   �L	`e�6��锃��r~~^ `P>'���{v�kwK��A��	ˏ��rԌ������ߛ�M FC>��3��   �B�   ����Bggg�����T��Vi���	�w�����<�ݣ��������������q�ͣ��_^��x�u�{������z�x��Ӛ t�+	�/--�۵$   �K�   z �og\]]����:��q҄����7�h󍷿���}�󡿇����A�w� !�>l�b   �/�   �Ci0[__/�������/..
 �{݁q��  �#�hO�}vv�   �}p  �>H����rggg���t:�   �Y0���T��  �K�   �gپ;���6�g���   �a333S�'ܞ�v   �5w   ���鲱�Q������qmu���*    �� ���|mk�"}   �'w   ����:a���tj����    �S�Q��=�(���	   w�   0D길�(GGG������    �Jv�[^^�����  `��  `��̔��Ͳ��V�����   �><x�.�O�}nn�   ��p  �!699YC�ggg���t:�   �)�!M�	�OM�   0|ܭ  @K�M-����V����   �!�-nee���  `�	�  @�LOO������~rrR[�/..
   @�������X��p  �6p  ��z��Am]�H�=��iv���-   �����</H�=!w   hw   ia��ܬ��	�'�~uuU   ���sss5Ծ��P   ���  `�LNN����:������a�t:   Myд�OM�    �~�n  `D��-���6������    �7??_��ikO{;   �
w   q���ecc��������v�+   �.eqq������}   E�   0&��V������=����    �kff�,//��vm�   �:w   CiyK���ښVw   B��  W�   0ƴ�  �p��  ��p   *��   0��  �'�   ��hu  ����   O�   x��V������~~~^   �O399Y���  ��	�   ��f�=��	�'��   >,�������:;�   �'�   �I��666j����i�w:�r{{[   ���zqq�ۧ�L�  ��p   |��ϥu.#M�	�����   �jbb��+'�>77W   ��p   >���dYYY�#����x���)   0fff���rmlO�   �4�   ��ʄ���f���(���5�W   5Y������   |>w   �'<xP�dϸ�����������   @[�~w~~���s�   �/w   ���b���V���Ymu�t:����   @dǲ���lOs;   ��   @_����q}}������   ��I��	�'�   ���;   0		����qyy�&�~uuU   `P<xP���k�}aa�    �%�   ���tY[[���쬆�3nnn
   �ZB��5О��,�   C�   *ss�{����p���TRKj���(���,#{��2�(3�$�A֑y�YA2��UR]��:o�Z-�պ��z8|�j���VI��N׹��*��nu��z�.   ����c[�p��   ߡ   )���؜�\.�F���g�Y  �����5j���  �\�   @z������u��y�c"|  �?QO&���=�   ��   ;%>>������M�c��z�.   �5�k�����i    ?�;   ����c���j�s{{+v  8`�ǖ�ۇC�$   ��w�   ���������r�,���5v��   ��#j���  ��%p   �J|�|���E����2��
   �#�������T�   {D�   ���w~~^g>�׭��G�  ��O�j��c   ��#p   �h4*�߿���#t��}�\   ���ze2��w���c\   �K�   ��x\���������=f�Z   �^D��������nj���   �a�   -����ݧ�i����z]   x=-j��=�vQ;   &�;   @�=���"&6�G�[���   /'�;::�D���    �M�   �%�FXq{D����u"~  ��D�   �C�    �nv�  <��   x,�;   �#��  O�   <��   �	��   ��   _K�   ���  �!�   �I�   �������z�  �"���L&����~   xw   �ҍ����M����r�,   �D�   ��;   �+9>>�suuUf��&v���   ��`�����;   �K�   ���x\����5p��}:��-�   oi8n���C�    �I�   ��F�Q�����X,������   ��x 7������=
   �[�   $�����,�����]�  <�^�W���6Q�`0(    �   ����ݻwuV�U���b���  �D��/�ɤF�q�k   �l�    ; �PbB�����f�  p��������    �	�   vP�)1���e�Xlb���z]  ���h4�< ;�   �.�   ���xvvV'���___��rY  �����6�G�>
   ���   ����65~���f����9  ��A���?�v   �}!p   �c�������|>�lw������ �����=w   �}�    b4�9??�q����f��b�(  @.�����mK{��/    �N�   p���ǘ�����=B���n�;  ��x���Ԣ�8   84w    �f����:�� ��-���i��mi   ��   �;���G�>�N7c�;  <]��vD�   �%p   �A�ᰜ���i��#t������   �����D�nK;   ��	�   x�������G�~ssSg�Z  8t���1�   �8~�   ���F�:����z6��	�c�;  ��x�	ڏ���á    |9�;    �&�������ͽ���Ƕw  ��g�t���`P    �zw    ^D��/'''u�r�,���5v�����  �+"`o1{li�S+   �K�S    ^EA-x���CY,5vo�c�;  dlm����"    ^��   �7/�������v��g�Y�  ����m6��D�   ���   ��1Qh�{���(x �9�{��hT���D��    x[w    ���W�U�����s�;  _$�c���������    r�   �^�G'''uB�٬L��:�w  ������A;   @~w    vN�I-R���� �	��vvA;   �n�   ����rYnoo���M�; ����=����=�q   ��&p   `��rrrR'�����]� �[�ƈ��    �M�   ���nx�G��b�8F @��b��c��q   `�	�   88�鳅R��b�(��t��5  �g8n6��q4    ��    ��A���Y��\.7�{�l6+  <�x�0B�6�ǧ�    ��    �1���I��Z�j��b�8�=  �X��j����q=F�    ��    ��Q4���f�X�	���yY�� ��E�>��lg�O�   ���$    x��޽{�����wƖw `��{��fv��   �w    x&��}2��ily �I�߉�=&6�G�>
    <�;    �����G���rY  ��-�m+{;�F�    /I�    ��-����]� ����{w"r   ��$p   �71���I�f�Xlb����w ���b���=&�   ��&p   ����a�n��6�wg�^ ��tc���=    �H�    ;�M�m��|>��6�����z��n�G��   �%w    �a-`�j��[��q ���F��> �16�   ��    �g����{����w  �����m�>    ��;    ���'�I�f�ZmB����}�^ �m��축���q.f   �P�   �@���r||\��E��M�Ţ  �'�oG�q��    p��    �-�;==�܋m��w��8.�� <,��Ո=��    ��    (�ɶ�+���=���� �����mc�ng��z    x�;    �d�M&�:]�w��6�w ��p8��qޢ�x     �:w    �ٵ͵'''w�/�:-|o�	 ����ޢv!;    ��;    �jb�m������w7�����w ^Z�׻�w'^    ^��    xs�!7f;|_�V���m��z�. ���י���V�s     ?�    �������ζ����cڵ��0�׍n�>�7׶�   �n�    ;�s[��}�{LD��w�ݶ�w7��k    �n�    {���i���1F���b�z<������    ��%p    J��'��'��V�;�߻綿<����w�   ���'�     �/���x\�>��{7��k ~���M�    p�;    �#�0������b�{��[��=�� �^�W���`�{�v    ��     � ���hT�s"po�{����xkm��v���    ^��@    ������7��~{ �T7\�N��W    ��;    @"-8}Hly_�V�D��^�����"Ho��}�z;��     ;�;    ��i1k�x<~��n����ǹr���#FoQz7P�>����u    `��    ��cC������t��n���p    �P	�    �"���F�������y�5�Eۛշg�~�    ���    �$_�~.~����]wϻ׶��Z�ގ���]o���:     /K�    ���X8�k���y7�o������u���v""����]o���h]�    ��     줯� �G���}�|�����4�?���5����b��w���^���������     �w     �"�    ��!p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�������o�����E  �q���?��(    �vyy�w���  �Z�����?�}!��?��o������i  ����w��    ��?��z�.   {j���mX            �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�      ���X���\ �/�������� R�����.�&p       6���?���ß �E>~���z��$�����UHM�          @
w           R�����_ R��z����K >��^       ���[ v���o��         ���           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
��k׎    �[OcGq          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          �B�J{bʪ�    IEND�B`�PK
     t$v[;mLP   P   /   images/ded7c6f2-b589-43f4-a4a7-c3e3242414e5.png�PNG

   IHDR   d   �   ��]s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��	�]C��;!��kD,!K;�S��6|��f��Q�,�D�UMՔ(�N�}�ˇ1�!�E;�� �.��b����o���sN�s���f�>U����s��~���O?ݷ�YBhҤI��m�m�'~�[�F�6��SO5K-1��� mF@ڌ:��u i3� �f��ͨH�Q�6� mF@ڌ�
�s�9����+n�Sυ-B����9��L�P[��r�-���m+ۖ�X@����ʶ������i3jW@��6ҳ!Ö25�R�k�������M�Q�2��i1��ѫ�q��ӫ��j��֟�v��9��ͯ����w�5�2+���O0n��_~q��v������ �ݻ�Yj��L�>}��K/�������7ߘO>�Ĝx���.��9��s����� 0��{�ܹ믲�*#`�?�� �YH ��2�������٦��,X����_l�( l@���m;ж},�FΟ?��}�,�U�L��g�Y���
����e�s�����g_t�E���G � b-���/L�� PtMh�2��׶-��tS�?m�ն�t��Ԛn�N�1�5nFx�m+�C������%�V������b>���	m�m������n��6@"Z��m�dj@�����
��~��|���믿68�����z9� r�8������_ެ���� �s����/M��0u`�1ݥ--$����m�m��w| ��/�tяu���~��1Ͽ���Eܿo߾Dp�.�[i��@P8�ѦfZ����m�珳����e�ٶ��^&'�駟�>���
��͕�:�����>��=��7�4�-��f�u�1����,��l��mg�8�1��� r�I'��f�v���34g�����;M�|&mi5��Ϟ=��0i�6C�q�M�* ��r�65�f�f+}KӀЙ ��l;�Df�����o;�@j}�Փ�k�1c��/��`�̀�4fOۦ����]���-M��~�]`���ub8NS��{�9����H�����[Ns�j��L[�j۶��dSKV6Je@0ֵ�f۶���0�̙"�v"$i�o�������8�;b�V���=�h�J�`le۝�J��8ї^zɽ�3���>*�@��{�9g^7�|s�ER9��dj��ʠ�$ cW��m��&�g@H�k���4���� f�9���;�������]�?��c�裏���/�I&���9�)�Q�R�`�mj`tY���D//���S�v�
0h��c7OA���k�m~�a7�^�����ѣa�G��(�FYP�	�����T?�M:��W_��ӧ�H�݁!�#F�p`�tF3��l�͜�@�/��(cǎu�	@A@�l��e@I$ cL�������駟v꾤��
q}���IH�(<� 
-����N�2@a�o��RH �PSӌ.s���t|I��H��k���}�B�Кp�(����K�d������6�\�@)�C��Z�m�M��fhn���Ɓ3!�ׯ���xe��O�  b�M7u��,��+x6޶�R��H�@;�Cf
��)0�4z�D���a�>��?���fԨQ.�B`B�(���Ds�}�Y��V[��cNZ���c�O��d��7�b���N30S�	����9 ��+�����̑��Y��`*}��"��|(S�Lq��ZK���^�F(�c� x��m��<PRL��.Uf�Т����!KF�R/�h�k�L��蟊�r�в���aR2�\Ä�Y<�Q����ڒq&E�e���P��*C��m���f�M61k������\���O0��Ѣ��Z���qϛ7��
R8
�c����s 37�q�9�����0KK�f`�H���� �K� l%�.�0��4?�����I:�����f���s�ꫯ��| k#E�,�d��y�����7�./����'JG�>1|�_|��J��a���nk��b��� �K&��l���h�߁�B3x�~��f�mܤMꩧ�y�>Uо�_~�	S�邧�mN��.����X�AG��Us��=ц]w���
�AR�N��  *����Oݛ&G�1SH3 �\`'O�����Rv����;n,r�O���jI��Py�{�$�����R-��
�]��^{9��>���3�/���jiL���x�	��v۹曵� �Պ̸��!L�w�h^�9�gv�]5#p��������KM}ߥ��#�j�=�9�}��c��x �RF�� um�P�p��E�#b�Wv�ֹ�&���j�7��3�j��� *~j��VsZ�u|>ǌ��=����*�#�|�t�7.�Rx�/����%�'�5�*�.B\�v�yg'���AHX�|�D�*&�1��.��A��18��_|х�1�Ì�\��G�?���T����c��#�<��~�����"�A�0�9��������4�\Q�QYN���6~���Rw�q�a�9- -aw��d���G}����07�%Y$pI2C�;w��&�>�r�-�@��>�B�.!�	���7ݓ<s��	�f�;����Ly1����t�����|_f
�Ǻ��B�f \��~���]�T���@ hX���otY�I}Bx�<���F�����wd�B詳���S��&9򬔂4&$��9�g�LqL�Հ��g0��O!����K���g4���������#������	izx~����i�`��7�!D"
y��������e�be5n���o��bbА,;�c��@V��+��Q��.̣oL������<P�t�]��7��<�T�G��@9�p�f�)�×�FyK�Z3@=��!  ��3�a�`>'���{� �]��ED��\��fHBF�{n��N�\�N��������a��rPxI��dUb��H9L��ƒ�0�|�>�}�?җ�� 8H
=��c.�mH~�O_v�eg-�*Y
Y|U`�}@0W{��Z�o�F�4�|
�%�'�IH��L�Ȭp_��Ic* 7�|��i��\N	�i�46@���I�WMq?��9V@�~ ��Z=n��f��A6f��:��.�.g���4S��q�p��&]��<�Lw=3�� �) ��av�5UEahY�~���Y�c��[o���l'`:ҍ�"(�ADe��l�=����g�}�����*I�-*���%�ce���Bs�,d9^�A��n�@�L��;nE$��h�R�=����㏛�/����M1]@~�h��dU�fLA�a|fP�����Ͳn@Z���<�=@���+j�� ��bz.��2'���"���U�I�裏̬Y�\hJ^�� �S�c�B��ZJU-��e �����Ҟub_�D+�J��7  �CI�*t�Yg9���FYj4�a>��Ѥ�tK�o�5W*7%h`��
)�B�v�ֶm(���}Y�_J��%�!A:�Xe�9�Gr�t�ĉ����wQs	���v\�V����k)`Ǉsg�X��Z�e���l��`8��Ȼ������G�:K���̙�U�|�mV���ou�g��T`��C�$���A���W!le�{>*� 2����!
 <��)�* ��T�s���e��|�2��HᡇJ�5�p�I$���{"D_��p��h�v��� CL�H����@+ &�UI!"L�����L�:�2o�}����F&��"8�K.�I��u�#��l��||��0\�/���Re�W5c�g�� Ht��B�2!�f�d4y�eC]�����>�g�ӶM�R:�>�:^�oW���4ҫ�����N[����3{�c-cٻ�lg�#LN}�Y�C�� 	?�����V�.�m|B*ʤ�a>QQ�xs�;�zx����ٙ�<b��+�oTڃc�Y�ʱ�� �`@�]w�3Y��wY�'�O�}� �?�& ��$�*ss�J�b��oU!�H�ځ��DIk�$a <�H�0E2m�;}ԨQ��|��,�p�gH`���[o5T˝Z@/�Lk�w�) ��Xk�"B�eT��':P�\��J���yHT}e��BG��������H!K�$ނpt�*B(�a�+
e��;�4x��`ۿ�G���̺^�{Z�`>㏓1�Y�&���!�hJ�� ��6���2NK��Ϊ1)C����P�:�A����{����Y·p���}oǆ9tBU/b6���A3��SQ؜�z��j5��-���('�<�:����}��M��ԟ�M���U�!�2M��>3�	&�`5��󯷭�� �F��h}<f)��ïY��*��{d�RV�B�>2�$!�r錎O*"ˌ�y�1U�.��P����e��z}ʔ)o�hm8�a�=�0/������ �/Lx��5e��ġ�!i���?�E�p��<88�{]u�U�}@ʙ��pI�S?v�y�чޖ�Tx�\��u��-_�F^�B�2N�DX��<߫�nm(�y$��y��h/E*i2%��W��A2b;�2�k{�O��1��09�AT��ߖֲڵ��Ϯ��T����rp��!�3\�E��#Y���Q�E ��TiR��h�'���*�%��s+E_��O-0�܋����V+��G�����o%q�3���f�Q�q�dM
�L����h@@�����*Bٰ���s&!�x�y����m�����^�U<���ٳ7����234�~�e)��Џ��V?@0��_̪%��v}�E�Q��4U%����r<��T<�ۛ��� ��n�7�j�6v������f��+v�]��f��S�eҳ4�mD��=�Jt�EU�� ��UE#9X���Xw��UL��P�U��J�H��R'��+�'��Ué��16/�B�4�E �B�Xu�
�p������g�-�_�y�V�R���q��Z@�d�.QѠ�9�m�v�mI}�yL�o��2k+8�d�?F𵴆� T{W����8;&�8^:�{*��H�0�f�� �Y��ϞY���z4�K��h�����H�Sy�H��ZIC�:�rZ)����{���=��Y)CHI�7�h��BƼ���X�W�A
a�v�}w�,�,*�� '3�<_E?A�T�� ��&�ʣ��߼I��=�X�&I�.�"�}�1����UZu��q��[V�'ˡ�O4�h�7
F��j��#��{���J3�Ѯت�w)�K%����_��0��Gb��\��G���bD[Y��"��l�$�2�������>��)��̏�l�t� �x�xƔ�Y��R"JA��"�	H�%yE�f}� ���3�8ô��#�R!�,z��W~�7���PY��|i��XTC �"���0�HM���[ːT�b��ʖ��cS�W)�� `[�! `*E&'� G�G�%˓e�T��p�����D�!
���
��8ѳ2q/2�D.)f�/�%�ͼ�1�V�Ę�*ά�����n�d�K�ْ�ԯ� ��j@$/��Rs��wI�4K�@�L��䐈��k�Du���RFDN,�T�܋yV���, H�h64�ͥԆH��g �w�1Ǵ�t������|d	��)D��k�#oU�`���Bb���OD2�vA@P��$���bj�Q�����Kv8A�?�F�b�LmX� p����_�|�V��ũ���7I֘5�
���	$�/���!��kb����H�}��g�)͚/ԟH+eSc(:\�~¬���\xᅍ
H�eR&e�2d|8s�!7�w�D�>_�����9B���ס1'�ud~���9J�R�����9	��f��>��;�f5kRJ�J���Mǈ�
�S�Nu蓼�FM��`��Pe�� ���b�T�;�P�4���q��$��R���s`:�0	ŧ  ۪1�����
Ig�^y�� �'2�:D�Y���������Q�O:*	&ss�×h;$9���T��馛�3�a`dU��(�c�5K�BH?�W=#E1?����� ���I�p�U��|��ᏋriI��DTY�Y2�U�L!Pb�#X?�S�QG��qy�NM%�-�REQ\{�w8��փX4��BP ��*�uR��'L�vg��*��5�����K;� /�t� &�=�Gq�370F�p�Pj�R�y��0��:��`(�c��CE�H���OAR��� �|�y��*�b)3F�E(��ZB�\����d����؂���K�3�׌󗳦�){���9�Y�>c|�V�Ul���^H?���y=���� ��Pe@��,��6�Ĉ�<��uJYT���	b��i<C~�_�U_ -��POEkh �'T�cf���o��g��3�����t��A�q���>��SK�u�}���ES�J�q�,����=�:'7��7ý���u�]�<b���H&Zb��H#> � e0��Cg)r��	LEs8RF$I	l(���=�Ȭ�c��������S��P��20:$�xpl��JK�L�?4э��&Y> :��ȧp���as��B@��:?�1c�`6���p�fU���AȂ��RӀ�ڝ�2P�+ԏ�@0��-΄$�D�	��F�ֹ�>I�y��X����J�fL���`�٬�S�������/��L�,��]2n���~z '(�S�߀e;Ơ��Dh�*��\���=+Y�M�� ��,�=�ֱ�|N�*WC���� h~�)}�g��'V���Uh�Y�ʼj���tVc�	>��*�4�E3d9V�I0s���g0Kg:����b2�k�j��H��7�nxm�I�r�8@B��/ӤL'raЄ��:�T	@���(-�)��/�pT����P���@(c��Tꖟ�&�J���*1P��07V�#�Af���2� �Tz��1���I�5D+����03���/{�%�k��u�g�p�g�{�X�݈9�UIR��S��F����V` p3u_P�h�JF�䪤-e̗N.���akwV�.��0/��'P B~��E�����B_�H�O#5�-��w���p�,�00��ŝ�Z��w����)s_�s�\�<TI+�N����*i+j�������c���\�͑�N )�a\㕾�͉���\��*ve����hU� ��{��nD�����>��f��q�����7��왏\���^
�am��@�$^������_g�Dݦ!�8�33Vфj�t.���D�BJ-4qM٭*�ù� ��0f�=�s�Ea+ �k�L-&�	L�}��iu �:�(G�Խ�b`�~\E��{0O�.V��+�20��Ι0�$���	O����vf�.ơ�e�ԭ��d��"�E�FU�1k� M�6�V�����K��C��V5eh�~FI'�����K]`j�zHap �U��\д��P쾲�e��c�� .�磱�8M<���<VmZ��� i��0�&G��=�P>Hztܑ~L����Vu�
���͟Y� @ `�V{Q�"b���o�J����11�����6�����]�������H1=RI�Ik�z���<���J�L�\�4*��)ӔE����iQQ����*`h��HfLK�0�_i�'�.��t��L#�z0>Ӷc����g�{J���%��,�=A> ��z'~���hk?7�N��Y�����W�+�r������Ib�C
h�m��=L퇙���ƿaM�v<n`��;�� ��v�����СC�6mڂ2��Iv��������y䨉�BJ��v;��7&�P�d��zҧ��5k�2�Z��j��DV�J+@T[�@V���� �vޤI��b C/�z�w��� �~��"a~I���?Ԉ�v`�mW�'E���ߛ�#v"�e�����s����%��, ��v���El�z�����Û���_��%���g�������v�F@ڌ:��u i3� �f��ͨH�Q�6� mF@ڌ:���/�5�a<�|�    IEND�B`�PK
     t$v[U�p�	�  	�  /   images/42e39361-2f02-4030-a678-a3271aadd3f6.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx�����e}���}�m���N�s�	!"�UD�R)�-D5t��9�s�N�ҩ����L[�N;��g�t��3gfN;ө��V.RDQ	&$B��U.I��H�o�����jEd�<k����Y�, �F�k��z���   p�	t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t x�kC��m��T:Y�YQ(dˋ���$���4)�'M;�$Kz�&I�����Wz���?ϲ��eI3�餓����]���C=��~�T����v�ggó�N�̒%#�O?��f  �@�!�B�yr��=�Ph_*��-[�BgA�Ю�J�z�6�i�`�h~��<�F�]��t�S���Vi{�Y|��L�v���]�_Z ��@`hm�z]��x��J���r���Tj�����X�]\*=8��-I�\��+���Bc����?���������fyo�Y����F�x�[����s�I� �Q'�
w�q���+��V��ˍ����B��������Q����=�}�s�5���f����j��u��ے���  ������ޫO-�����̞].���uE�>yT��ǫ�V*3K�G���=����3�<6��o]�cv6��ʦ����/��  ��@_۲�ݥn���W*��j�g�jS'�J�.�,�B{�V;p�wV���{���;Ϟ���=:=]���L��'���q�7t pDt ��C�Re����ڋ�����FF�>6M;���+���g,X�|���sk��>��o��V��,}�'�	v x�: ���������5���E��w��hQ>���PhW�����?�-����#�\���TmӾ}�.�覇 p�: �ٶmCyzz�򱱙+k����jO�Ȳ,����.����珕+û�z�=���[fg����}ڴx ��: Qز�]KK�}׍�M]Z�=tb�v��m=�}�;��.a�e���x䑟�Ɓ���t�G�<�CS �����/_�bE�����k�?�,�V���.t�;��㏿���~��g����n� : �l����ΞkE�3�5�m���7/���O���<��8p�vS�1���L �!%��s�_��p��gll����N�R�w�i��p�޵���)��C]t_/�?�v��7 2�9s�W��ti�����Tj���+��hў7��������-�ܾ}�?���� 0: Gԡ���w��=݂O�B7�"�J3��/��vٲ��<r�_<��Cg�y�ǒ���  J�pDl�|�I���?��R�� ��$��w�n��;���m�.�mϞ�zӛ>�x �#�xY�lY�����=:�詽?tW9s�T��W՗/O����o�o�ޅ���s��K �@�E˷��p���[�����Z}bu�y�-|g����ַ��Ԟ=�������3���w��v�]��~q��'ޙ�p��j����{����k_��SY��ߟy�ܫ@_� �D_��[_�l��{���,�� 2����+�������_�m��c��v�'w �#���/]qҊ��5>������ �+���K�����sE/�?�o���\p�'� �: ˦M׬^�p/�w�9M�~V�wҴ]���/�u�7�q���]�[B��y����u׆c-���ŋ�uE8�\�v�K�캬�}����-�n�>��K.�Ԟ  � ��n�z�ʕӿ�t�#W�¼`�������.ݶ���<�d�;��}�@ ��t�!�u�u�R���/Y��[�9àPhV�/�y��xy���_�������	 �0�����_����\,�.
0dJ������_\��~��w���sι� �2�0d6n���c���۵���r##S�7�?��߽w���}��� p�t�!��[�x��.^��M!dI ��^�J�~�>x�''W��ڵ� `�	t���C�T����o._�ȵΙÏ�-,^�����]��o~s��;��|� l˖+7����E3�8,�bst���^�h��[�\��k�~��  �@����Y�lپ?�Yf;;����1k�<�?��ok4V�ʙg~h* �� &��>1���S��, /K7]�d�e�恍��s����7}, �� ��;�>aժ�8:��kpD�ˍE���z袷8��"�\� }.�ޗ>����Y��w
� ̉��ȢE{�;�����_��[�k �#H������5O>��?��8�� ̋B�Y?昧��#��i���/�ŵk?�3 � ���֭W��+�|O���4^�$YV(�+v�;;��3�ڦ����^����{���g�}� x�:@�ٲ�]K.��.|�� G�t�\>$O��Y�=��t����n��d��^�k��Ph�֬y�>x�x��O.��6��x�:@ٴiݕ�V=���� GH�M���@7IBH�$Y\(���R.���1��z��}�쏷�����l��Ż.��kwl�r�?wo: /�@�۶m(��.]���z9�^s��|��T��G����	�T?��?�҃�N���wY6cy��R�^�z������/��k^��%��}���"�"��}����&�0G����N-��M��B����Qɷ�w��v��GZ��C�^�u��i�81�����������^x�c �@�X>nb�_I�N)��vw�_�ߙ&i��X.��Y���j=��t���v�m����O<����������9��xK �� �"�e˻K��#�t�S���[̱nwo7˦�IRK_�N~~�\>��9#���N��p����P���J���{�?n�v��N?��� �'� �ٴ��K������NȜ�ee�3�$9�����4]Z�=���y#��V��v��V�!���˗�����������ڵ7� �:@D6o^��ի��w�RcA�y��+������$I�եJeu�\����y���<�l��h��m�=kdd�����p���? �� �"q��W����O��|�T����}�%�C?|IRI��S���T��i�h�Z�Z!���+���V=v��-W|`��[> ��xp�m�z]}t��?]���sE��s�,keIR���i��P._T+�������֖Ơ߱^(�G֬����ח�u�i��Ul |?�p�u׆c���p�z���nȲg�I�z^oH�rR*�Q)�^S�Ϫ7�[��Σ�����%˖=��G���7�|�Ϯ[�� �@8j6o���ի���Rifq�H:���(]�w�����R����j�3{h��`��Ͽ�կn���/�ׅ��d `�	t��`ӦuW�Y���U(4�"�e;����H�e�Je]=?��j}��n�����ju�W����7���.�� �P� �l��+~qbb��G���J���y^Ρ�$�9�J�Z�|^%?��nokfY'�r��������-���ڵ7~* 0��9�G��鿞�x����(���f�������#$�X�\��Z����ln��כ���=w�O�ۯ~��5g�u� ��~��m�6�K��:>��"���.п+�C+�g�B}�l���VI�-{��������N��/ �N�?|ɖ-�j;?6:��� } ���k+!bI���W�K�״��;g;�gb�{�e�ҥ�^���/<���Wװ�0�����-Y�������Ng{��ǡ��?Sl��v�gپ��ŋw]��#wܰmۆw�~�� �P� sd��k��^��'�����H�MeY���$�/$I�xB�X<��jmm�Zw�� ����}�@�ᡇ~�ړN��F `�	t�9p���^�f͎�+���P>ͽT�@��BR*�=R,�Xj6�i�뛝 /d����=x�ܺ����y懦 M�a_���w����|Y�>u����Ї�dA�Ry�h��V����,;������������t�mW��K>�' 0�:��i��N[�zǇ�{���nwG߯>�[���+�Zw϶�_m���z��q'��}r��k�y��|. 0�:��q���{���V*5G��nwo7˦�IRKCK�RR._P-O)7�5��<۷�^�M�Y�z��k�;�?�����#���{��ԕ+��I�(��}���	}�ߕ�K
##׎���juj��>��͛7\u�7< (�eڼ��&&���b�� � �vw�C8�ơ!r��+J�Vӟ��JχO�^s>v�]�v��7� ��2|���׬Z��#�RcaIRM�l&�C��O�.-����h~6�ټ���7�&��q��7l�z��Lw�%��9?�؝�W*3K�P(&��*�ҙ�F�3S���2���y�,ke�9�0p���7T�����[���`�Uz�~�����[o����.�M� ��l��˖=������0
�W�*�7U�d���+�+j��G'�Ab��Y�l;IV�6������������L��h+��z}���zU��m�~��74 }M��H[�lX�t��V�V��y�|q�X|�Z%Y_����d��X���S.n�RͿ�k���V�3�6@nll���n�^���s�7���� /­�^R_�d�'j����X<�T�\\�c�G��$Y\�V��ff>9Տgx9<����f!�����%I�tF�PX^���y:���7�{^�ɟ���� @�� �)�ޗ>��v����J�zR.��V,�WM���R��Ƒf�K�����<ݞ��oK��J�]�I2^,M'���ώ���6��<�W[�/�}Ѷm������{ }I�����K��]X�tj�T���$��^--���v�t��v�u@�Ԛ�͍�Q(�*�g���K���0��#W���Vk�l￁�/V�xf�׾v��׾�� �;�0|�k��wɒ����$��O��������rq5��w����@�tv��G����TzM/�O�|wx�`I�r���4]�6�΄��Jϲ,������{�c�s�g }E��w�}�;V���À*V*��kI��el].�]mf�/&���./M�Mg�V��4
�S���ٕ|.A0��	�4����짧��{;I��c����M���q�y7� ��Ǹ���oX�f��	�;p��{J�sG��s*Gb X��ґ���gf����Xm���'�����7�m���J�.��i��P��k�Ѹi�_v�
�5k����o_w՛�|���0P?@��;�������Ӵ���}�,I�I�|y�X|��>+M��;������.GB���Z��íb�U�PϷ�/��z��IGF��7���y���N���[�^wřg~h* =��#�w�/[�ԟ���.�P��E���$��x*O(u�獴Z_1�}(��p/�����r����^��Q��T�3��֦�����&״�O|���7\�t��	t��_���c���jujU0���*��G�z�v�m>��t�����C���N��b��J~�"I�0����$Y�6��M�����?���G�m��{ Q� ?����������$�^4��Z,�:O����R���e&;�g�����z�uo���f�\�`�T:���>W*�Z�?ph6o���c�t�3Wmݺ��3ϼ�� �� �g˖u�NL<��0@��֋�+��1���_��?wf�/fٔ�Co��l�:��l+��W�|z~�#M7���>��x�b���ܼ���=��[ Q� �q�W��j�S�!��ս�:t�|}=IF��=��Yݑ����ُM��*#s���ޞ����b�ryme��[̵4�(����韘����B�]Y����eˆK֮�a  :�g�������I�Ь��_yU�\V�W���ב�+���%�F���w��e6&W�^VM�e}�~��5l�����T�S D�R�^>>�����= ����p���n��A
W*�]�����͏�b�r����jmi��,�ݙ���d���J�t�H?��'�x�V�vtf��Y�?�H�s���_��g��W DE�C�k_��7,�q^i(�/��JgDww{��A�����<j�;ߧ��͍N��v�ry-I����$Y�V�����0�e���g���-��_���O �!Ё��{�z���S?��I��j��	��|��e�^�Lf�.��������'+�7W�œ"����;߫��33���}Gz7]�r���~�����曟 DA�C�_�jQ���%I�oW��F9yk-M�-����RU�o�E��'�`�5�57Ow�;����~��G�V�ދ�E�ݽTj�����,{�eI��h�N�a"Ё�u�1��s�4�8��$����m�|[��
��ȕ�H��T��~X���ً�Ρ�^�C������G�7:�����o��:���x3p��w���h��熾7����"fq_�H�ե��|���� ?B��\gf�#+�+���|�rh��5߹f0�#+V<��l�r��׮�ԝ���/��_��'ML<��}w��_�j��lo'_-�#�Q�h|r�\��Z,�:����#��md���#�(#=?�b���u�u�y懦 G�@����o({��T(�GB���ޯ}�ߕ�3>4���v�!�3�Ѹm����-��8���>����J�aC���JezY���{O! p�t`��z��[�8!��Cq���o�}����\^���>��m�ֽ��{���Z?�˷��W�"��hg/,Y��[��׾�u��> pTt`hl�x��+V����wV�G���a`Tӑ������'�)�^@���V�;=��K�o}�X<��e?]m6o�u�B�{����ڰ���o� �w
��zI}͚=��TK�ZR�^ݷS����n����h|z�dw~��8D����\w��N�3��k*��k�֖F�P��]��������y'Ё��zu��+��%�O�J���6���(_Qʲ�G��;g���3���O�ғ��w�^._0�Gz��p+Dh���_��t����_ �J�o˖�߸l��W�>�$#�8�h��\�tv%��t��~�,�ݙ��W��>���$��,;0��<�Ը���޳y�Ϝ{�� �@Z>�}ٲ��_��'I!�����鲾��_�<\�R�v���eG��B<��=�C���.��U�'I)�T�V����d/ԣ;�Q(4������? �7h�������ա/%�\^׋�ե0T
�pɇ�}�.��G���'�j���ݙ�|�?�~�Ѐ���H_�x��[�\�a�ڛn ���M��v���O^�T�|Q�X<��P�z(\>��vt�B\�lWgv��S�J�ݽ������B��j�q�t�L�e�ʕ�~c���n>��M �@֊{�}�v�r��\>�R*���X���R��.���E���������v���b�r����j��d�Rifq������� ����@ں��_�׷��P��z�T:o$��pɇ�5����s�
�ۦ+��j�>��G��7�t��:�����%Kv]�q�_p�-� �)��M��Y�bŷ�A�C�B�|I���\�?��v����4ٝ���~��$c�����W����ff>r0˦"�2�MW���;�_���k����F�9$Ё�3>���
�>\�M+�����΁�sh�{��w2?k�'h��i�颴X|u_I��5`]}v�㓽(1�V�V�|�_�=�` `�t`��y��7��?u~�;ŤZ����A�-����[�33q0˦#[]$F���g�t������N~�Z�5�BaY!��ї/���7^�g\��� s�o~h�U����|;f�3���s��K�$ґ���gg?6�eѵ�ɿGfg?3U��k,��	Q�f��n����?�!y�g�L�>
�����{��� �@�W�z�?}�U�ϔJ���J��uj/V��,�Jo�5��Fw%�Ƀ�Ѹqjd���|����*zݝ��v:�u�!p��3�C���y}��%{�r�]��:��� 8�:0�kCuŊ'���BaU1��8l��Y�\�WR�<���;g��js��ʷ�g��^��!�����v�֎�nab��zO� �8�������x�#IRO*�+k�vgs��G���N��xtWR�Vkk3M'���)Gl�J~^����-���6GFG��~�=�������� �%Ё�w���^�t�ΫC_I����^�Gv6�_�߾�����d��w(�������L����$_䬇n�eS����v�m��cG{؇NL���m�6|���oh ����c����4m��uJ�ҹ#izl)�2T�J����̇�0ԭ�aif��-�##F_x��`��K����N��{{O' p�t��m�t�ً=}n�#���b�|N_}��4]R(�+�����t��4��4���F����Z�|���l��Gk�ް? pDt��-]:���t�Z�T��5;ߢxY�l��j�=�n?!�9l��g�����s�Ph�+�����_ ��������;#��r��j����
qjg�����ݍ��"u�8?r�.�}�m�]��K.�Ԟ ��&Ё��t��ik}�X<�\,���,���o��;gC�X�B�]]�j*_E�� ��&Ё��y��7��=��O�O�d,�T����y��h�1�e���,Y���7^�\��� /�@�Ҳe��z�e}�z�_�vY5�:x��f���Vk[Ӥv�S~������{����E�}g˖����=yb����J�-��jW��H���Z���3Yv�vv����{.߲嚕k�~rg �%�@�Y�d_��������ÖeS�f�3��C� �|�^?�[���8 �	t���}��o�ן<!�J%��^���v��f���١����dӦkV�w�'� �$�+˖��ՙb�R�x��퇥�5�_�m��m�/�i��`�d>��=��D�}c�����ן89�$I�埲��0t��;��-S��g͡ύ����/_�n�g ^4���˧�y�{�K��G��fj�OphK��f�� ��B�U;������ ��&Ё�p���^16����
��R��r�eY+k6o�6�ҥ��y��~��ko� ^��+�����>x�JB���ji_�����F�3S��3޼� *�f������� ���ov�a��g�uI���i�B���/ �v���?=¤��0��,y����y	Do����f\+&��y#���~��h�2�9�z��q�7����so�l �	t jY��t��[�}�T:��$c������f3��\�ðX�d��~� /�@�v����5kf��荦���*��e��fZ���*<���ןr�7> 8,�������@�|�H����ݬ���L��M��P���_�=yO �t Zw�y�	cc��"�$�
��ɥ������^���8�!�p��7o����ڵ�ŕ� �A������
L�ܡ�p�U��^���s �JͱBa�����3 �	t J�_��0>���C�
��B�x���������8X�߶p�����@8�TQ:��ɟ)g���o�7�B��}v���N�Qq|����W�G����O= ��:�ŋ��"W(�*��p��۲o�9����M-�|w�ɯ ~,�D�_|�+GG�|u�\�x�kվ���4k �B-z��,{�o$����$Ё�,Y2��+���5^CC�4��͍ ���Ƣ{����ӏ ^�7�@t��\"W.�Wq�<�v��f���� ���O�� �~,�De���o.��X"��K�4}�П=�t�����N����dll�7�|��u�>{  �#	t *L_"W,����Y6�m4n�ʲN 8i�)�\��L�� �H���؁sCĒ���J'��y~��-�Y6m�xQ��&����:�����r��E!b�♕
C�z�l~i&�� ^��у����Z��?��� �@�Q��"�$�P*�^C��~��j}�uj�K������������ ��"Ё(d���;n�z{{�pJ9IjQ_�6���ݝF�s&�/���3���#	t 
�7�s���7���J����,kf����
���9����O۲�]K׮��� ��@-�}G�X�����ˇ�5����L�����)I��ry~'� ���}�	������	+����n��V��͹s��=�os� ?D�G��w��ӯ|es4D��
'e�gY#�����޳ p��jOں����g~h* �=8�FGW���J����<�W��ZwLg�A[ہ#*���j�}[��G �#Ё��^��|{�)C�z�n?�j���
 s`ll�-A�� �U7^��V{lu�T���i:QC&���l�> �H�>yf �tਪכ��������<�Ði�6�fٴ�����Tf��u�U�9��O? �6�U���E!b��ɥ0d�lo�ݾ� �X�>{U���8j�s�ګC�
�U�$Y8t���/�dY' ̵���7 �G�G͝wn���O��z�Ba�V���G���� 0���n����e���5� Ё�h|<[���b��!�v�l~q6 ̓4�/.�Wm~,  Ё��^�:;D�PXYH��h��ͅf�F�p�90�FG��m8*�m�P�V^"��'�����j��W��]�6�,��&Ё�bjj����;�n!/�^5T������,�q�0�FF&W;�p�P��Q�5�"�$����C3�=˚Vρ�&I�����O��� ��@��ju�!R��+�굱����sਪכ� Ё��Z�>!D�PxE�[�4��@���3 ��6��R��(�?O���P��������W�<!�ޗ&���$5�̻Z����BaM�u������Z����G]�Ю~�+���{�� 0�:0�*��ׇH
���n?�ʲ)��@j�v~�@��м�Q�Μ"U(;4������ �Zm�� 0��(���ۑ�疇(��I�p(Οg��N��� "Q�� ��@���h���i�P����yMl�h�2= Ģ\�]��C�T9�?2ZC�f�C���"�����51�Z���z+ D$I���{<�� 0����(�j�ur�T��j(��w:5ChX>�S�w�s�Z�W���+C����$ɂ(��i���Vρ(���N CL��jddvU�P��*�\�Mw;���Q���0(j�7_���5����Ba�Ploo�i�� 1*���`�t`ތ�&�H
C��C���*��c7^���>�\ B�7�R�!JIH�e趷�˲,)����� ��@���H�U!BI2��P�q���`d���+Ё�$ЁyS*�&B��t�����:�Gmo�W.�� CJ��X�]"4��κݧmo�W.�W�!%Ёyq�]��҃��4]2�����lgY' ĮXl. CJ��Ph��il*����N��9����x R�i�:5D(I
�7�:��:�Ҵ]q�0�:0/���+C�����Q��)Y�̺�g�o�F�6O��"Ё�#Ёy���!B������p��+##�{�� ��@�E��\"�$����v�ہ�R(�� CH��Tj-J�a�g,�}�\� ��@�E�܌r*o��A���@_)��`	t`�]��B���Z�РOpϲ��,��@)�����;����^*F8)=�z}����c��;�R'�u�@�\�يt@\-�F�����e���'M�� 0�:0�Ҵe�;�^�W�kC���o�	 CD�s�XQNpat}�@�R�3���X "�s�bwi�P�����^�gY�|7 ��J��Or��P���+���C�Ҵ>Ё�eӽ@������ր�#Ё9���E!JՁ���t��@�*��%`�t`�
�(=I�����t�9зҴ����#Ё9W,v�B�F|���t�o�~vDy<
`.	t`�%Iw$D(M���[i��:��R�Ri��w��e� 0d:0�$+�%I%2[܁~�$�~�0w:0�z��kMq�W�ChXA�V�g�@�N�o��A��qz��|��;Ё�U(��(�4���Qnq����i�[I�}*0|��s.�3���y2�+�!�:з�A��@�A7�@O�4>[܁�%Ёa$Ё9�{�]�g٠���ZVЁ��e�������̹}�ϟw{�m���+�� s�0��O>�[�]���l�?I�[:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@� ����n%˲�h~i�t+�� x �t:Ya׮沣�5��|v��ʳ��'� ^@�^�n6�����^ `�	t �c|��������c �@ �	�.��k��F�; `�t �� IB�bEe׎3+��P 0: �aH�Н��E��D�
 �0� p��Ť�bE幝;�?<�ׯ0x:� ˲�LOw���H�(��|���;ɗ-+�>�ׯ0x:��j4��]�K��P
0�j�t�^�L��?��k ��0�ff�#;w6[pp##�����G���5 �4�0@:�N:5ըu:-�x�J:�OV?�_��� 8�:��h6ۥ��F-�(��F���gG��p� G�@�sY�%SS��v��9C�X�+ʻ�k�B\���"��X��.�[ڃ���^w&&*��������5 ��Ч���f�mK-C�q^,�Q��w�+���*: /�@�3�v����gY�I��
u���B�zQ�>�lc�8��� }dv�Y��m�Ͱ��=W����<ο3$� ^����n:99[�v3�s�l��򮑑�"�e!y��r�8:@�\��0[����V+̄�q�쳍e�f� �� �r}�n��Ҟ���t��s�5���v� ��!ק1�-*�[��8"�kWc��L�� �(�ק1�za�Ѣҁ�={Z�SS��  G�@���� �z==�xq����{[�l/ 0:@\�!T����e��!R����h/ 0G:�Q��48�RIg�/���������k/ 0�:�Q����	��1���11Qy.IB"45թ���\ `�	t�y��4��RҌ9�gf:#�v�s �@�G�O��Q,�V�i�!B���ʳ�6��`�t�y��4��(�LL�<W($��F��g�N������V���[-ɒ�o�`v؆d�ea	��H�,����xϙw�L�03gNf81�I�Ֆm6�%��a��W���ޫ�k�����V�mY��ꮪ���~Nn��2������S33M� �U: tǧ�en���ض዆</�U�G��5 �* :��Ӏ�Z��T��DC�Z��ͩ0NV  t� R�Գl<F�eKj�u͖h(�rS�yp �~ @��!Sځ5�q��Xѐ��S�/�� �  t�ؘ���Zu�P�13Ӝ���M =E� ����CCvE4���f�^ ��#� @��K##βhjv�9�h� @:  �\�,��:%���|k�^� �&t  ���8�LN�����o�R	� �Ft  ��2����h�X��eH  ��  6�뚍-[�y�T��J%D  ��  6E*e6�nugC"�P��EL  ��  6̶��9�k� 3?ߚ  4F� ��,�mKϘ����z=H�ζ&  ��  ���Ql���X�����=�  �9  �Ðpjʝu��Z�33��Eb
  	@� ��8w]�%�О�nN� �$!� �zE[����i�)
��Rq�b	  	B� �u��L�g�V]4G�y�`c*�� $?�  �qsr9�&Rq����)�G  H   ���84dWDCQ$��Ls2��  �P:  8�8�K##βhh5Λ�0-  $�  �P>o��Ɯ%���\s��3 @��  ਲY�:1�,���8��  �t  pD�Y��tDS���H� �>A� ��I���Ԕ;g���Eoxy�  ��  ö��u�;�k��J^�T�G �>C� �G�q�mۖ�5M	EC岟+�1 ��  �-��`jʝ�,#�jAfa�  ��  �0$ܺ՝q���Azv�5?5 �>E� 0�V�<�2=�P���s �  � l����fK4�y�=3��Eb
  }�@ `pE[����i�)���:x��5�   � ��w�Y�.
�Ț�nN� �AB� 0�FG��B�����(7�8����  �@ `��K��NY4Eb�8��(%   �R(�ˣ�NI4��|f�9�j��  0�t  D.gV�ǝ�hjv�9�h� `@�  �LƬMN������x�f �F� ��\�ll��΋���j5�  �@ ���Rfs�Vw�0$-.z#�?$  �@ �_ٶ�t��R�+,/��  �t  ��e��m[z�4%��~�X��  <�@ ���Ql���X����� ���M  x �>b�8w���Azn�E� p:  �#1|ߏ�аLӐ���}����k4Bwf��%~j  x ��e2�R����i�ѡh�2���,k5�W~�\��ff��9  O�@ �d2aɶ�ֱ��0�0\�d����W��*�x˲N8�=/�U�G���<  �( ��s�`9���f��(����m��]��;���Wo;���Ț�nN��X  �� @��nXN��z���8���j?���SW�]=���c������ �~ ���L  *�
+�U��{��)7�Z��  p\t  �q�U�PI��H�  �� @��v�H�òh�^7���L	  X �����vlM���p�  �u#� H�[�l�$����!�7�  N� @XV�e2��y�a|��  8a:  �3���f�b�45�f��̬  �!� ИaD�J�GZ�y�edZ-3/  `�t  ��*��HEC�g��MsH  �� � �P��¢iF�h��M�^7�C  �&!� Ќ�s5rnY�/�}#U��8�� �L:  zQq�dۑ'��ܩ���: `��  h$���8o������u� �N!� Є�ˎ5DCahX��9*b�  :�@ @��S��.�"�$� �< �s���J�5�P�Y���q�[  :�@ ��l;���aE4Eb4�H�/  ��� �Gl;jd2�hJ��ǹ#  �+t  z�4�V�%��J��)  ]C� �eq�{�s�T�n��
  �* �.2�ȏ�h��k����  ��#� �È����{��  �:  ]��\�Gz(j6͜�9  =C� �qz�y�edZ-3/  ��t  :(��q^4�(y��n6�!  =G� �!*��n���!�7�z�6   � �l6*�v������M�  ��  t@:�q6ECq�;��9�9y �Ft  6Y*�'j������u猝 � �M�J�׍j��04�Z�1L  �!� �$��\7�����0�s  �F� �	'���aY4Eb�8�#�  �- �������hH�y�n�����|  4�k � �0�؄k �f�Rg����n�q�;�����T�m[�  �� �(���f�o�L��eE^&�{��)A���+�R-�N��\�� зt �$j���|3��f�| �f�g2A�0$���p�)�
�F�Ѳ=/��y�c4 �� ���<F��aDA6j獆5��FZ�w��j4=�q�l6�h: � 6@M=m�<+CF�F��y��f�a�=���Z�޴Ջ��|�3MC��  �G��	bJ������\.,�f��#�yfN0��5����;���F ��!��0�}�8W#�i9���22�g�E��Y^�3� �� �������|ɶ#O4�yf��4�KMyW#�B�)� �`: '���L&,�q����6�`�Y=j�{��f�w H( ����*�-��q�`9��h(��tj5c��%#�f��H���^:�h�W ��t 8֛�T*(�RQ]4�]����A���Ն��˹�K�!��(Xo>�R���QM4JZ�9���h��bc]: $� G�z���JE5�����S�Tq.b0�Ǵ�.}h(Ӳ,�H �� p�j�\0�l;j�nP�8�Vͱ���O��u�j�8�K �� �q>�,+l��ECQ$F�n��8j6�:/=I���~��w����~��?�z�A��!l7�L3l���EC*�k5s$G�P�ǅadd��lZ'�t��������Mo��  � �qn��FPj�mG	��C��.r�P�i��i�4Bӌ�������כ��3	;���o��q�߾󝯾��k>��>G�h��S�m�-q�y�Q&h���o娷@���]�l'.��û���ϧ=�\.W7�ƾ��w�{�)��M� }�@0�"�Q0��M��/2���T���{n��-��{�[���E�Hꦔ80��q�j�������m������ş�O� �S:����R�;##�9 �����Hߵ랳���|�o��W	 �!�@Qq^.ם H%zC8 �LI�t�P���W����5�}@ ��� �j��Q��s x��HWk���I�R�15�����O�z�?�S�>B�*Η�� ����S���W�>�>4T�j�~����2Φq �	�����W��� p,������[�,�}���?}� @� ���r��R7� 8.jw�J���~N��]?}���_�WW_���* �t }M�`�M ��:'�0�(�s��BnY�LM�����{n����{ �@зT��L ��F�e��ٔ����׭r��w�O� �@Зj��M�����M�4�(�v�Զm����_���/�� @�� �N��Y�R  ��Zm8�eD�c����O��{׻^��o��- 	�,���6�S7� �T�r�QǯY���l;0FF~���o�G8z@R� ��:�\�@
 `�EQ�{ljx8�T��u41���}��w�O�. �@:����:�PϻF �A�#]�3�w��Ʌ�_�'W\}���' �0:���vl�s �<ut�ڈSם�'���o������k���) � :��c�v �.�wv_J�J?�z��"�!�$��a�v �>�!��X�����������/~�o�� @BpS �Ԧp�J�M� �G��"���h�qcx���ȵQ�� �$��1dS8 �����^�ϧ=�жm��]/�����W $ � ������� ��� ��Ɨ��ѷn��+��~��u��xX @s:��Q#6�S�@�jӶm+Tǉf�����x��ӳ 4G�H�(��\n� ��ܨ\�k�}۶��񶷽���^��� h�@�(�j�u� ����Mz���8������ ��t ��n�8� ����t];������{�;��/���O�/ M� ��� �?]�^3M����5~J��� ԴI�����l�Fó�iG�]�'&�w������_* �!���͞�6) �D�՚�:zM�]������o���=�ڭ� nxhO�# �Ĉ��PS݇�2�Mu]v~����O_# �nzhMM�T#� H��Mu9��f&'�~���RF��@��0��z���) H�J�錎�M���Ȳ���uk��U �����8�� �K}�wø�_& ����@��1z I��qj������W_��� 4��/ -U�M�<�>�6�S3�r9W���CC?����@��vV7 @_P3��4w�2�E���˼���?o|�'�Z @: ��jLm�~���
O4�������@�n�hE��s� ��V�W�f�miu���ԃ�o{��_x��� @�� ���9 �/��{>�W�[�S(<����� =ƍ0 m0z �����L&���7'��m�s�^{KU ��t �`� �_�޲���Vk�3��i۳�Z ����F�`0�Q�l��u;}x��? �1��u��G 0 Ԏ�o�2���W���o�� =�1������s :���f$�����O	t =C��9���  J����F���c'w =E��9u6�  ��,N�@�Yo�%o~ӛ>y� @� zJ���ah `����jy���Z����|}�@��	@O�u� Hͦo��cc�� �@Ϩc�8Z ������u��o�_��M��� ]F��6� đnf2)�֢��/�t ]G���c� ��(T�@��& �:��P�9 @-u
�а,S�i�CCe��o�K����>- �E:��P	  ��3!�M��	Èo���?%�t��'�� X�fU��D'��̓ ��@�uLo �����ad贛���l����u�����( �%:��k�= <�n��;N`4��%~�F�.!�t�ڱW  XC���]�� ]D��*�S/�� �S�ܣ(���GD6;�S ��t ]��p ��Q��8v(�Y̼�W��\s}S �t ]��S/  ��ya�M��R�E��>~�7 ]@��*�	t ��xܚm/�Jt ]B�蚕ctX 82�[K���	 t	��k|�8 <� �@�5
��� @�� ���� �c�m��P�y��v箽��� @�� ���� �cQ��E#���T��O�N ��t ]�ζe�9 �X�@���Y~�� ��@���V#"  =�s�Fq��)�+ �:��`�8 ��RŉFR�� @� �B�)�  =����Ϗ׭� ��@��m� ��ʲ(Kt��չg�|����' �Kͺ2}�u=����']sͭw t��+�� p�ԋ��>}�E՗�:��"�t�� ��P/���ݼX ��t ��9 `����Q�. �a:��c �^���0�Ƙ @�� :.$� �E��Ķ�� @�� :. �.���kY�� @�� :." �.����R F�  @;����#�t\|��: `]t��aY,��y:���m ��2��@�q:   ��ۋ��E��<@ǅah��  �t �@�   �`Y� @�� �!�e�a����C��
 ���3L3�e E�^A�:�n �t�ډw��۶�	���Ʉ˂�C����� �t����M���m @wGt@:�n�& �.:�AD��C��ZL �Z��C�@7���t �( `���`� :��, �	�g��C��8�v� �O�c� �t !� X� �����t �@���&�b�" `=|�w@��>� X��
tF�t���<Ϗ=%  �8�)b �@�q�0M �.Aj茠�@ǱI `=|�{T ��o~ :�i� ��C�D3���@Wx�8�#�  p�f��ft �@��
ϋR�c� �c�{T �o~ �����lV� ���M_�{TF�t�V�� ����- pl��kU�:�n!�tE�峓; ���@,�X�"��#�t���=�4M	 ��h�h�@�-:��QŹ��  �"�Y��z(���@�4�a�� 8�z���)���7@ ]�t9CC �httF�t�V� ����ˊ�L{)�  p�VK�H���:�n"�t����<I�R�  S�{�hF�n
 �B��F#pS)�@ <N��A��F��Z��b: �H�R(�q��t ]�h�L֡ �����t����N���i�.  R�yi����猦�@�U*�8�] ��J���� ��@�u�J�w�� hS'|x��U� z�@�uLs �U�z��J��@O0� �J����t =���OL� l�f���v�t �@��	5ͽш2Ls��V������1k ��@�3�r+�4w l�r#��Q�:���T���x�2�( ����Ì�ڕ/���
���*?74d- `�,/7��F�����J��;4T �`�}�k��%�a�@/� zJMmd�8 <���� z�@�sj�c:�&�`�,/׵���� z�@�s�j����cۑ' ��W��� ��a�:��{�Y�: -,-5�nQ  }�T�kw���:�^#�h�\�;##�m�� �o�ja����[�}��&C� :�@��r�ˏ�:K �[KKu�VS�hz�Eڽ� �� �Q*�R��#�iF�  �N�ft=?���a��w �G�Іڀgy��qJ �;KK-�V;���
���<�V��j����iQ( ���lF�F����r<#�o�s	@�� ��Fї�ZC�E����Xϋ���9܊ H� :�@����j�P�\t ���s]GϏoz�
t��Q t�@K���-�E $Z���X�r���=_��Ec G��R�ڰ�M7�FC  ����|?�r��=W|�i
 t�@[����9 *�*ki���F��1k�e�#�hK����-�rfU  �S,6���:Z��.ˮ t�@k�l6;\��5 H�VK�r��;z�AzZ ��t Z��XXhOL�E $��|� �:�@I�B ��t �S#0�B��  !J%oH-S�87���Yg���
 t� �檅;
���=  my�8�n��w���4�� �0@"x�o����QgI  ښ���1܉MmW��f���zOM ��t ���TM���D�E Z^
�FK˩�ʉ��+�F�% �:�D���mߞ�7�sx ��ھ�XɈ�N4���5 ]A�H�V�3��<���ft�ڮ6�;����� �@⨩���p6�1X (��~�ھ*
� �@"�Ζ�;w7M3
 �3�z�Q/���������V�?& �:�D
�Pff��۶e� �A ��\%/���y��	����o
 t� ��t�R)5<<l� �u���� 76<�A*�7:z^��UD� �@�-.V܉��=����� �-��?\�576<�A�nU�5�� @�� -����r٬�j�� �q�z�U/���6:�}���A��!�$���Ţ����s��R�h|�% ��Q���,k��\��otj�Ej���� ��@�X�3&�ܙ��a���a�YX����� �b��TFt=�\Qa�Y���Hk߾��H �Kt �52�tu#����f*��� ����P  �jv�>�y����)��J�6uP�� �B�H$�J��Г��V˴��K�j��JaX�w� fq�5R�77��Zm���U��� ]D�H�����������.ɗ����N��-/�R���m��v%����! �E:��1KFF����L���
/�*�OT�� ���V���B9#���8W�ձ���7�B ��t �S(<Il�p�9���X6�}AT�~�*t X�f3J��.�Ds*�7sj�R�o}P�^�n"�$���E���EQdx��\>���R���  �[�%����C�9��\]����� @�� %�=E\w긇I��k��YC�|U*_j
 ���Y�?\��85e�ם�
;?�? t� QFF.^��FE��Gz�T��kK  G˴���Gt�s�q��'_���� ��@��Ըd�������}�0�:���Z�D: ��==]��@�ΕN�;_�h����w ��@�j����ݘ�y�m?-���T�����`���������y�֝+jz{�1� =@�H��J�pކߏI���H�J hS#�.'b�S��W�J'_��	 � � ���&��lʍ��t���u��2����8Wl�������az;�^!�h�0�8�/����"}y���� �ڭ}z�<B��+
Ñk z�@�����㛲ܦ�<A`�H/2u�0�߮ 6���ڭ=IqީM�V�J'�����!�hΐ���:��Ez�P�6L� @��,%�(5��;��U�����w z�@�5���ю�����j:���e�� @�ף���r>)q����j4����^��"� ���<�$~R�m�$2�c�'��H�5m�� ���rPXX(g$!:�c�Z������%om ����VF>N|�x������lݪ"����r����Y�q,�I�W�8��<-	��ӛ­
CC�-o �1@ǭ�~��锕���H�t�/�x�W*�T6�6\�i	 $\���XXh���uG��q�,-�Xz�k?�e�#�t����}��~����25���Gz��p|?0s�4�$V��Lu��hu~�&�f�+�ک��|O ��t ]��^.�$��l�֭����Ho�<+�tuV:ǰH�3���塤����q�h��SN9�M" �5@W���*�7beM�?�פ����O��{�TͰ�;�$�V���\9����Wu����g��%/y+������V�n<�%?|�l���8�S��[��=�M{�K��R�^\���0��s�w�fs�n M� �n�"�^�?��ɶm��,+��:�.=B3�uY�@;a(��l}�^o&j��ҋ8W����W�|� �&t =�y���<��-�}��D�3��f��^���g�i���q ����(=;[)$m��ҫ8C;j4v� ���g6+�[��8�đ���u�:~��Q*U2�|��y� z-i盯ի8W�����W�� �� zj�"��+��CnOw�dvt�nO���)�)� zA�6;[M�v��q���j;� �������8>�-q�D�lyA44t~W��Ԕw��Քwvy�5�F���.��K��^ƹ��p��W^y� �!�hc3�I�"_ff>���G�㿣n ;~��bc�w �{4���ᥥjJ��qE����� �nt ZٌH�o��X�S<oI��^���W�]�=/�r9��|&sX��Z-qgg+C��'n#8euIS�-,�zpϞ�>+ ������lN��5����,۶�,��|Wnh=�3���,�� 6�5/���b�����W��A`G��{D� �Q�S��� �����F�!y��e�֗E��I]uR�魖o�r�&Ǳ8Q�g�33�Ď�+�Ĺ2?�O^��[�, �)=�[�X��~�h����~����v46�̮����o���M�^�0j�������^k63A&s� 4F�К��S�/j4}#�(���;ڛ�m��ҭu�
�� ֣Ւ��\��jy�5W��o�XX���{��� ��t �S7x*�7zV�R.�$�����[/�R�Ѯ����n�ɤ87���X�bs�\�;�p��y�<�ܵ�i,� :#�$��F5�����͙��tu^z�pnWG����l���\�s� �aaa��I��k���#YZzʻ���ߺ�Wy��t ��雱�{6ez�SR��ML����ݵ���c7*�Z�q;�u��0ut��|��lz�7� �6�[�X�Uܿ���( � �}�cP7��5*A�j�u����ј��[_�Rc]�QG��J^&�I��� #��t���Z⧳+:m����Q�t���
 $� �\wL&'_,���(���7����i�������D##u}^f�ް��w����F�i �!�iz	���0�� �/���֛�57w�׮��ß H@bY�kl���hq񛲰���N�'*���F�_�Z�u45�b��\WC}u�{|��c�u��:�+RC2P� �JN��	rq�g}?�k����|���d}��g�"�$ �:�D�o���gK:�=:x����Z��r�����E���]�������X������@�5�Q:�|?�3_��|�L��%�ʅW���l Yt }!�;�ص�8��A��7����*?|����D[�� �	Mw�T�O_Z�2��Rǲšn��\X`����ZX�j��~��7@���k�Ξ�ý{o�� @�� �F*5G��hz�������J��8����ߏ���z2L�l��ǲ�RN�ͦ[������)�J��w�Y:Oi_U���\����� @��� ��0lc۶K.wZ4;�y	��-Q���<�	zJ41�����+��g�W�P���a����Uah���oٿ��* 	�w?@ @:��dN������o��-/�H��_���󢡡�{v���L}����/.���j�/㮝0�}���y?ۿ���S  ���	 (�3d���g���w⛶/Kzjm���g���hr����?ܳP_���B=�N�L�`D�*3���axV~n���(J?J�U��d��Ӟ�4�� ��@���.K:�#:x�S�y�~���/�V�OFG���=+�3�^�z�q�0�I�,��ث ��i:Eg����m��c��H�X,�)�BE����}'�V/��g?��u�K�w^ ؀Lf�q�)�Gss��Q�(un�����X��LN�^��������=�Җe���9����1�L�5~~A����,���w�0���/��d�=�����S��ۯ<$���o}l�ޛ>+ �p:��a��15���͞��~���F5������B��&r�]�i�A�>G�0'��$e����_�������);��+ƩN�e��_�CC����}��f��鶤�����?�{?�j�>���� �A���F6{J47�%)��ql�g-�r��T~ٞ�>:�L1M���E�E[SQ�m<�}�E��5��o�a�M�cR#ȧf㼬al��n=�gם4v����|�}TcR$q�\�Ն���SK� ��@0�,�5�n}��MOnSF�V����?���߉����kे�P�VK��3d���������փ��_�X?�
j��FZ��	+��ʛ�Y)��	תi��/--m�����_�����Qs%�hq�^�U� ���� �$���^�>?������M�����LOR��m21����O_�Q�q�Tj��N���_I�~w������&o�}�0�8����a����'~�j��g���G�ӟڔ%5�-�����.��e�}� }�@0����-[�/��Y���Vk~S�o�q��>=�?+WH�j�a|��g�I.w�����Z����
0gg|���a��
C���\��Ν�"��]���� I���������
 � �dv���?ZX�S�ٞ��q�T*?k�64��hl�9=�Hn���w���c�%��c���e|��,WG���a�geE�JG�p�(�§�m獓Nz͡���^}m���*̓r��єJ[�Ap��"_ �7: �a�11��dx����l��O6��FQ�T�@��*##F��ϊo�3��%��꾯���,�ԩq���x�M;�}�(@r��>=-rFFd�E���գ�\wk4;�������J������s�� }�@�#p���}�K�Z}J|3��M���F��o�w��(�.�o�Ӣ5^č�s$�9/��v�7���[G�0\ò�p�LmwD,m^+�1\w�}[����?�_�\	'*���q��H �O� �r�Sڛ�--}O���ksSޯz?��_����đ��C����9��:?���ď����p���'�g�/�,�GʣhgZd��F�#MWi�RƎ{�8б���e:����y������ �� �`�1:z����D�����g���7ڡ>4�Qg��v^t�2�>־���AԈ�v0��ټ�=��#��Ȯ��N7�&앓
��D��=R,~�cq���ُdz��o���W �9 ����~�I,�����ܗ���7�}���*�������#�3,�Z�	>%jͺm�{$A�b��8��-�=�:��3W\wg�;�k��d��0���凄a3R_��8�N��O���ZX8}zϞ~� �  �`�2��Ʈ]��Z�M�_��tv�޷Z����S#�q��s��Dg*�[������5����{,���`"��yӛr�<�m�Ɨ���k*��
�;���:�\�(W���|M7~��ȟ��\]�3��Q���Ү]�:]�N�A@��r�������gr�S�l��hy�'2?������-��n_�̎���l��D܀�q9���T���ǯ�Z�C~.��3��M:���4s��Ͷ�s}��Q�n�2���YF�j-F�65jީ���[g�X��[j�Կ?��Ͼ�)9 ���J��4ﾑ�������~�ڙ9*��>?}�6�[U�?_/��E����Y���H�L�W�V�ݶ��ڶ��h�3�����}q�OQ��m�G��e�jF���r�sG�Q�UQ�V�U{L�v�t�c��0W���V��ԧ_q�u�s� $��㮼���7�|Ź���^(��u��&������<5ZXP��}�G��T������;dh�8�/��$Q��_��gL]Ӽ J���0�(����8������*�:q��ş�*�'������6 \�䌒�
�V����������MQA�:������ࡇ.|��^w�� ��+��y߃7ݴ�9���������cYYc˖ߕ���D��w�g�o���Z�Z,�������GF�&��)�M��̈���PW�0�ϻ��f3��y�0f[�7��� +D{��v!���A9~Nďc�߹)����'w�fs���[���M�:_kP�\��tX.?g��^w� �oo��g��|����R���?�����jx��ϕ�ы:�j�z�����F�ը�:�Ͷ��� 7��<C�I���W�4���G{�P��5}_E�\�Q������R!>ҾLs"~�����W�<ٯ���ru�b��i4��5Ha���MO?�͗]v�G ������#���z[:]��HWVC}d�鑚�ډPW<oI�"��_�\��8ԟ*���kTWF���_Ċ+e*���v��R*�U���p/������]}1d#�ΰ�B|ǟ[�q8�k�=2E�#1��<�OVF�$��O::Z�Z�+*�gg��_.��#� `:���#�����WLL|��3���tŶ��F�/�T��M�:q�RR���}��Ņ��q��/�Ը��G�]���?���I�8h"۶"�5CèaX
D��Ȓ�y�H�m��R$�J�0n����W�F�е�Qdɣg���_��ըR�[����<N�h1������˽{?�? ��'���S*�''����0��ʲ�q�����?;Z^�'Z\���juf�b�/K�����Noo�����c�~��݉Ʃi���S�nY�8����d5���o� �yO��Z�">J}9ov|���?��+�w�ǿ���g�!n��8��ǌ��Jڮ�'"��Z�e{��V�u{)I�®�Gsh��?�q��  ���o��K'&��f׭ԐQJ����U���=��V����yj����y�j�{�p��rg�1��Aqh�]�$h�=?d��Q��q���Nݎ�Fh�8�[�G�f�Fߣ��a=~_�8���q�ף�����7'�҆eL�U����~��~�����Z�0��j�H�ϣ�O$��Hg�F���{:>�}��h� ����n87��o޻�CLk�Ct =�o߭��w��ǿ~[&S������3�W�1-���jGB�F��y�˩�S���'��~Z
��#AmPw(\��R���x*�V�^�������㞏��y���Rq�-Q�M�^{�~e�>�����Z�������`+g޻���oS�C���<�1n�~����Tl�������7+�D=�������>ծ��*�Ո� �<7��}����л ������&�����ߛ����ܲ#*��*۷�4�q�)�-��?��:�U*W�����c������AY?Q*�U������!jBH����P^�#����G�{�F�7��Q>��ˏD����s߸���s 8�@W^y�7�x�s��ί��Ł�C�u���俏#������NW�(o�|w�R#���)q��՞oY�J���~ԺruA��� �/?�V+��>����?t�  �@��}�|���sa}绅�|��dv�Ԇ^j���Z�QG<�J��診�F��oJ:��=������ ���J���}ҋ����x�ڰW,>�%�]v�� 8"�V����{�?O�o�;6����M�69�<QG�ukT]Qk����ۗ�����l��8�O�L�dYY�����6A��~G��ԙ�ҋ��-?�ju����g]~��
 �t ڹ���o�s��z���w16���G�U/���1gRw�畤T�^�R��Ԗ�txue2;�1b���%�"U{��
�n�~$��?�Rig�X<�IW^yˌ  ��@K/z���n{׍7����o����z�TjDl�~�Ȭ#��Ijt�ٜn_�����ը����]��7!�f���#�9T��@�A?"�x�̜�P�z�iW]�� ��@��ھ}_���[���[�|����duZ��z�Z�v�V�bYYI�Oj_�̎�q#�8n+A�`|�[|=$�ּ�b��Z�ľF�|{��~��7 p|t �۽�3/�馗�cr�Ϋ��p�8<փ �����n٫��)�(7ꮻ-J����,+��'$�8�gE�#WW��@�e�Q�~ah���şڻ�_& �u!�$�޽�M7�櫣�w}8�Yfg���BM�WVG�{�+C�����}��J�=�q���ś�M��1�9�yq��/�D�������.����]X�V+��>�_v�G��  ֍@�{�~���y��׾��JAp�֎ ��+���q�Z^�q�-j
|*5�\[�G���K�'����|{W�Vk���y/7t;��(g]���VǚKK��e���1j p�t �r���vo��{GG��۸�^'=c}�E]����W?>�VCg(J�&��ͭ<N�����߿Ԇ�j�6�[��������ڿV��+��o���ӧ��w�啷.
 ��� ��Ko��;�|��sz���ED�	Z'��`�E����U��r��U�G�3?����<���:�ϋM����o����X�j��a���E�����W}�Y"w
 `ct �u饟~��7���'�|�u۷?�2FS7���V�]���ǋ��>��-u^��w�V���8�w���s�ߗϗè��}�Ő�ǵ�u��~,L]� pù�g�}Ϟ��V  ��@�h{��z��߿����?��3��s�q��7�ڨQ�ƺ����(�Y�~$�a�H�>?���n����ee�Gęf�������:�0l�G����v5~��wI_y��w�W�Ö��g�z�����E���[?+ �MC�H��/��7��ڱZ�?:��]g�rg&:�tt��֫���t���E� =���Ê�u�}\�i�=�����N�z%]��l?>���߯�ȹ��㉢�Ʊ��G�o��_��M�zb%�ըv`��o�����V�\�s����#䌒w�z}nq���K��]uխ� �T:��p�U�Qr�-����:���y˖���]��#��ў�`"jm�iV��6�	��	�T4?�Gw���k �:���{����}��ӏ�_��i�]�w��޻�h���)��k��P�N4���������i t���\q�G�Eo��G���������'sW�e���M�v�A�C��s~s�i�{�%���& ��"��%�x��k�̛nz�_�|��ꤓ�c�f���9|�j��m�4u����ʄ�xǥ����|U  �G��k{�~���r��_���ϙ�dvP X�ã���am|32����R�r���w�[ �@�۽����n�q���Κ�bj�����h#��{r0"�|��D��S���|�E"� @w� ƾ}�]u���=3�寜}��#�;E=$�����s<����x�)�w�J��^v�e�C  =A�(W]u�ㇱ[n�}�����ɋ㶰��:�4�U���6�đ)�׾�籣�� @�� ��ݟx�{�{�SFG���s�=k2��I}����#E�ڷ�<���q�G��������\¨9 �@0������⇩�oο�S~�o۶g���P*b�qzx�kD~���H皷Eơ_�8��
��.�̥�~��
 @:���g�ǯ8p�򿞟��g�y��L��t<���K#�Թ����g�d�ޛ�#  �� �����2~������SO��۵��)�.P` �F�:�-,\�7�_~��+r�  �C���}�mo��׾����~�����OL\$�a� +�hi�I?n�����ߺ,  m� p���z�?����==��O�~��c��D:��)OYX^>��W\�
 @{: ť�����a�����c�����/tm{�P��F��/-=����kD�- �d ������������ٟ��g�o��o�^��
C��<gBP�G��Q�J��^��5K!AP
����3�ܶ���9����6�x)*xk��V���*Z_���઼_	y�d����!	��>��~k��7���f�,�?�w���ם�$irrvc˖g}r��W�Z�qv�V#����cﯾ�s���ί�p�	��pቡ�.� 0��z�w<��1�^p�'n �$��V���]qz�UW����x���?��y���i�����~�+��� @K� `ժ+�.NG\v���_���zg�>R���֭G�������}�'�!|= ��:�p��W0N���~�1���|��gwu-��A32�`|���>���=;O���0�:�?�󁋮��w\כ�.}fW�8_��ftt���m���ŋ���Oߞ @�� �$�qz[���W��˖M�~�Q�������۽{�Ķm����%ǽy�Ja��:�4�
�����-��s��>�l��K�
u`�<2��<S�t�p��Xq�d�ޱy���u�~�c©Bx<##���_�{��3��x�Ct��l��oj>��я~�˗�8ꨧ���Z ԁ�ٵk����v���ҕ��3	t�Cd���s�㪫��ޥK���^�3g���\�w�{ǎg|�3���S�� �C	t��jյ�V���喇nZ����=='�︩���(��~ʽ##���Yg}���qi+W�u ��	t�42�$���K­��
K�~7|?��!��������������w�Z��/��  ?�_� 	�����9�{&�G�(��X8�ȧ�bq~ Z��Ȃ��۟�,;�g�� <
���<�
?��3�a������?��(̛wL ZK�Q[�.۶{��8�����r �@H����p�-KÏ~�+}��Ó�</>!�s���ў��[O����Q�:眫�·�;��  �G�$�����w>+�FX��|��8��,+ y^۷�u׮'t���3ϼv2 �~� -��m;~���aɒ��󛏿o��سg�Ķm'�\(,?�mo���� �@	t�466/�s�s��91��	~',^��P,�������ؾ�����sŪU���-`�t��k��{�}��z{o�{X���!�<a�er�v�\�}Ϟ�_��>�W������<3 ��� m��(�m�N�;�w,��� ��a��;�����b�/9�[�?|�[?��!�{ ��E�����Y�ᇟ�w�����6�����< �Jv�Z<�k��GG�{�;���� �P� mnllAx��s��s��`���E��Y��:�y3ʗ��޽��y~ğ�\y�u!|? ��&�:���8��n}^����1Կ,�%��c�O�yޕo�~��ݻ��j�pD�ʕ���N9 3M�t���ly����5�����;����G���z���[��YvC���r���' @B: ab�+l����㮻1�����{k�y�QxZ�ԣ룻w/�q���ŋ���X�=!|# @�: ?'�
?;����_��Gc�����aX���0k֎ ��;�c��-�v-���X�'��|�G�h��4>>'l��zZ���C�����ϟ{��C��'�Li4f�;v�ctt�d����q��׆pG �V$��/##K��|��G�����̹#,X��;b���:Ϟ=s㟿�a׮e{
���>u�ŧ�r�?t ���k>?2r���|3|3���(̝{g��;COϽq�=~����,�⟭��Ν�����Ʊ<�a?��]�r��  mD�0m���{�{G�������1��
�������y�,�Y�_099'��ud���0:z��0��� �St ���yq<=��������J�}�̓����ŭ/�={��<4��kL�w�Fc���G�}d}t����w�1 �s	t �sι��q��O����s�o�i�]]�����vbw��K��yx��ٻ��S�oeͧ*FG{c�/��{���cc ��: 3�7~��q�|j��g>s޲��zvW��W
�O�={��ٳ�ϝ5kWW�	��c|/�{W|Ϟ�c�G󅂋B�w ��	t ����o�;N>5~��N;����My����'vw�8��k{o�ٳf������]1�{�X�����aa|��x�$��.�H �@��}�u��#S��\���<^�h��<�w=��{dy���q�[,�=g�h�qt~�;ݣ���{a��h�aS�E{�8�q 8x: m�S>�+N35է?�����1��,��ƞZ(�>�X;�P�3?��vu��*G�f��S(&
�zL\�FcV��1���������9&&z�M3ʛ_�(: �$�@�y���-N�q����o|���n+��]O˲Ʊ��c˳l��<�X�e�����Y�&fOL4fŹ{r�1��{�899�������'�
�f͚�٭��k͹�k2k4��_�b�h~mt����F��������u6Y(�l2ϋy�=29�5Z(����MN��32r�i�����5�ǻ���K� �� ��1�tҵ#q�yj$iÆGŚ?���y Z�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@ ZN�� �� ��,�W����JeW �6!���T(N��� �	� ��F��� �h# hIY���� h hUϭ�j/-��_ �: в�</�I��: в�,{��������� ��	t hqy�P*�腍y��<�z ��	t hq1��g͚:U�������c Z�@��`��=������y~���f͚{ �(� -����ɳ(t���/����P��y��V%���N�j���rQ�`1�_����� �	t hy�?��}ʆ��q6: �H�@�q~G��:\܇�<�?q饗��=�y�� Z�@����8^hF�����O�rpppw �!���(�n�{7�#����������~ � ���8�9��N�����7o�fw Z�@�60>>~swww�����j����  �� �֭[��Z�ޙe���ω{�'1��-���; @�: �����/���}�z��R�tm �D	t hY�}>�G���h4>^��f��� H�@��qC�8
�_Ҍ�<ϯ�V��J�rU ��t h�r��Z��oq����������zV*�� �� m$���b�
��0���Gb��@J: �������c���j�Z�T*� H�@�6c�1:��Ł������k����r� `�	t h3y�D�OY��1җ�J�u�2 0C: ��y��}|dddC�͞�����K�� 0: ��.�`g�Z�Tp&��z{o�q���W�^�' �!&����Z��838}�i||�s1�O���= �!$���Y���Z����<-��^166�š������� �� Ц&''��P(�a�Eh쇸e�+��>����; � m������j���|u�@](��V���\._ � � �Ʋ,�� П��8�6F�;b�, �A$���Ũ�1����5+�����*��{ $ �����{���N��y�2�9��Z�vloo�y�x �i&��ͭ]�������(�D��}��c6n��{�a`�	t � Y��o�������������O]�v�] ��@�P*�F��j%.�L�_����r���V*�� � :D�O�j����7�Ó�,�r��7���/ x�: t���<���O
L�Eq?��Z��l��  O�@�R.���j���u�i�e��韨���J�� �@�#�oc�_���"Fz1F�_�}=.���  @�@*�����<60����j�Ν;�=88� �: t�/���z���F��/�G��&����������> `	t �P�R���j���L���H/�H?C���: t�J���V��(�<�����7o>���� �8: t�<�� ˲�����v��1w�ƍo^�z��  �A�@��T*�j�ڛc�5��a��v�����1��"�x, h���j��Ƹ�>�Y�������k��3� �* ثR�|1F�fY������������c���6 �@ ~&F��c�?+������zFoo�X����< �#t ���ܹ�#�<-p0�]�׷���  � ����|��Z���e���%���=�Z�r��� �t ��4��^��_���?��g���V�[�^�U � ��_�T*m:�X,~9^86����w] ��	t �W���'�
�B3җ�U�e�8��V��S�T�5 ��: ����~T��^���bL�n����%�\�/�� @�� ��*���644�?���?��E��tbb�_|�o�[�nk �#	t `����{xx��B�p}��L�,˞����77n<y���{ G� ����﫵Z��q�� ������} �o t� �r�|����k�,�\=�i���j����J����"�������������3"���thh����/ :�@ H�R�b�x���;��&�gw�P��V���\.� � 8`1ҿ#�1�?�rI`���|R���^:88�; ��: ��4�`����h4nhFe`���|^ooo��g ڞ@ ��R�t����oM��~L`:��Z�~�R�|8 ��: 0-���C�Y�5�IF`��=�4<<������ �-� L�J�r{�^?��h4��~R`�̉�y�����|�}	t `Z�J�-�j�丼6���E�{{{/��s mI� ӮR���ݞ���cX�-0]~�V��s�\�X ��t ����2F�Ob��L�<��?<<����� ڊ@ ��8��V�����Y�	�[� ����暗�X�b2 �6: pЕ���z}k���Qa���Ľ���oO�����/H ��(�JWV�խq��,�����ذa��֬Yss �-t ���T*���뿓������X�e��ƕ�7o~�y�7 hy 8�J���6l��[1.�.^>9�D<ǎ�8�e ��	t ��k>�=44tR�XlF�s,�����gJ��M��&�����ϦM�^6::��xyj��4uo�|o``��So��E	t `�\p�;������M��]������3� �,� ̨�����V�}�Y�.n��j�z]�R�I �%	t  	�8+�yxV`��@_�n(.� �$� $c��������<,���^�ׯ���O��#���T*�/lذ᥍F�����>k~< ��M�7o~���Z�@ ��<��^���<+=6��gm۶��8_ h) HR�T�{�ƍ/�6^��g�B�/���/�� -C� �Z�z�����S{zz6eYv^`_>11�.����!���N��]�j��8_��}���q��_�Tn �� ���C18�k��;�x����q�
 �� ���W��S�7��>�>44tI�� �� @K����|�^e���c�<�B�X�8Χ �'���S*��~�%��lbb�,˖�ɵZ�r�|c  i hI^x��b��t*ҟ���<o������	t �e�H�mxx�e1Я���xTq^W��^P.�� H�@ ZZ__�}_|�+���>C�ŁG5u�� �� @�[�n�֡����B3�_�%q_޸aÆ׬Yss  I h���;b��6F��b���E����?����$	t �m4#}�ƍ�����,��[֯_߷v�ڻ �� @[Y�z�������j�8���X,�� �� @�Y�v����|�e/
<һ6n���W�� H�@ ��T�����uC�|a`�,ˎo���c��t �m5#�^��:��������A�$G� m�T*mٸq��ccc_β�遦�lذ�7֬Y�� @2: ��V�^�@�^?5����#arr�8	t��t �#�J���P(�K�\:\�e+�=888 H�@ :F__����76����:;t�E===���3�$t ���J��V�g��zIZ!t�3�@H�@ :N�R�D���Y�����������6�v �q �H1��_�Վ��R�\s������� ��� @�ڱcG_oo��婡s�-t�$t �c6����V,o���(˲�޴iS�\�3 0�: �����wT��7���c�.	�g����o/��q �x�J��Z��2.?:���	`�	t ��\.__�V�,˲��a���� ���  Sv����===/��zJ�,�=�����#� �4_�q��U���߉�G��eY�1w�0�: �#�^���Z�vV����h�B�(
��ӥ�#� ~A�\��Z��?.�"�� f�@ x;w�����}e\>#t�,ˎZ�~�1k׮�+ 0#: ���=<<���_�G����$�f�@ �����R��>��`*�? � �1dY��h4��#B��9t��%� C�T�R���g\~0��,˞ �1 �q{챗�~��kb�>3��E�z}q�J 9� �8V�X1Y�V���m.����$�f�@ ��r��z��..��X�e���[�CN� ��y�Z��+C�����  �h֬Y׌�������`�t �}�z��=�j���,�6�:���  �!˲�Cz�� f�@ ��R�;�z���\��� ���  �����Z����<=�'�0C: �~���_c��e�ǟ�7 0#:���������-����
����	��t�"�f�ڵk����h9Y��m�ǟm��͛��;�� �!%� �S�\�1N١�}7m�Գcǎ����{�1� ��@ h\p��C���[�. p�	t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H��,�ST�J��    IEND�B`�PK
     t$v[񐼛�  �  /   images/a4af1710-95e2-4b5e-9600-8e4d90487313.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  ~IDATx��	��yǿ�������=uK @� !a#d!@0�A�B)8��VJ>��*�\I��8���l�vbLى�KBh.��B�J{��5GOOw�|_���JZI���z�UO�3����~�]�_?�P�T��L5 ��D2ՀH��T"�j@$S�d��L5 ��D2ՀH��T"�j@$S�d��L5 �iB پ�2H�{��LP�2p�c�����Bpp]>�p̘��a����D��@�o_uu��8hZ�"J���VnA����؊�w���3�2�X�s�i%�~��6�駿A�y�K!��-�%���L��B|
-�"���"�qS������f��wu��ἁ�e�6�4Ͷ���|��9s^�%�}���Νg�%�	Ӧ�AG��+�W��Z�o� �x��(�9��A���T|����s;�j����ѳ��;Rp�ٯ���Ȼ�^	���<�A��-�3�؁�B`6��Qv!*�q>
c�!���JV#��_|�s?��gESSƙO�K��)r ۷_�0���.j�͛�QU��V[	[y|{rAQNSUu��8�ʮ���ZF03s�_�����M����لy!̚�dR�@v�x���(��d[��`�t=�e�N|6��	Q��ؠ�yY�q����-9��9h-W���O�S��ݽ�;�޽ �g�%2 [�^�������#U��Pa�p�8�8�+�
��qިp��u}fd��Pt�m��Z����//X��RK�.t_��}ɑ�E���ï�E�H&�,e��뗛��Vɶ�\bL;����6��+EM�0��4�=�`,���3p?/crэ�x� ��;;�ܜHbvw̟�"D�H�P@u]��,���EW�Gh�C�/���r��z=��En�P��޳������k��&c&#kӴO �$����8YK
��A�)���@*�2(t �7_��NrS��'o@�qeP�1�aV�Z�G�X��gr����hR}���u��XlU���}����X�A�������[[������H�B2u�A(���J3��߄�������Q�d���U�ڄe�:'DA;�3���\w�cY��c������X�qނVGY��1E���\�׺^z��"D�Ё���X��rY_��8|W�뚪��ef�����&"/ƛy�]��U��+|!���,!y_+�b���v���ܹ *�
d׮�`�ѝS�U�A���1V�����MU��V.��eۯ����*h������y�S�<]�o@0��~�R����#W�ͻ;a
���|�|����0HT��V����Qձ�o%7���z���Ӆ*�b1�<s'������ �h*����(_�2�0U����x"+9wڴ���T��u֫�B�q㵠��p�-?��?�c�W|;�(�2�����p�����S,��8Z�%�{oN�r�Rh@����t��B0rk��U�l���h[l���]~dB�%.0�d���B�˥�LB�s`��,�����J��l�:���D.��l�%�	G"Rh@��tY.i>|A�a�燺+�̩�x?!�5�F����8��(��y��Lm�J�&wD���-�;D�G�bPu�&:��� D�Ѐ`%�� whCB��-��m���H�
�U��q��"$�OF�X�R�uM����/�)t�C�>ڠ�ԥB5�G�7��y��J�R�0n�$��B ,�1���*;�s��t"��5�9���~'U,z��0w�L�@�����eٱ����͖�d�4�TJͩX�����aR:�@� a���P(�����IU'�q���թ��f=C�9��BI��u|�T6�U8����Oa��n���2c`�M��5U�KfIdX'�[�4ya�P������x&c7��d@N\�bDk�ރV�<��gvw�-��{�	�I�Þ:��RU�_�*]c�� M
 ��4ݾb��D��\�d���M������q�?��u�R,*��6G`&4�A��(�LnK�-KI�㄄A��@D,������𣆖�F��o
�!Y�9��?��z#��{�:��C���4Q����q�ױ����-5�4�C#��)�rف��|�r�[��ϱ#����U�s�0���=aXՁC��:�/z�h߅֣a��XVY��I]�Y��O��{�麳m������K��;� LE�ajj�B�13�F��i���y�q�O�>�4t�[���b�׻.�����00P�S��MP(?�����O��а�V$@�3�R(xj,c
~L������nC_@�2�+j�;hG3	����o\q���=��"X��mK!_1�'�	�B��2���ɶN���t�Z�w���ϭV�	��xB����#�x��r�)�ሠ�����H�1gͮ]6mڇe�lh�*�W^�K����	�Nj>T�yaa9t� �Es�l_Ƙ��|!�uW87��
��ŋ�\�.�U��R=62��+T���wnF �Gh@ǃ�� ���t��O���Ӕ�:���nMG�a(4 �a�2��pP�����ňdh���e�<���&�ЀX��� ���î�QG(
ǂD8�)X��x'p�[�F뺗��X�x�a�!q��7�Ԁn�K��d��`�Z��qu�)�A'1Q)ڎo	�q�sJ$��kF����;�]]eN����A���[h)�uuZ��zc����#��P:�� L�>	�'��!���DB��*Yg�X�=����Z�3��p�#Դ���.,��Z��h���@�4X�U���4<���� ���%��ٶ��aJ���R"3e��10P21�Ы�K�:�P�:��{閖p�;���jc�O�!��xl�U�Y����l4?��؞���Pu�O��$�������)ɨ�w<䪀ww�i�^5v(J���|���A��[�&4 �L�����2���
v�f�:xag]d4#���PO�|8�sjX�����/x��<��=��
�������٧��t�O���r��;&���ahNXP��K%W��Χ,�C�Ac���tzώ����/� a)T�5mZA(T�A6�-�WL�r5+F��*�i�X4V��+;R�P�,��I�QR��-&���0dZǿLGk��ܐ�E0u]k���={��+Y2y��8�b��`��6QQ]]��Ȣ�?�k��8��!A���e�qi%!�Nĺ����:�ʨ�P�&yW��>h���hIYϣB�}K!a��0u!<���55]==�����
ӜMM���9��9u�rm�u? �����q^���V����/km�ST����91��6M3����Tz]h�kcD��<O�488�[�������jU�3OB~7����8�x�~B��,�:]�����ŦC:�����0����s�0%=�
��83H˿
Z�CGG	�!h��X��L�0EiLc< ���T{���d��|W�w�ˉ���"�s	�<I��mхB�<s׷w�n��e_�����/ףK�@o�����4����\l��aL�Tu�F�Ș�>'DY룐kS��i�[���׵��W,����}aY��BP*����C��a\���>E	�&��_B�
Hw�g���%صk,X��o���ݮ[�vr�\u,�1hl\��vh���13{;1.T�l#��LU���7!�$A����M���D/%�<.HeU�O��ê��>W*�Q�s�10p�|�z�B�Y��qX��o1N��6=	�}��\.�9�HU�e�5������iY���ta'�ҲB����*cP~SUrI�A���E�"���.m���^����$���|t���e�~������w���߁�[���SO��%7���t�������>� �v�G�
VB���������ןd��|��֗!JE21�����fϞW_�WUc�f�������`)�ĹEř��򉏬��4<cX�l�v]�Q��l��6����֊�U�BԊl�ڪU���/��Ex�|��g�ԺU�	���J�Ĵs7f]�cs��`�����K�G �h�s���w����L�v���oAE>u����x ;�@�O��1�τ\n6�(c���@��#S�l��^���,�pO��RQ�s��f,�@Lb���j�f!�϶��mI$��[���o��s_��g�M7m����c)r c��+�odع41�t��W3f��]�������2�����t�칡�����x�7�9�jP�`�0��'�5̈́�k�|�6�QRV��4-�wt\�.� ƞ<ZM�͍޿�,�Vp|�R$VaR�"'u�u#��=Id�n��χ���_����>yM( 	��L��2?�S&w�=���,@F��#E�g�-ؾKO&����+�.lc-I}�_��e��͈4"I��9clB.�)�g�'���i�Y�dӄ2�j��ݎm�����	�����^f�ȧ	$����YЁ�nl�Ñ��	�!����ׄ�v�Z�c+��;�=v���6Zm�R6(�:t��!��BP�����;h]�^�C��
���A`���؜�#�.�6(��L �C�����a�9���Q��=�nV�T@H��/��
���c�/c{f��~���{!jM: �C�������/J�Wb{Z+�ȑ�я{��!P����؞cS���A��nS�z�4�5��sB�%���n�h_�??��J�
�u� �$�J�?��c9PHo��VU(,��x����'��S!)���ߧ�sBX7��� r�k�{�kx�h�HMê�L5 ��D2ՀH��T"�j@$S�d��L5 ��D2ՀH��T"�j@$��'FS��+"    IEND�B`�PK
     t$v[��r�  �  /   images/022fab5a-d187-48c2-96d7-20ad2a5d1671.png�PNG

   IHDR  �   �   
VS
   	pHYs  \F  \F�CA  cIDATx���ylTe��񧥅��E��Ũ�W��+"����K��Ƹ�5�ܪx}��z�AM4z5��B"�DAcQ$���EEJY
]�=�c��t�zf�s�sf��$��az�<g&�g/3���m�q����S (o~(o2Q��P�dJry#	`  �9  `   � p�  �  `   � p�  �  `   � p�  ��D�y��)))�WSS��$Pmm턖��;l��&���&�M�D���N�~L�.�Z������{a֬YM.��̙3K���/�~��w;�{^֎My)o�(/��WW+o�iFx�d��ի�޷�'�����1c��8��w�*�ż���ƻ��(/���-��ZS(�r�w��֭�yߺ���s��_�<����nhh��w�[��7񢼔�*�+�[���l���-ee�����������y�i�̆��ݻ������:��۷�xo(�奼aQ^w(oq����n�y�������{��޽{�BTZZj?�p3d��e��z�j+�9r�8p�IZ�奼����@y����җ�2}�(� N�1h� kǳy�(P�p(o�P�p(oaڵk�)S5����y�  ]ASS��|^������6u  �={�e�?�����   �Ai~ ��4.�Nm  �LY����DWTT  5?+s�u��#�
��~��q48̅7�|3����Fy�Ay;Gy�Cy�᪼��ωn`�ۢ&�B����㓆��}|�P^��O�k��Qk7��m����t���   �T9M�B���j�0  �i�t�~�>}�  `W����V�(��  H2�f��JZՂ+++�Z� �bSWW�u_V k0V��b  I��Uښ p�  �  `   � p�  �  `   � p�  �  `   � p�  �  `   � p�  �  `   � p�  �  `   � p�  �  
2�{��m�8��k�.�z�js��g���#�4Ç7��S__o6n�h֭[gZZZr����sꩧ�ϧ���ذ{�n��n߾=���ٳ�5j�0`@��777�m۶��>���ٳ'�c8п.zN�ijj2[�l1�6m�@�
.����o}�Qs�A��^�b�y���<�1cƘ3f�nݺY;�����ܹs�o������z���s�5��ݻ��y���� t���7����O=��Y�lYNw�'�9s��ݻ��wk֬1�?��ٰa���\ O�8�5|e�ر~��~���\v�eV�W�?�x?�o��6����>}�D��@�2e�����x})��RUUen��v��\Bx���9���v�ifĈ��3˗/7 ���}�f�ׯ_?'U��!�b������z|{��&]ߠ�l�n���\�2pst��R^^n�O�n���̧�~j ����$y���=��c���_F��p�|��G���/7Gq��c�&|�)���A,]�Ԍ9�TVV�}�iӦ���o4 t� aժU��o4Æ�W]uUƠ%4�158(�Kε�T���͵�^k��~?�|*C���ǏϸOc ��5�馛�Ar=z����r�-�ٱc�Y�h�ߕp��G�	&dbSw���� �� I#fm���袋�F+0�y�f��[o��w|p� ����&���6�s�Q���^�߶`�lӯ�֭[�ԩS3� ~���Q� `KV �����d�s�f�{��[!�p�B �d��j����4�TMwQ�qI���臰�}ӥj��{ 6d%kj� U릦;-4���E��z�7��W�]�����` ��� N�fi-Ƞ�BXF1��j������3��K���Ԃؐs�}����� 3PH*�R-��Cm�O��K/��,X�� @Xyu��i�v�ի}�	���c�����W��4�K�ඣ�'M�d^}�Uj� B���k�D-t���HmV����;��ˍv�a�����|�� �a��ڰ�X�.��aK{�8�0I>t�_|�_�;��_쯂��= �+#���/E��;w��W?b�V��u���j�z��I�x\y����)��=�u� ȇ��[�4�X��tŚ���w��v$L?������/���J�5��P��y�gN>����~�q�{Z�]-��N+t� °>z*ª	w�>����W\�1b6,�4�t����~��6Asݵ���c}1�={v^���i�^--�?��_SZ�&E{����� �+���
���>�b�����m�ڵ9=^s�/^��Z�v k S�������~ڸ�k��?�c�=��>M������ @>"�?���T�U�:묳"	_}�)���amذ����O��p[���2XM��Ԉ�0�RT��u��ĉ�S������3��O>1�ƍu�#F��$����ƅA�e��\` ad$�6`H��X5��a��۷�)F������݆O}�6m2˗/���-&���m�Gp�Z�9���c:홬�����СC�j�ڶ��Z1 �a�T��ԇ�>�4�(� V�h��F�����y衇�}���-(r�3gNF`+��;�8���_�8]p�Y�}��� ��6��Q_��4���)�MJJX��|��W��DZ{9ݐ!Cb`�lo���)H �
�9��Ԡ*M�� �\�֎�w�,��͛7g��{H��m�0���o�5 FΣ�R�aM�E��Z0���կ��d���/ +��ɪkQ�\jª+���/ũ�����oV�Ze  ����&�2��� F!д#-7ٖj�6��@�	��9�A��h�F
�Y��ꫯ��ib�~`K�240K��V�s1���§���sN���-b�g ք`�fUS�O+���:ujV+�ւ^�r� [�������<b .Gy�;vl�������&+��BЭ��T�>��k�k��H�����j�+V ���.	
Ԡ5�<}���i�_~1.4�|�M��P��y�P�C�F+==�����qҨ_�)֘1c��ɓM�~�B���*�\^g��h*љg��a�����5�����q��y���6��y���Y�z��������>}��8ai������{���E���Ԅ^�⨣�2w�}wd#�7n���Z�R�ng�ٺu�rZ� ����|p'�6Q]]�o��f��OŜt�I�5�k��a�:|��硫U�j}�\Z(��|�n�G1�~D�I 'u!��5�3	��p�ש���j�6�Ɩ-[�ܹss�&Z����O��|z<���y 
�8I�Q���~_���۝>��_�ޯy�I�~�s�4i��ի��v���%K�>�j�꿞2eJ�}��z=�����s��K/���5�_:�3zOn۶�����fٲe���q�;�k�`}H����Aj�:G�ӑ�x�	���]w�)&
`��R`��Q���~� @Ym�f�#  ��  �p{�';B  �:��"� ]�� ���A� ����fAk�
_ ��Y	������%| �������~<�  `!�{����	`  B��7���� ��w k�sG{�v��/  �+���m���"� �S������τ/  	�
\mX�K�o
�_  2�m +xU��\�|w;R�2� ����
Z��U�7�6�����d  �_2X���]--iko���F  2e�B7�>ގ(|iz  [F �\(C��� �}l+0�4= �1�5`����  ��Y`j�  c-��|M� L�>`�r�<_\ \�B
Ԡs�S�l��   ��
`����LjmgV�  ?�ր;�jnf�  ��n��T��� ��vk���W�g誆��}����'��� (Y���D郰����ҥ״������iLZ�Z;4�]5  I�����U�TM���>��a=N7m�� .--5  "g��ٳ'�)LZ�R_���a @Ar�
�ݻw��[N���� ��X������]�c)���  *��}�����ci WEE� �P��QmU� ��,�� �"� �r�`�Z0 �P��QnW�c� �B[ ��9�]�R+v1 Pb�8����  Ik8�s� �B[ �4 �_�*��� (�p�H  
E�5`�Ϧ���M;8�� (���jU�~0
qm� ���Vyy��l���jzV� P(b`5����z-X+`�� ($��۪��~`[�B�x�Y PH�t�VVV���MMM���~_ �B�l�RUU��7����/� (TN���VS��Af���G�� PȜ��Q���hm)��m�X�R�c� �$&����
aV� ��p[/ ��%6� (f0  �  8@  �  �0  �  8@  �  �0  d�m��݉  ���O���
��;w�;  ;��A�~�2������  ˴ß�5}׿� ���7  �>Ur;�{�  `��gϞ��n���f�? �}j�VStj��� �Y��ݻ���466��x[M蕕�9=�����y)o�(o~(o�(o~�Zy���G݊�
��� ���{�}�jjj�g��٦P��P�d���������������  DL-�ܒ��?X�_�  ���U-�G�0�� �GF 3� �x�f���Wâ @�����b���0_|��]��>��$O"��M��-L��X������矛w�}�lݺ��q,X�/�=n�83j�(k��¢�vP^���#��͕�^58������Q�y�~����.^���(αc��t�R3~�����O�\�xw�7P^�(/���Qy�f�V�,3�{a�~<�=�'g̘�3�sN�6m����y�E��{�����8�My�Gy)oT(o�\�׆�`�~^ZZ�?�v�za֬YN�K��;�x?��9s��VWW_���/�>#�sQ��Q^�k�_��)�콰˼�8ϻ��LBxo0�?�jkk'x���9N�ql��奼����EY�($:��v�I�����y/��>oʛ,�7ʛ,�7y�  +  `   � p�  �  `   � p�  �  `   � p�  ���i��x+��    IEND�B`�PK
     t$v[6ah    /   images/39d025b2-988a-45cd-b457-87e73cc458ec.png�PNG

   IHDR   d   )   �$��   	pHYs  \F  \F�CA  �IDATx��[hG�Ǹ&�x��FATP�H�T�R��iT��!�>zA��ڂ�WERP�S
���/�A!Ѩ�&^� jLLb���g;ߗ|I^�����Μ��=g�3gv=������ͷ)��7�4æ{[�n5���L��ܦ>~�6�J&�Mr����L�h�݁8U�U3���7۷o�������+�&�c��7�|���bΞ=k�N�j&O�����K�)�Lyy��7o��ݻ�inn���3g�>��3��}����|��Y�`����A��B�}hǰ|o����{���	�=;�2%(--m3fL���2,z���M�oig<��Gj����O��ɦ3�AN�T9�6�j̰��6��Їr�?|��<���;M˼ϟ?���E������oߚ!C��d}dZI�1b����3)@X#G�4���.�"�v�mgPvFF��0@�YŬ��"tc���z���FCC����������!���ӧ"Gm�4�p���2�޽k�3#hC�����6��#d��{���"u�ŋ���:���m����MG�^�@�>�>lc�t����x,#�'�$zh����.��I�Ĩ�$�)$�K�θ���Ϻ���,;ϓ+�
��w��s=��>�~(s�d"�S����cǊ+k�a>�ĉ�p�Ǐe�	����gf͚e���������1c��}����Ҽz�J��2e���L���
�@� ���y�f	�\�zU68
�5i�$�z��`F�7������B���ev��!n"u�F�2�?6;w�W{Ŋf�С����Č�J���6o޼�q׮]2F�{��b��h��
UA��Nf��k�DP�ӧOf۶mf���" Vƽ{�̖-[��˗/7K�.�jۻw�����Ǐ7�w�6}����8qBVбc�̆��ŋ͹s��D���!��e�c���x�X�C00�v��P=�
V�NUoz&�\�u$��������K�.��y�x��0�p8p`�c'�̙c6n�(�H���G��p�ܹ#�k-��Ø0!���I쌄jS[�L��͛7ͦM�Ė=x�@Vl����a�f5�q�m<���O�<1�O�!��O�t������e�e_��0���� �ANN��K
�i	�Ǟ$�a���C��.�\U
���!�Fʸ�
�~�C� �� ���X�v��0�QM��n�:�S�_�N|ucg0�'�1S�j�*3}���K��7��hs��EqU]��̞6m��!T\bM(�6Lht߲r�J�DD>�>|8�U��sg-�A������Em�����`Piii������,�G�LYYYT�SW�l�Cm^4x\555��zK*5��G�� T�֭[�ƍQu��<���S=1l�ɓ'����K�V���x�����2���	Pu�Uf��0^G� ޘ�OcE&��v�3��!x�}��EԳI���S;��p���}I�g�i��UU* �B�ӓ�~xz��2aF�ՂZ#���3���6��aW��X9��l��{Ѯ���5x�D���@to��rVO����
Az��;��@zq��rl�"��z^G�lR=WAD��P�N=�v?щGw�B��B�������o����r���Dm���Lǥ�86����������2~Z�G�1�{��e�8T�?��;w�|���t�A/))�j<{�l�hѢ6��^�O~�E8?_�f��Pl(?�c�8�v��g�~p�k�D"yuuuK�Qii�WTT{ߒ���Mt�h�������TMMM��ͷVUUe���۾��ȍ��nԞ�����}P�Q�[�ϱ�]Z�8�^29��7؅�O���{{���;�[��������ۺBۦ�����U�Z��p�8]v��������4拐�ׯ������]�~b�gϞ���}��G�~�Џ�Qe$��b:�,����B�bl�1�v�����;�"�u�6�=B�4��r    IEND�B`�PK 
     t$v[e�{��~ �~                  cirkitFile.jsonPK 
     t$v[                          jsons/PK 
     t$v[��2��  ��               D jsons/user_defined.jsonPK 
     t$v[                        *b images/PK 
     t$v[z|S�wq wq /             Ob images/b949fd05-6e10-4256-9d1b-e11f1f9900de.pngPK 
     t$v[Ìs�    /             �	 images/01119c27-1bad-421a-afe4-dfb48490a906.pngPK 
     t$v[��Н�� �� /             �	 images/0657d52a-d145-430e-bb7e-5d1be0618b5b.pngPK 
     t$v[T��T$  T$  /             U� images/8ade0660-1c92-4b58-a3e7-adda420d3982.pngPK 
     t$v[��4k� k� /             � images/fd3ac6b5-800b-45c8-a4ce-2476671127d4.pngPK 
     t$v[F���9  �9  /             �� images/915d9337-ea3e-4fec-8caa-7acd53f715e1.pngPK 
     t$v[���HT T /             �� images/00941d67-c746-454a-b945-4fddefc776b2.pngPK 
     t$v[�īd}d  }d  /             @P images/ef87c5cc-d843-475d-a868-97060fb00c54.pngPK 
     t$v[t���?  �?  /             
� images/e2e2c934-b375-45fc-834c-534243cbf361.pngPK 
     t$v[e���  �  /             �� images/6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.pngPK 
     t$v[�;� � /             �� images/31959ea2-aec5-42cb-a646-ec7cb3b6e41e.pngPK 
     t$v[�Ƚׇ  �  /             9
 images/ce527fa2-4558-4370-a5e7-21077342728a.pngPK 
     t$v[�c��f  �f  /              images/cf4cf9a8-07ab-469d-9c7b-0a7a38725bdd.pngPK 
     t$v[��EM  M  /             ;z images/48e84d7e-67ae-4bb6-ba3f-a958722ffd1d.pngPK 
     t$v[������  ��  /             Ս images/27b84e47-6648-4cee-a869-6ff1a6fc12fe.pngPK 
     t$v[�����  �  /             �r images/50196d33-890c-4789-8115-a73c306e50dc.pngPK 
     t$v[��� � /             � images/f158dbb6-f78a-4fb5-8a82-0ff8626242d4.pngPK 
     t$v[��e�/2  /2  /             �� images/0956fa89-558f-410d-92be-91de6d3dc59e.pngPK 
     t$v[�����  ��  /             u� images/2c98734f-75db-43ce-800c-ea69461525e8.pngPK 
     t$v[���z"  "  /             �w images/d4c851cf-9fb5-43cd-809f-e1699313b4d2.pngPK 
     t$v[�e�e�  �  /             -� images/3d0a314b-f708-4b2c-819f-35c414b123ec.pngPK 
     t$v[�kZ��  �  /             �. images/6608fa58-7afa-4488-b64c-2b761d69d6bd.pngPK 
     t$v[9&��ސ ސ /             �B images/b01488b3-8551-4b4c-b09f-2812c4acc168.pngPK 
     t$v[d��   �   /             � images/d3b73945-fe79-451b-b309-b64aab767520.pngPK 
     t$v[��9PN  PN  /             �� images/779eddd4-9cc6-4216-b155-89a4f50be07b.pngPK 
     t$v[w�'<�  �  /             wC images/44e1934a-57d6-434e-9b76-9cc9cf9f98cc.pngPK 
     t$v[wJ���  ��  /             �` images/f9728bc6-2422-4ead-9082-90351081a874.pngPK 
     t$v[	^�G�  �  /             { images/9ba3df0f-d630-43f7-8169-617793654d93.pngPK 
     t$v["1^FHo Ho /             � images/e2a053a3-24a6-43e1-ac97-395cbc045e87.pngPK 
     t$v[��n  n  /             �  images/6b551873-9f16-48c5-b1b9-2fc6ab10f815.pngPK 
     t$v[�9�L� L� /             ٟ  images/b9037746-96b4-41bf-a651-5749520ed4a9.pngPK 
     t$v[;mLP   P   /             r}% images/ded7c6f2-b589-43f4-a4a7-c3e3242414e5.pngPK 
     t$v[U�p�	�  	�  /             �% images/42e39361-2f02-4030-a678-a3271aadd3f6.pngPK 
     t$v[񐼛�  �  /             e>& images/a4af1710-95e2-4b5e-9600-8e4d90487313.pngPK 
     t$v[��r�  �  /             ~R& images/022fab5a-d187-48c2-96d7-20ad2a5d1671.pngPK 
     t$v[6ah    /             |g& images/39d025b2-988a-45cd-b457-87e73cc458ec.pngPK    ( ( �  �o&   
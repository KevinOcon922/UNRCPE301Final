PK
     �9s[���J�O �O    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_0":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_0":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_1":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_1":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_2":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_2":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_3":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_3":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_4":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_5":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_5":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_6":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_6":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_7":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_7":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_8":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_8":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45"],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_9":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_10":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_10":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_11":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_11":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_12":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_12":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_13":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_14":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_14":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_15":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_15":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_16":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_16":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_17":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_17":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_18":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_18":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_19":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_19":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_20":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_20":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_21":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_21":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_22":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_22":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_23":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_23":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_24":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_24":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_25":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_25":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_26":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_26":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_27":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_27":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_28":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_28":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_29":[],"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_29":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29":[],"pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_0":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_1":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_2":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_2":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_3":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_4":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_4":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_5":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_5":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_6":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_6":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_7":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_7":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10":["pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_12":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13":["pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3"],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_16":[],"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_16":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg":["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg":["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg":["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg":["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos":["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg":["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos":["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg":["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-neg":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos":[],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos"],"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-neg":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg"],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-pos":[],"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_0":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_1":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_2":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_3":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_4":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_5":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_6":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_7":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8":["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9":["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_11":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_12":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_13":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_14":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_15":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_16":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_17":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_18":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_19":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_20":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_21":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_22":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_23":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_24":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_25":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_26":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_27":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_32":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_34":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_35":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_36":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_37":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_41":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_42":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44":["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45":["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_50":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_51":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52":["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53":["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54":["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55":["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_56":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_57":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_58":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_59":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3"],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_68":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_69":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_76":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_77":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_78":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_79":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_80":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_81":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_82":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_83":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_84":[],"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_85":[],"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"],"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7"],"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"],"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9"],"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3"],"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4"],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_0":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_1":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_2":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_3":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_4":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_5":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_6":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_7":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_8":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_9":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_10":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_11":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_12":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_13":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_14":[],"pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_15":[],"pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg"],"pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55"],"pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg"],"pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53"],"pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg"],"pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52"],"pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg"],"pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6":[],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7":[],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_8":[],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_9":[],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos"],"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_0":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_2":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_4":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_6":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_8":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_10":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_12":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_14":[],"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14"],"pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10"],"pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13"],"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8"],"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"],"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"],"pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_0":[],"pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_1":[],"pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_2":[],"pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_3":[],"pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_0":[],"pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_1":[],"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"],"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"],"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"],"pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_0":[],"pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1":[],"pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_2":[],"pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_3":[],"pin-type-component_14263f90-2499-4c11-88fb-601766524db5_0":[],"pin-type-component_14263f90-2499-4c11-88fb-601766524db5_1":[],"pin-type-component_14263f90-2499-4c11-88fb-601766524db5_2":[],"pin-type-component_14263f90-2499-4c11-88fb-601766524db5_3":[],"pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_0":[],"pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_1":[],"pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_0":[],"pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_1":[]},"pin_to_color":{"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_0":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_0":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_1":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_1":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_2":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_2":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_3":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_3":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_4":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_5":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_5":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_6":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_6":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_7":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_7":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_8":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_8":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9":"#735348","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_9":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_10":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_10":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_11":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_11":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_12":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_12":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13":"#735348","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_13":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_14":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_14":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_15":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_15":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_16":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_16":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_17":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_17":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_18":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_18":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_19":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_19":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_20":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_20":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_21":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_21":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_22":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_22":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_23":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_23":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_24":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_24":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_25":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_25":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_26":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_26":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_27":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_27":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_28":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_28":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_29":"#000000","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_29":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29":"#000000","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_0":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0":"#FF0000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_1":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1":"#48a1d1","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_2":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_2":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_3":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3":"#189AB4","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_4":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_4":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_5":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_5":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_6":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_6":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_7":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_7":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8":"#90FB92","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9":"#7E2DD2","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10":"#ff3232","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11":"#189AB4","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_12":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13":"#1464c8","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14":"#BDD393","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15":"#FF0000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15":"#0023eb","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_16":"#000000","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_16":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-neg":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos":"#000000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg":"#189AB4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos":"#FF0000","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg":"#189AB4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos":"#FF0000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg":"#189AB4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos":"#FF0000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-neg":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg":"#189AB4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg":"#189AB4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg":"#189AB4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-pos":"#000000","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg":"#189AB4","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_0":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_1":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_2":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_3":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_4":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_5":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_6":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_7":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8":"#dddddd","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9":"#FF6E41","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_11":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_12":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_13":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_14":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_15":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_16":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_17":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_18":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_19":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_20":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_21":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_22":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_23":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_24":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_25":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_26":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_27":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28":"#E85EBE","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29":"#010067","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30":"#9E008E","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31":"#0E4CA1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_32":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33":"#90FB92","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_34":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_35":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_36":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_37":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38":"#FF0000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39":"#189AB4","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40":"#189AB4","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_41":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_42":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44":"#735348","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45":"#735348","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47":"#48a1d1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48":"#BDD393","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49":"#7E2DD2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_50":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_51":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52":"#caca24","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53":"#519355","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54":"#ca2424","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55":"#3885c1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_56":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_57":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_58":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_59":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62":"#FF937E","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63":"#95003A","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64":"#005F39","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65":"#FFE502","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66":"#010067","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67":"#E85EBE","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_68":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_69":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_76":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_77":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_78":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_79":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_80":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_81":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_82":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_83":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_84":"#000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_85":"#000000","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0":"#1642b2","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1":"#ef9cdb","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2":"#eed145","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3":"#f2681c","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4":"#cc1212","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0":"#E85EBE","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1":"#010067","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2":"#9E008E","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3":"#0E4CA1","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4":"#FF0000","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5":"#189AB4","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6":"#1642b2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7":"#ef9cdb","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8":"#eed145","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9":"#f2681c","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10":"#cc1212","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_0":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_1":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_2":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_3":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_4":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_5":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_6":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_7":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_8":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_9":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_10":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_11":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_12":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_13":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_14":"#000000","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_15":"#000000","pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0":"#189AB4","pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1":"#3885c1","pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0":"#189AB4","pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1":"#519355","pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0":"#189AB4","pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1":"#caca24","pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0":"#189AB4","pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1":"#ca2424","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0":"#189AB4","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1":"#FF0000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2":"#FF0000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3":"#E85EBE","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4":"#189AB4","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5":"#010067","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6":"#000000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7":"#000000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_8":"#000000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_9":"#000000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10":"#FFE502","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11":"#005F39","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12":"#95003A","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13":"#FF937E","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14":"#FF0000","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15":"#189AB4","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_0":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_2":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_4":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_6":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_8":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_10":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_12":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13":"#0023eb","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_14":"#000000","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15":"#0023eb","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0":"#ff3232","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1":"#1464c8","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0":"#dddddd","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1":"#FF0000","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2":"#189AB4","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_0":"#000000","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_1":"#000000","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_2":"#000000","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_3":"#000000","pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_0":"#000000","pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_1":"#000000","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0":"#189AB4","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1":"#FF6E41","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2":"#FF0000","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_0":"#000000","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1":"#000000","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_2":"#000000","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_3":"#000000","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_0":"#000000","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_1":"#000000","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_2":"#000000","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_3":"#000000","pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_0":"#000000","pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_1":"#000000","pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_0":"#000000","pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_1":"#000000"},"pin_to_state":{"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_0":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_0":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_1":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_1":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_2":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_2":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_3":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_3":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_4":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_5":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_5":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_6":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_6":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_7":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_7":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_8":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_8":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_9":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_10":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_10":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_11":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_11":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_12":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_12":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_13":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_14":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_14":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_15":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_15":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_16":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_16":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_17":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_17":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_18":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_18":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_19":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_19":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_20":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_20":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_21":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_21":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_22":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_22":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_23":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_23":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_24":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_24":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_25":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_25":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_26":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_26":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_27":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_27":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_28":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_28":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_29":"neutral","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_29":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29":"neutral","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_0":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_1":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_2":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_2":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_3":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_4":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_4":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_5":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_5":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_6":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_6":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_7":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_7":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_12":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_16":"neutral","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_16":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos":"neutral","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-pos":"neutral","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_0":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_1":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_2":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_3":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_4":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_5":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_6":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_7":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_11":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_12":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_13":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_14":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_15":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_16":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_17":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_18":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_19":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_20":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_21":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_22":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_23":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_24":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_25":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_26":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_27":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_32":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_34":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_35":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_36":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_37":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_41":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_42":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_50":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_51":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_56":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_57":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_58":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_59":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_68":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_69":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_76":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_77":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_78":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_79":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_80":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_81":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_82":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_83":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_84":"neutral","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_85":"neutral","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0":"neutral","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1":"neutral","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2":"neutral","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3":"neutral","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9":"neutral","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_0":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_1":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_2":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_3":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_4":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_5":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_6":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_7":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_8":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_9":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_10":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_11":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_12":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_13":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_14":"neutral","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_15":"neutral","pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0":"neutral","pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1":"neutral","pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0":"neutral","pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1":"neutral","pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0":"neutral","pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1":"neutral","pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0":"neutral","pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_8":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_9":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14":"neutral","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_0":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_2":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_4":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_6":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_8":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_10":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_12":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_14":"neutral","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15":"neutral","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0":"neutral","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1":"neutral","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0":"neutral","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1":"neutral","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2":"neutral","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_0":"neutral","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_1":"neutral","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_2":"neutral","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_3":"neutral","pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_0":"neutral","pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_1":"neutral","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0":"neutral","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1":"neutral","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2":"neutral","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_0":"neutral","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1":"neutral","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_2":"neutral","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_3":"neutral","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_0":"neutral","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_1":"neutral","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_2":"neutral","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_3":"neutral","pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_0":"neutral","pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_1":"neutral","pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_0":"neutral","pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_1":"neutral"},"next_color_idx":9,"wires_placed_in_order":[["pin-type-component_d90b98ea-ec54-40fb-811b-0a8df63d2651_1","pin-type-breadboard_c9f5ccf4-1899-4000-97c5-bc5e34b6c93f_0_0"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_0"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_5"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_6"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_7"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_8"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_9"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"],["pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"],["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_1"],["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_b9b7af04-f5f2-421b-a03c-fefac4376a25_0"],["pin-type-component_b9b7af04-f5f2-421b-a03c-fefac4376a25_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"],["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"],["pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_15"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_15","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_13"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_13","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_12"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_12","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"],["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-neg"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-pos"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-pos"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-pos"],["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_29_polarity-pos","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_29_polarity-pos"],["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_29_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_29_polarity-neg"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-neg"],["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_1_polarity-neg"],["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_1_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"],["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"],["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_1_polarity-neg"],["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_2_polarity-neg"],["pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_3_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_1_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_4","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_10_polarity-neg"],["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_5_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_6_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_4","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_15","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_14","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_14","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-pos"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_15","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-neg"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_1f1f15d7-582d-46c6-8062-134460c0cfb1_4"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg"],["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos"],["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg"],["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg"],["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40"],["pin-type-component_ae8acd73-fbc2-438c-bd1a-16ad65be65d2_3","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15"],["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg"],["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg"],["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg"],["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg"],["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52"],["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53"],["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54"],["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg"],["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63"],["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"],["pin-type-component_c034544e-ef8e-4127-909d-5c85a081ec0e_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"],["pin-type-component_c034544e-ef8e-4127-909d-5c85a081ec0e_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"],["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"],["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"],["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg"],["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos"],["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"],["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg","pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_3"],["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"],["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_0","pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_0"],["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_1","pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_1"],["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos"],["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33"],["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"],["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"],["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14"],["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1"],["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos"],["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11"],["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15"],["pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4"],["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20"],["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45"],["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"],["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"],["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"],["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"],["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9"],["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[["pin-type-component_d90b98ea-ec54-40fb-811b-0a8df63d2651_1","pin-type-breadboard_c9f5ccf4-1899-4000-97c5-bc5e34b6c93f_0_0"]]],[[["pin-type-breadboard_c9f5ccf4-1899-4000-97c5-bc5e34b6c93f_0_0","pin-type-component_d90b98ea-ec54-40fb-811b-0a8df63d2651_1"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_0"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_0"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_5"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_6"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_7"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_8"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_9"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"]],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"]]],[[],[["pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_0"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]]],[[],[["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_1"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_1"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_b5fd5d86-c9a9-42df-91a5-a8683ed12120_0"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_1"]]],[[],[["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_b9b7af04-f5f2-421b-a03c-fefac4376a25_0"]]],[[],[["pin-type-component_b9b7af04-f5f2-421b-a03c-fefac4376a25_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_b9b7af04-f5f2-421b-a03c-fefac4376a25_0"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62","pin-type-component_b9b7af04-f5f2-421b-a03c-fefac4376a25_1"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"]],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"]]],[[],[["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"]]],[[],[["pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_15"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_15","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_13"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_13","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_12"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_12","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0"]]],[[],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_12"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_12","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_13"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_13","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_15"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_15","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_16"]],[]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10"]]],[[],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_0","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"],["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_2","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_2","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_3","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_3","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_5"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_4","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_4","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_6"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_5","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_7"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_6","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_8"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_7","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_9"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_8","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_9","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_10","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"],["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"],["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"],["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_11","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_1_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38"]],[]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_12","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_13","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_14","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15","pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16"],["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_15","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]]],[[["pin-type-breadboard_2c0029e7-54e1-4817-822e-cdaaeeebc81e_0_16","pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0"]],[]],[[["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39"]],[]],[[["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0"]],[]],[[["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-neg"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-pos"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-pos"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-neg"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-pos"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-pos"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-pos"]]],[[],[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_29_polarity-pos","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_29_polarity-pos"]]],[[],[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_29_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_29_polarity-neg"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-neg"]]],[[],[["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_1_polarity-neg"]]],[[],[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_1_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"]]],[[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_1_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"]],[]],[[["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_1_polarity-neg"]],[]],[[],[["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"]]],[[],[["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_1_polarity-neg"]]],[[],[["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_2_polarity-neg"]]],[[],[["pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_3_polarity-neg"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"]]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-pos"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_1_polarity-pos"]]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_1_polarity-pos"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-pos"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-pos"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-pos"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_4","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_10_polarity-neg"]]],[[],[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"]]],[[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"]]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-pos"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_4","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_10_polarity-neg"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-pos"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_5_polarity-pos"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_6_polarity-pos"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_4","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_15","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-neg"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_14","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-pos"]]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_15","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-neg"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_14","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-pos"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_14","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-pos"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_15","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-neg"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_13"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_12"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_11"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60","pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_1"]],[]],[[["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62","pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_1"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63","pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_1"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_5"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_3"]],[]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"]]],[[],[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"]]],[[["pin-type-component_ef32751e-db38-4691-a34f-2587734b054d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_0_polarity-neg"]],[]],[[["pin-type-component_730f6843-7c62-43fc-860e-8f09589d638d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_1_polarity-neg"]],[]],[[],[]],[[["pin-type-component_e70cd174-2eb7-448e-b301-6cb6ab1d5bfb_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_2_polarity-neg"]],[]],[[["pin-type-component_f07feec7-27f2-4fc8-8cd6-79c12796e38e_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_3_polarity-neg"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_1","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_5_polarity-pos"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_0","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_4_polarity-neg"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_2","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_6_polarity-pos"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_4","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_7_polarity-neg"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_14","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_8_polarity-pos"]],[]],[[["pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_15","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_9_polarity-neg"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-pos"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_0_polarity-neg"]],[]],[[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_29_polarity-pos","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_29_polarity-pos"]],[]],[[["pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_0_29_polarity-neg","pin-type-power-rail_58b0017f-e758-4a6b-9e36-e6b051240d70_1_29_polarity-neg"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_3"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_5"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_10"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_11"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_12"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47","pin-type-component_964f8ed7-2d56-4f26-97a9-ab33e355803d_13"]],[]],[[],[]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_1f1f15d7-582d-46c6-8062-134460c0cfb1_4"]]],[[["pin-type-component_1f1f15d7-582d-46c6-8062-134460c0cfb1_4","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0"]],[]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"]]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4"]],[]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"]]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2"]],[]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos"]]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg"]]],[[],[["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos"]]],[[],[["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg"]]],[[],[["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_ae8acd73-fbc2-438c-bd1a-16ad65be65d2_3","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15"]]],[[["pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15","pin-type-component_ae8acd73-fbc2-438c-bd1a-16ad65be65d2_3"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg"]]],[[],[["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg"]]],[[],[["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg"]]],[[],[["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg"]]],[[],[["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52"]]],[[],[["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53"]]],[[],[["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54"]]],[[],[["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"]]],[[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"]],[]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"]]],[[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg"]]],[[],[["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"]]],[[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos"]],[]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64"]]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6"]],[]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63"]]],[[],[["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"]]],[[],[["pin-type-component_c034544e-ef8e-4127-909d-5c85a081ec0e_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"]]],[[],[["pin-type-component_c034544e-ef8e-4127-909d-5c85a081ec0e_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"]]],[[["pin-type-component_c034544e-ef8e-4127-909d-5c85a081ec0e_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"]],[]],[[["pin-type-component_c034544e-ef8e-4127-909d-5c85a081ec0e_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"]],[]],[[],[["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"]]],[[],[["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"]]],[[],[["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8"]]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos"]]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos"]],[]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos"]]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"]]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"]],[]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10"]]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"]]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos"]],[]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"]],[]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10"]],[]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"]]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"]],[]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg"]]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"]]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg"]],[]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"]],[]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg"]]],[[],[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos"]]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos"]],[]],[[["pin-type-component_5aa9b9e9-ad09-4d35-b1a8-7a7b8e670cfb_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg"]],[]],[[],[["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"]]],[[["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg"]],[]],[[],[["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg","pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_3"]]],[[],[["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"]]],[[],[["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_0","pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_0"]]],[[],[["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_1","pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_1"]]],[[["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_0","pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_0"],["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"]],[["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"]]],[[["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_1","pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_1"]],[]],[[["pin-type-component_8c10ff73-740f-4886-be5b-c94a7bcbfbd0_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg"]],[]],[[["pin-type-component_350eb403-34b4-46e7-be78-ea7d63f1f722_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos"]],[]],[[],[["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49"]],[]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33"]]],[[],[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"]]],[[],[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"]]],[[],[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1"]],[]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13"]],[]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14"]]],[[],[["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15"]]],[[],[]],[[],[]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49"]],[]],[[],[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos"]]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos"]],[]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg"]],[]],[[],[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos"]]],[[["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos"]],[]],[[],[["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11"]]],[[],[["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4"]]],[[["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20"]]],[[["pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45"]]],[[],[["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"]]],[[],[]],[[],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"]],[]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"]],[]],[[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"]],[]],[[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"]],[]],[[["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"]]],[[],[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"]]],[[],[["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos"]]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos"]],[]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"]]],[[],[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"]]],[[["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2"]],[]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9"]]],[[],[["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_0":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_0":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_1":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_1":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_2":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_2":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_3":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_3":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_4":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_4":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_5":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_5":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_6":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_6":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_7":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_7":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_8":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_8":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9":"0000000000000061","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_9":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_10":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_10":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_11":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_11":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_12":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_12":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13":"0000000000000062","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_13":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_14":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_14":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_15":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_15":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_16":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_16":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_17":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_17":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_18":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_18":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_19":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_19":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_20":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_20":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_21":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_21":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_22":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_22":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_23":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_23":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_24":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_24":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_25":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_25":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_26":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_26":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_27":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_27":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_28":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_28":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_29":"_","pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_1_29":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29":"_","pin-type-breadboard_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_0":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0":"0000000000000040","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_1":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1":"0000000000000042","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_2":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_2":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_3":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3":"0000000000000041","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_4":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_4":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_5":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_5":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_6":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_6":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_7":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_7":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8":"0000000000000054","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8":"0000000000000046","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9":"0000000000000055","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9":"0000000000000047","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10":"0000000000000057","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10":"0000000000000048","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11":"0000000000000058","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11":"0000000000000049","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_12":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12":"0000000000000051","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13":"0000000000000060","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13":"0000000000000050","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14":"0000000000000056","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14":"0000000000000052","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15":"0000000000000059","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15":"0000000000000053","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_16":"_","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_16":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos":"0000000000000009","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg":"0000000000000010","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_0_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg":"0000000000000016","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_1_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg":"0000000000000017","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_2_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg":"0000000000000018","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_3_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg":"0000000000000019","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_4_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_5_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_5_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_6_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_6_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_7_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_7_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_8_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_8_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_9_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_10_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_10_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_11_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_11_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_12_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_12_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_13_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_14_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_14_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_15_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_15_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_16_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos":"0000000000000002","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_17_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg":"0000000000000001","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_18_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg":"0000000000000041","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_19_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos":"0000000000000040","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_20_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_20_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_21_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos":"0000000000000038","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_22_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg":"0000000000000037","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_23_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg":"0000000000000032","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_24_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos":"0000000000000031","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_25_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg":"0000000000000029","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_26_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos":"0000000000000027","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_27_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos":"0000000000000026","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_28_polarity-neg":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-pos":"_","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg":"0000000000000025","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos":"0000000000000011","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg":"0000000000000012","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos":"0000000000000011","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg":"0000000000000012","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_0_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_0_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_1_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_1_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_2_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_2_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_3_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_3_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_4_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_4_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_5_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_5_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_6_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_6_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_7_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_7_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_8_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_8_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_9_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_9_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_10_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_10_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_11_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_11_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_12_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_12_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_13_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_13_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_14_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_14_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_15_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_15_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_16_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_16_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_17_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_17_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_18_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_18_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_19_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_19_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_20_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_20_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_21_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_21_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_22_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_22_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_23_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_23_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_24_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_24_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos":"0000000000000005","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_25_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg":"0000000000000004","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_26_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos":"0000000000000059","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_27_polarity-neg":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg":"0000000000000058","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg":"0000000000000013","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg":"0000000000000014","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-pos":"_","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg":"0000000000000014","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_0":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_1":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_2":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_3":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_4":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_5":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_6":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_7":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8":"0000000000000039","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9":"0000000000000000","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_10":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_11":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_12":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_13":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_14":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_15":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_16":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_17":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_18":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_19":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_20":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_21":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_22":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_23":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_24":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_25":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_26":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_27":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28":"0000000000000003","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29":"0000000000000006","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30":"0000000000000007","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31":"0000000000000008","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_32":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33":"0000000000000054","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_34":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_35":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_36":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_37":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38":"0000000000000009","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39":"0000000000000010","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40":"0000000000000013","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_41":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_42":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_43":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44":"0000000000000062","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45":"0000000000000061","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_46":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47":"0000000000000042","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48":"0000000000000056","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49":"0000000000000055","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_50":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_51":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52":"0000000000000020","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53":"0000000000000021","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54":"0000000000000022","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55":"0000000000000023","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_56":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_57":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_58":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_59":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_60":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_61":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62":"0000000000000036","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63":"0000000000000035","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64":"0000000000000034","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65":"0000000000000033","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66":"0000000000000030","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67":"0000000000000028","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_68":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_69":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_70":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_71":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_72":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_73":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_74":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_75":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_76":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_77":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_78":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_79":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_80":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_81":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_82":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_83":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_84":"_","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_85":"_","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0":"0000000000000015","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1":"0000000000000024","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2":"0000000000000045","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3":"0000000000000044","pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4":"0000000000000043","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0":"0000000000000003","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1":"0000000000000006","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2":"0000000000000007","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3":"0000000000000008","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4":"0000000000000005","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5":"0000000000000004","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6":"0000000000000015","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7":"0000000000000024","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8":"0000000000000045","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9":"0000000000000044","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10":"0000000000000043","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_0":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_1":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_2":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_3":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_4":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_5":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_6":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_7":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_8":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_9":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_10":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_11":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_12":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_13":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_14":"_","pin-type-component_88075651-101d-4b77-9d5b-8861a83896c1_15":"_","pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0":"0000000000000019","pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1":"0000000000000023","pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0":"0000000000000017","pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1":"0000000000000021","pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0":"0000000000000016","pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1":"0000000000000020","pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0":"0000000000000018","pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1":"0000000000000022","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0":"0000000000000025","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1":"0000000000000026","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2":"0000000000000027","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3":"0000000000000028","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4":"0000000000000029","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5":"0000000000000030","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_6":"_","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_7":"_","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_8":"_","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_9":"_","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10":"0000000000000033","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11":"0000000000000034","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12":"0000000000000035","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13":"0000000000000036","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14":"0000000000000031","pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15":"0000000000000032","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_0":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1":"0000000000000046","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_2":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3":"0000000000000053","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_4":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5":"0000000000000047","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_6":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7":"0000000000000048","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_8":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9":"0000000000000049","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_10":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11":"0000000000000051","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_12":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13":"0000000000000050","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_14":"_","pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15":"0000000000000052","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0":"0000000000000057","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1":"0000000000000060","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0":"0000000000000039","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1":"0000000000000038","pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2":"0000000000000037","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_0":"_","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_1":"_","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_2":"_","pin-type-component_aadcf1a0-67b3-4a34-8461-766def044c41_3":"_","pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_0":"_","pin-type-component_912f99f9-1a7b-4d96-904c-46d72b192ca7_1":"_","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0":"0000000000000001","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1":"0000000000000000","pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2":"0000000000000002","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_0":"_","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_1":"_","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_2":"_","pin-type-component_c37a5152-d1df-4c89-bbc1-31eea23fe6a5_3":"_","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_0":"_","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_1":"_","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_2":"_","pin-type-component_14263f90-2499-4c11-88fb-601766524db5_3":"_","pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_0":"_","pin-type-component_d3b14dfa-8357-4d45-8fa7-81e44c3574de_1":"_","pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_0":"_","pin-type-component_f9a354fb-a5e8-4c85-bf60-2ac09a3d1443_1":"_"},"component_id_to_pins":{"802528b6-1c68-4132-8eb3-ef45339a8beb":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37","38","39","40","41","42","43","44","45","46","47","48","49","50","51","52","53","54","55","56","57","58","59","60","61","62","63","64","65","66","67","68","69","70","71","72","73","74","75","76","77","78","79","80","81","82","83","84","85"],"e5348ec8-9804-4ec3-98a4-c934e85c4b49":["0","1","2","3","4"],"59718622-87ae-47c5-ab64-77f43e28c079":["0","1","2","3","4","5","6","7","8","9","10"],"88075651-101d-4b77-9d5b-8861a83896c1":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"d31a6738-5eba-41b7-bcd4-00ce53bb91e4":["0","1"],"317b37d2-20d2-4d51-9e3b-72e93df3ce83":["0","1"],"e33041df-846d-4953-b931-56a7b8227815":["0","1"],"29b8e01a-285a-4675-b6e8-5a3c24817ccc":["0","1"],"fd8f8cb1-e823-496b-ad06-7cf0fbacd90f":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"22bfc2f4-ec74-4e25-b5ac-80edc339190c":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"127fe76f-620d-42d3-bc33-d5252ff1a787":["0","1"],"d1c6c4d4-8ab8-4ab8-a980-754c86362baa":["0","1","2"],"aadcf1a0-67b3-4a34-8461-766def044c41":["0","1","2","3"],"912f99f9-1a7b-4d96-904c-46d72b192ca7":["0","1"],"ea1a6d9b-043c-42f4-95db-9fdb3e699131":["0","1","2"],"c37a5152-d1df-4c89-bbc1-31eea23fe6a5":["0","1","2","3"],"14263f90-2499-4c11-88fb-601766524db5":["0","1","2","3"],"d3b14dfa-8357-4d45-8fa7-81e44c3574de":["0","1"],"f9a354fb-a5e8-4c85-bf60-2ac09a3d1443":["0","1"]},"uid_to_net":{"_":[],"0000000000000009":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos"],"0000000000000010":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg"],"0000000000000011":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos"],"0000000000000012":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg"],"0000000000000016":["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg"],"0000000000000017":["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg"],"0000000000000018":["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg"],"0000000000000019":["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg"],"0000000000000020":["pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52"],"0000000000000021":["pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53"],"0000000000000022":["pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54"],"0000000000000023":["pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55"],"0000000000000013":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg"],"0000000000000014":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg"],"0000000000000025":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg"],"0000000000000026":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos"],"0000000000000027":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos"],"0000000000000028":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67"],"0000000000000029":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg"],"0000000000000030":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66"],"0000000000000031":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos"],"0000000000000032":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg"],"0000000000000033":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65"],"0000000000000034":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64"],"0000000000000035":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63"],"0000000000000036":["pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62"],"0000000000000037":["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg"],"0000000000000038":["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos"],"0000000000000039":["pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8"],"0000000000000040":["pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0"],"0000000000000041":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg"],"0000000000000046":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8"],"0000000000000047":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9"],"0000000000000048":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10"],"0000000000000049":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11"],"0000000000000050":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13"],"0000000000000051":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12"],"0000000000000052":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14"],"0000000000000053":["pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15"],"0000000000000042":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1"],"0000000000000054":["pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8"],"0000000000000055":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49"],"0000000000000056":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48"],"0000000000000057":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0"],"0000000000000060":["pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13","pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1"],"0000000000000058":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11"],"0000000000000059":["pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos","pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15"],"0000000000000061":["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45"],"0000000000000062":["pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44"],"0000000000000000":["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9"],"0000000000000001":["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg"],"0000000000000002":["pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2","pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos"],"0000000000000003":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28"],"0000000000000004":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg"],"0000000000000005":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4","pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos"],"0000000000000006":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29"],"0000000000000007":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30"],"0000000000000008":["pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3","pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31"],"0000000000000015":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6"],"0000000000000024":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7"],"0000000000000043":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10"],"0000000000000044":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9"],"0000000000000045":["pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2","pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8"]},"uid_to_text_label":{"0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000021":"Net 21","0000000000000022":"Net 22","0000000000000023":"Net 23","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000025":"Net 25","0000000000000026":"Net 26","0000000000000027":"Net 27","0000000000000028":"Net 28","0000000000000029":"Net 29","0000000000000030":"Net 30","0000000000000031":"Net 31","0000000000000032":"Net 32","0000000000000033":"Net 33","0000000000000034":"Net 34","0000000000000035":"Net 35","0000000000000036":"Net 36","0000000000000037":"Net 37","0000000000000038":"Net 38","0000000000000039":"Net 39","0000000000000040":"Net 40","0000000000000041":"Net 41","0000000000000046":"Net 46","0000000000000047":"Net 47","0000000000000048":"Net 48","0000000000000049":"Net 49","0000000000000050":"Net 50","0000000000000051":"Net 51","0000000000000052":"Net 52","0000000000000053":"Net 53","0000000000000042":"Net 42","0000000000000054":"Net 54","0000000000000055":"Net 55","0000000000000056":"Net 56","0000000000000057":"Net 57","0000000000000060":"Net 60","0000000000000058":"Net 58","0000000000000059":"Net 59","0000000000000061":"Net 61","0000000000000062":"Net 62","0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000015":"Net 15","0000000000000024":"Net 24","0000000000000043":"Net 43","0000000000000044":"Net 44","0000000000000045":"Net 45"},"all_breadboard_info_list":["c9f5ccf4-1899-4000-97c5-bc5e34b6c93f_30_2_True_939.4999999999993_-529.5000000000002_left","2c0029e7-54e1-4817-822e-cdaaeeebc81e_17_2_False_241.99999999999994_317.99999999999983_left","58b0017f-e758-4a6b-9e36-e6b051240d70_30_2_True_205_399.99999999999994_up","08c4f86b-8832-45bd-8fa3-b796555329d7_63_2_True_235_460_up","246c73ed-c3aa-4493-99a9-e79818341acd_30_2_True_235_295_up","2622c028-5eeb-487e-a780-ae7d5e5671cc_30_2_True_309.5_745.4999999999999_left","d229e1a5-25f8-4573-81e5-290fe5d1779f_17_2_False_655_280_up","7425f490-20e5-405c-8f1e-bcd16b84ce42_17_2_False_842.0000000000001_-282.0000000000001_left","7cabb3b8-0cac-490c-b7b1-faa9382fcc19_17_2_False_812_828.0000000000001_left"],"breadboard_info_list":["246c73ed-c3aa-4493-99a9-e79818341acd_30_2_True_235_295_up","2622c028-5eeb-487e-a780-ae7d5e5671cc_30_2_True_309.5_745.4999999999999_left","7425f490-20e5-405c-8f1e-bcd16b84ce42_17_2_False_842.0000000000001_-282.0000000000001_left"],"componentsData":[{"compProperties":{},"position":[1165.936459,830.0020834999998],"typeId":"de09217e-3b73-b82d-0145-70b2df9a4b72","componentVersion":1,"instanceId":"e5348ec8-9804-4ec3-98a4-c934e85c4b49","orientation":"right","circleData":[[917.5,800],[917.5,814.9979165],[917.5,830.0020835],[917.5,844.998959],[917.5,859.9989590000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[816.2844175,866.1994415000005],"typeId":"ecbd5bee-2226-4f1c-8fdb-aaff666e8628","componentVersion":1,"instanceId":"59718622-87ae-47c5-ab64-77f43e28c079","orientation":"left","circleData":[[767.5,815],[767.5,829.4904139999999],[766.0509640000001,842.531792],[766.0509640000001,855.5731115000001],[795.8902765000001,920.5741939999998],[781.4944090000001,921.4738984999993],[844.4762799999996,803.6079139999999],[843.5765154999999,816.2042525000002],[843.5765154999999,827.9008865000001],[843.5765154999999,839.5975205],[842.6768109999998,853.0936220000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[126.9183789999996,972.1184914999994],"typeId":"307d45d2-aa1f-05de-326e-55c453eb206e","componentVersion":4,"instanceId":"88075651-101d-4b77-9d5b-8861a83896c1","orientation":"down","circleData":[[197.5,1115],[197.5,1100],[137.5,1115],[137.5,1100],[197.3499999999999,846.1999999999989],[197.3499999999998,830.899999999999],[137.61942699999986,846.1847134999989],[137.63471349999986,831.019426999999],[181.89999999999986,1025.3000000000002],[166.89999999999986,1025.3000000000002],[151.89999999999986,1025.3000000000002],[136.89999999999986,1025.3000000000002],[181.89999999999986,1010.3000000000001],[166.89999999999986,1010.3000000000001],[151.89999999999986,1010.3000000000001],[136.89999999999986,1010.3000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[388.78038849999973,72.50001799999981],"typeId":"972688b5-e2a3-1d53-e820-bc24d2f5082a","componentVersion":15,"instanceId":"802528b6-1c68-4132-8eb3-ef45339a8beb","orientation":"up","circleData":[[542.5,215],[557.4999819999998,215],[572.4978805000005,215],[587.5020295000006,215],[602.5020115000007,215],[617.4999115,215],[632.4998935000008,215],[647.4977920000003,215],[407.5001574999998,215],[422.49805749999973,215],[437.50220649999983,215],[452.50218849999965,215],[467.50008699999967,215],[482.50007049999977,215],[497.49796899999996,215],[512.5021180000001,215],[617.4999115,-70],[602.5020115000007,-70],[587.5020295000006,-70],[572.4978805000005,-70],[557.4999819999998,-70],[542.5,-70],[527.5021000000004,-70],[512.5021180000001,-70],[218.4982974999997,-70],[233.50036299999977,-70],[248.5003449999997,-70],[263.50032699999974,-70],[278.5003104999997,-70],[293.5002924999998,-70],[308.5002744999997,-70],[323.50025649999975,-70],[338.50023999999974,-70],[353.5002219999998,-70],[272.5003164999997,215],[287.5002999999997,215],[302.50236549999977,215],[317.5002639999997,215],[332.5002459999997,215],[347.50022799999977,215],[362.50021149999964,215],[377.5022769999997,215],[482.50007049999977,-70],[467.50008699999967,-70],[452.50218849999965,-70],[437.50220649999983,-70],[422.49805749999973,-70],[407.5001574999998,-70],[392.5001754999997,-70],[377.5022769999997,-70],[662.5019410000004,-70],[677.5019245000005,-70],[662.5019410000004,-55],[677.5019245000005,-55],[662.5019410000004,-40],[677.5019245000005,-40],[662.5019410000004,-25],[677.5019245000005,-25],[662.5019410000004,-10],[677.5019245000005,-10],[662.5019410000004,4.999999999999943],[677.5019245000005,4.999999999999943],[662.5019410000004,19.999999999999943],[677.5019245000005,19.999999999999943],[662.5019410000004,34.99999999999994],[677.5019245000005,34.99999999999994],[662.5019410000004,49.99999999999994],[677.5019245000005,49.99999999999994],[662.5019410000004,64.99999999999994],[677.5019245000005,64.99999999999994],[662.5019410000004,80.00000000000009],[677.5019245000005,80.00000000000009],[662.5019410000004,95.00000000000017],[677.5019245000005,95.00000000000017],[662.5019410000004,110.00000000000031],[677.5019245000005,110.00000000000031],[662.5019410000004,125.00000000000011],[677.5019245000005,125.00000000000011],[662.5019410000004,140.0000000000004],[677.5019245000005,140.0000000000004],[662.5019410000004,155.0000000000004],[677.5019245000005,155.0000000000004],[662.5019410000004,170.00000000000068],[677.5019245000005,170.00000000000068],[662.5019410000004,185.00000000000045],[677.5019245000005,185.00000000000045]],"code":"512,folder,{\"name\":\"sketch\",\"id\":\"47fa4ae5-8c4a-447b-a0e7-1e0b4e1aec2f\",\"explorerHtmlId\":\"13443a0f-75f4-4f9e-8ab3-f4f93fa01743\",\"nameHtmlId\":\"591d9dd3-ee94-4962-9f7a-6b0f401a3ef5\",\"nameInputHtmlId\":\"f8285722-3ac9-4555-85bf-85447299cb63\",\"explorerChildHtmlId\":\"7870fa5e-e923-4166-b0d8-19e3144686b6\",\"explorerCarrotOpenHtmlId\":\"9b1f7211-e75f-48c0-8b93-b555b65ffa4e\",\"explorerCarrotClosedHtmlId\":\"4429e12f-176a-47b8-beb0-a5cd97894707\",\"arduinoBoardFqbn\":\"arduino:avr:mega\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"feb43c4c-7472-47a9-86db-a1ef8cd6ebca\",\"explorerHtmlId\":\"1426fd4a-ab41-4e9b-8ace-bac64390decf\",\"nameHtmlId\":\"19d457e9-b845-4325-8134-185a2f11ad0e\",\"nameInputHtmlId\":\"b66b01d2-f19d-4d99-aaa2-ffe51becf8ed\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"e812fc5e-467b-4844-924e-dc6f4209fc94\",\"explorerHtmlId\":\"0ab4292a-45c5-4745-b729-edc2179e3445\",\"nameHtmlId\":\"611279a6-db2f-47be-b806-ee42712a99ff\",\"nameInputHtmlId\":\"13f8e070-def3-4a62-a251-7dde8b6d0e66\",\"code\":\"\"},0,","codeLabelPosition":[388.78038849999945,-84.98588200000015],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[565.0478665,-292.79700099999997],"typeId":"5f0a7f7f-5908-4e39-94d8-2714a0462581","componentVersion":2,"instanceId":"29b8e01a-285a-4675-b6e8-5a3c24817ccc","orientation":"up","circleData":[[557.5,-265],[572.5,-265]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[627.5000245000002,-292.4999934999999],"typeId":"117aab52-1b06-40f5-98b6-df63a601b0e6","componentVersion":3,"instanceId":"d31a6738-5eba-41b7-bcd4-00ce53bb91e4","orientation":"up","circleData":[[617.5,-250],[640.7613849999999,-250.12790800000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[507.5000245,-292.49997549999983],"typeId":"a70bb5a8-99ed-4f1b-882e-eac0873b75ef","componentVersion":5,"instanceId":"317b37d2-20d2-4d51-9e3b-72e93df3ce83","orientation":"up","circleData":[[497.5,-250.00000000000006],[520.7613849999998,-250.12790950000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[432.5000245000001,-292.5000114999997],"typeId":"1310de1e-180e-4aed-a1c6-f80032a2bfde","componentVersion":4,"instanceId":"e33041df-846d-4953-b931-56a7b8227815","orientation":"up","circleData":[[422.5,-250.00000000000006],[445.7613849999998,-250.127908]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1296.0726505,-200.6876064999998],"typeId":"7115dd0c-9076-1603-96e1-f4f66aa483df","componentVersion":7,"instanceId":"127fe76f-620d-42d3-bc33-d5252ff1a787","orientation":"up","circleData":[[1112.5,-250],[1112.5,-151.1619999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"","type":"string","value":"10000","displayFormat":"dropdown","options":[{"label":"1000","value":"1000"},{"label":"10000","value":"10000"},{"label":"50000","value":"50000"},{"label":"100000","value":"100000"}],"showOnComp":false,"isVisibleToUser":true}},"position":[542.4531325000002,303.92501600000014],"typeId":"7013093c-3557-9fba-53d2-85a05ece47f1","componentVersion":1,"instanceId":"ea1a6d9b-043c-42f4-95db-9fdb3e699131","orientation":"up","circleData":[[527.5,365],[542.4958405000001,365.00416700000005],[557.5093914999999,365]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"181","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[1256.4770755000002,306.53440850000015],"typeId":"23598c1c-7607-4538-b177-9ab948fb1937","componentVersion":3,"instanceId":"fd8f8cb1-e823-496b-ad06-7cf0fbacd90f","orientation":"up","circleData":[[1067.5,215],[1082.5020834999998,215],[1097.5,215],[1112.5,215],[1127.5020835,215],[1142.5,215],[1157.5020835,215],[1172.5,215],[1187.5,215],[1202.5,215],[1217.5,215],[1232.5020835,215],[1247.5,215],[1262.4999999999998,215],[1277.5020834999998,215],[1292.4999999999993,215]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"PTS645SL50-2 LFS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"C&K Components","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[280.00149999999985,425.2295000000002],"typeId":"232ac546-6e45-4194-9a27-0fa614949a21","componentVersion":3,"instanceId":"c37a5152-d1df-4c89-bbc1-31eea23fe6a5","orientation":"right","circleData":[[302.5,440],[257.4999999999998,440],[302.5,410.0000000000003],[257.4999999999998,410.0000000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"PTS645SL50-2 LFS","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"mpn","unit":"","userVisible":false,"required":true},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"C&K Components","displayFormat":"input","showOnComp":false,"isVisibleToUser":false,"name":"manufacturer","unit":"","userVisible":false,"required":true}},"position":[280.00149999999985,485.2294999999999],"typeId":"232ac546-6e45-4194-9a27-0fa614949a21","componentVersion":3,"instanceId":"14263f90-2499-4c11-88fb-601766524db5","orientation":"right","circleData":[[302.5,500],[257.4999999999997,500],[302.5,469.99999999999994],[257.4999999999997,469.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4700","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[370,470],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"f9a354fb-a5e8-4c85-bf60-2ac09a3d1443","orientation":"up","circleData":[[332.5,470],[407.5,470]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1300.4165050000004,512.7833300000005],"typeId":"97784b10-4dcd-a3be-9167-75f1272c8490","componentVersion":1,"instanceId":"d1c6c4d4-8ab8-4ab8-a980-754c86362baa","orientation":"left","circleData":[[1127.5,530],[1127.5,515.0000000000007],[1127.5,500.0000000000007]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4700","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[370,410],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"d3b14dfa-8357-4d45-8fa7-81e44c3574de","orientation":"up","circleData":[[332.5,410],[407.5,410]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[940.0000000000005,-151.49500149999994],"typeId":"155f7657-2d2d-eaf2-280f-5c76a41d0679","componentVersion":1,"instanceId":"22bfc2f4-ec74-4e25-b5ac-80edc339190c","orientation":"up","circleData":[[887.5000000000005,-130],[887.5000000000005,-172.9900029999998],[992.5000015000004,-130],[992.5000015000004,-172.9900029999998],[902.5000000000005,-130],[902.5000000000005,-172.9900029999998],[917.5000000000005,-130],[917.5000000000005,-172.9900029999998],[932.5000000000005,-130],[932.5000000000005,-172.9900029999998],[947.5000015000005,-130],[947.5000015000005,-172.9900029999998],[962.5000015000005,-130],[962.5000015000005,-172.9900029999998],[977.5000015000005,-130],[977.5000015000005,-172.9900029999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[789.9999984999998,-279.9999159999999],"typeId":"a76bb123-3d3c-417d-b1f3-c8417efb7bc7","componentVersion":1,"instanceId":"aadcf1a0-67b3-4a34-8461-766def044c41","orientation":"up","circleData":[[767.4999999999999,-220],[782.4999999999999,-220],[797.4999999999999,-220],[812.4999999999998,-220]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}},"position":[768.286318110109,-195.8785402787413],"typeId":"1c569fa1-772b-452c-b113-493dd976b9c0","componentVersion":7,"instanceId":"912f99f9-1a7b-4d96-904c-46d72b192ca7","orientation":"up","circleData":[[767.4999999999999,-205],[782.4999999999999,-205]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-365.00006","left":"32.43015","width":"1475.16825","height":"1493.61460","x":"32.43015","y":"-365.00006"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_38\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"332.5002460000_215.0000000000\\\",\\\"332.5002460000_245.0000000000\\\",\\\"137.5000000000_245.0000000000\\\",\\\"137.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_39\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"347.5002280000_215.0000000000\\\",\\\"347.5002280000_260.0000000000\\\",\\\"152.5000000000_260.0000000000\\\",\\\"152.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos\",\"rawStartPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-pos\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"137.5000000000_740.0000000000\\\",\\\"137.5000000000_777.5000000000\\\",\\\"407.5000000000_777.5000000000\\\",\\\"407.5000000000_740.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_29_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_29_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"152.5000000000_740.0000000000\\\",\\\"152.5000000000_792.5000000000\\\",\\\"422.5000000000_792.5000000000\\\",\\\"422.5000000000_740.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg\",\"rawStartPinId\":\"pin-type-component_e33041df-846d-4953-b931-56a7b8227815_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_1_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"422.5000000000_-250.0000000000\\\",\\\"17.5000000000_-250.0000000000\\\",\\\"17.5000000000_320.0000000000\\\",\\\"152.5000000000_320.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg\",\"rawStartPinId\":\"pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_2_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"497.5000000000_-250.0000000000\\\",\\\"497.5000000000_-235.0000000000\\\",\\\"2.5000000000_-235.0000000000\\\",\\\"2.5000000000_335.0000000000\\\",\\\"152.5000000000_335.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg\",\"rawStartPinId\":\"pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_3_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5000000000_-265.0000000000\\\",\\\"557.5000000000_-220.0000000000\\\",\\\"-12.5000000000_-220.0000000000\\\",\\\"-12.5000000000_350.0000000000\\\",\\\"152.5000000000_350.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg\",\"rawStartPinId\":\"pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_0_4_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-250.0000000000\\\",\\\"617.5000000000_-205.0000000000\\\",\\\"-27.5000000000_-205.0000000000\\\",\\\"-27.5000000000_365.0000000000\\\",\\\"152.5000000000_365.0000000000\\\"]}\"}","{\"color\":\"#caca24\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52\",\"endPinId\":\"pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_52\",\"rawEndPinId\":\"pin-type-component_e33041df-846d-4953-b931-56a7b8227815_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5019410000_-55.0000000000\\\",\\\"662.5019410000_-100.0000000000\\\",\\\"475.0000000000_-100.0000000000\\\",\\\"475.0000000000_-250.1279080000\\\",\\\"445.7613850000_-250.1279080000\\\"]}\"}","{\"color\":\"#519355\",\"startPinId\":\"pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53\",\"rawStartPinId\":\"pin-type-component_317b37d2-20d2-4d51-9e3b-72e93df3ce83_1\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_53\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"520.7613850000_-250.1279095000\\\",\\\"520.7613850000_-115.0000000000\\\",\\\"677.5019245000_-115.0000000000\\\",\\\"677.5019245000_-55.0000000000\\\"]}\"}","{\"color\":\"#ca2424\",\"startPinId\":\"pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54\",\"rawStartPinId\":\"pin-type-component_29b8e01a-285a-4675-b6e8-5a3c24817ccc_1\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_54\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"572.5000000000_-265.0000000000\\\",\\\"572.5000000000_-190.0000000000\\\",\\\"647.5000000000_-190.0000000000\\\",\\\"647.5000000000_-40.0000000000\\\",\\\"662.5019410000_-40.0000000000\\\"]}\"}","{\"color\":\"#3885c1\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55\",\"endPinId\":\"pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_55\",\"rawEndPinId\":\"pin-type-component_d31a6738-5eba-41b7-bcd4-00ce53bb91e4_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5019245000_-40.0000000000\\\",\\\"692.5000000000_-40.0000000000\\\",\\\"692.5000000000_-205.0000000000\\\",\\\"640.7613850000_-205.0000000000\\\",\\\"640.7613850000_-250.1279080000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40\",\"endPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_40\",\"rawEndPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_28_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"362.5002115000_215.0000000000\\\",\\\"362.5002115000_260.0000000000\\\",\\\"460.0000000000_260.0000000000\\\",\\\"460.0000000000_792.5000000000\\\",\\\"557.5000000000_792.5000000000\\\",\\\"557.5000000000_830.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg\",\"endPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_29_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_1_29_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"572.5000000000_1100.0000000000\\\",\\\"610.0000000000_1100.0000000000\\\",\\\"610.0000000000_830.0000000000\\\",\\\"572.5000000000_830.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg\",\"rawStartPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_28_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1067.5000000000_215.0000000000\\\",\\\"1067.5000000000_177.5000000000\\\",\\\"992.5000000000_177.5000000000\\\",\\\"992.5000000000_725.0000000000\\\",\\\"422.5000000000_725.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos\",\"rawStartPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_1\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_27_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1082.5020835000_215.0000000000\\\",\\\"1082.5020835000_162.5000000000\\\",\\\"977.5000000000_162.5000000000\\\",\\\"977.5000000000_710.0000000000\\\",\\\"407.5000000000_710.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos\",\"rawStartPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_2\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_26_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1097.5000000000_215.0000000000\\\",\\\"1097.5000000000_147.5000000000\\\",\\\"962.5000000000_147.5000000000\\\",\\\"962.5000000000_695.0000000000\\\",\\\"407.5000000000_695.0000000000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67\",\"endPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_67\",\"rawEndPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5019245000_50.0000000000\\\",\\\"677.5019245000_57.5000000000\\\",\\\"1112.5000000000_57.5000000000\\\",\\\"1112.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg\",\"rawStartPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_4\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_25_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1127.5020835000_215.0000000000\\\",\\\"1127.5020835000_132.5000000000\\\",\\\"947.5000000000_132.5000000000\\\",\\\"947.5000000000_680.0000000000\\\",\\\"422.5000000000_680.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66\",\"endPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_66\",\"rawEndPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5019410000_50.0000000000\\\",\\\"1142.5000000000_50.0000000000\\\",\\\"1142.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos\",\"rawStartPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_14\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_24_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1277.5020835000_215.0000000000\\\",\\\"1277.5020835000_117.5000000000\\\",\\\"932.5000000000_117.5000000000\\\",\\\"932.5000000000_665.0000000000\\\",\\\"407.5000000000_665.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg\",\"rawStartPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_15\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_23_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1292.5000000000_215.0000000000\\\",\\\"1292.5000000000_102.5000000000\\\",\\\"917.5000000000_102.5000000000\\\",\\\"917.5000000000_650.0000000000\\\",\\\"422.5000000000_650.0000000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65\",\"endPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_65\",\"rawEndPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5019245000_35.0000000000\\\",\\\"677.5019245000_42.5000000000\\\",\\\"1217.5000000000_42.5000000000\\\",\\\"1217.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64\",\"endPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_64\",\"rawEndPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5019410000_35.0000000000\\\",\\\"1232.5020835000_35.0000000000\\\",\\\"1232.5020835000_215.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63\",\"endPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_63\",\"rawEndPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5019245000_20.0000000000\\\",\\\"677.5019245000_27.5000000000\\\",\\\"1247.5000000000_27.5000000000\\\",\\\"1247.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62\",\"endPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_62\",\"rawEndPinId\":\"pin-type-component_fd8f8cb1-e823-496b-ad06-7cf0fbacd90f_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5019410000_20.0000000000\\\",\\\"1262.5000000000_20.0000000000\\\",\\\"1262.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg\",\"rawStartPinId\":\"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_2\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_22_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1127.5000000000_500.0000000000\\\",\\\"1037.5000000000_500.0000000000\\\",\\\"1037.5000000000_635.0000000000\\\",\\\"422.5000000000_635.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos\",\"rawStartPinId\":\"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_1\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_21_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1127.5000000000_515.0000000000\\\",\\\"1022.5000000000_515.0000000000\\\",\\\"1022.5000000000_620.0000000000\\\",\\\"407.5000000000_620.0000000000\\\"]}\"}","{\"color\":\"#dddddd\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8\",\"endPinId\":\"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_8\",\"rawEndPinId\":\"pin-type-component_d1c6c4d4-8ab8-4ab8-a980-754c86362baa_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"407.5001575000_215.0000000000\\\",\\\"407.5001575000_245.0000000000\\\",\\\"475.0000000000_245.0000000000\\\",\\\"475.0000000000_605.0000000000\\\",\\\"1007.5000000000_605.0000000000\\\",\\\"1007.5000000000_530.0000000000\\\",\\\"1127.5000000000_530.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_0_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_19_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"767.5000000000_-175.0000000000\\\",\\\"767.5000000000_-167.5000000000\\\",\\\"872.5000000000_-167.5000000000\\\",\\\"872.5000000000_590.0000000000\\\",\\\"407.5000000000_590.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_3_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_18_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_-175.0000000000\\\",\\\"857.5000000000_-175.0000000000\\\",\\\"857.5000000000_575.0000000000\\\",\\\"422.5000000000_575.0000000000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_8_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_-175.0000000000\\\",\\\"887.5000000000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_9_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_-175.0000000000\\\",\\\"902.5000000000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_10_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"917.5000000000_-175.0000000000\\\",\\\"917.5000000000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_11_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"932.5000000000_-175.0000000000\\\",\\\"932.5000000000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_13_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"962.5000000000_-175.0000000000\\\",\\\"962.5000015000_-175.0000000000\\\",\\\"962.5000015000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_12_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"947.5000000000_-175.0000000000\\\",\\\"947.5000015000_-175.0000000000\\\",\\\"947.5000015000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_14_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_15\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.5000000000_-175.0000000000\\\",\\\"977.5000015000_-175.0000000000\\\",\\\"977.5000015000_-172.9900030000\\\"]}\"}","{\"color\":\"#0023eb\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15\",\"endPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_15_0\",\"rawEndPinId\":\"pin-type-component_22bfc2f4-ec74-4e25-b5ac-80edc339190c_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_-175.0000000000\\\",\\\"992.5000015000_-175.0000000000\\\",\\\"992.5000015000_-172.9900030000\\\"]}\"}","{\"color\":\"#48a1d1\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_1_1_0\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_47\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"782.5000000000_-175.0000000000\\\",\\\"407.5001575000_-175.0000000000\\\",\\\"407.5001575000_-70.0000000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_8_3\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_33\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"887.5000000000_-115.0000000000\\\",\\\"827.5000000000_-115.0000000000\\\",\\\"827.5000000000_-160.0000000000\\\",\\\"353.5002220000_-160.0000000000\\\",\\\"353.5002220000_-70.0000000000\\\"]}\"}","{\"color\":\"#7E2DD2\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_9_2\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_49\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_-100.0000000000\\\",\\\"812.5000000000_-100.0000000000\\\",\\\"812.5000000000_-145.0000000000\\\",\\\"377.5022770000_-145.0000000000\\\",\\\"377.5022770000_-70.0000000000\\\"]}\"}","{\"color\":\"#BDD393\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_14_1\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_48\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.5000000000_-85.0000000000\\\",\\\"797.5000000000_-85.0000000000\\\",\\\"797.5000000000_-130.0000000000\\\",\\\"392.5001755000_-130.0000000000\\\",\\\"392.5001755000_-70.0000000000\\\"]}\"}","{\"color\":\"#ff3232\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10\",\"endPinId\":\"pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_10_0\",\"rawEndPinId\":\"pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"917.5000000000_-70.0000000000\\\",\\\"917.5000000000_5.0000000000\\\",\\\"1075.0000000000_5.0000000000\\\",\\\"1075.0000000000_-250.0000000000\\\",\\\"1112.5000000000_-250.0000000000\\\"]}\"}","{\"color\":\"#1464c8\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13\",\"endPinId\":\"pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_13_0\",\"rawEndPinId\":\"pin-type-component_127fe76f-620d-42d3-bc33-d5252ff1a787_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"962.5000000000_-70.0000000000\\\",\\\"962.5000000000_-2.5000000000\\\",\\\"1090.0000000000_-2.5000000000\\\",\\\"1090.0000000000_-151.1620000000\\\",\\\"1112.5000000000_-151.1620000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11\",\"endPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_11_0\",\"rawEndPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_28_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"932.5000000000_-70.0000000000\\\",\\\"932.5000000000_-25.0000000000\\\",\\\"902.5000000000_-25.0000000000\\\",\\\"902.5000000000_755.0000000000\\\",\\\"640.0000000000_755.0000000000\\\",\\\"640.0000000000_1145.0000000000\\\",\\\"557.5000000000_1145.0000000000\\\",\\\"557.5000000000_1100.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15\",\"endPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_7425f490-20e5-405c-8f1e-bcd16b84ce42_0_15_0\",\"rawEndPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_27_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"992.5000000000_-70.0000000000\\\",\\\"992.5000000000_-17.5000000000\\\",\\\"887.5000000000_-17.5000000000\\\",\\\"887.5000000000_740.0000000000\\\",\\\"625.0000000000_740.0000000000\\\",\\\"625.0000000000_1160.0000000000\\\",\\\"542.5000000000_1160.0000000000\\\",\\\"542.5000000000_1115.0000000000\\\"]}\"}","{\"color\":\"#735348\",\"startPinId\":\"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_9\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_246c73ed-c3aa-4493-99a9-e79818341acd_0_9_2\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_45\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_440.0000000000\\\",\\\"47.5000000000_440.0000000000\\\",\\\"47.5000000000_-100.0000000000\\\",\\\"437.5022065000_-100.0000000000\\\",\\\"437.5022065000_-70.0000000000\\\"]}\"}","{\"color\":\"#735348\",\"startPinId\":\"pin-type-breadboard_246c73ed-c3aa-4493-99a9-e79818341acd_0_13\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_246c73ed-c3aa-4493-99a9-e79818341acd_0_13_2\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_44\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"227.5000000000_500.0000000000\\\",\\\"32.5000000000_500.0000000000\\\",\\\"32.5000000000_-115.0000000000\\\",\\\"452.5021885000_-115.0000000000\\\",\\\"452.5021885000_-70.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9\",\"endPinId\":\"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1\",\"rawStartPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_9\",\"rawEndPinId\":\"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"422.4980575000_215.0000000000\\\",\\\"422.4980575000_237.5000000000\\\",\\\"490.0000000000_237.5000000000\\\",\\\"490.0000000000_387.5000000000\\\",\\\"542.4958405000_387.5000000000\\\",\\\"542.4958405000_365.0041670000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg\",\"rawStartPinId\":\"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_0\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_17_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.5000000000_365.0000000000\\\",\\\"527.5000000000_560.0000000000\\\",\\\"422.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2\",\"endPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos\",\"rawStartPinId\":\"pin-type-component_ea1a6d9b-043c-42f4-95db-9fdb3e699131_2\",\"rawEndPinId\":\"pin-type-power-rail_246c73ed-c3aa-4493-99a9-e79818341acd_1_16_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"557.5093915000_365.0000000000\\\",\\\"557.5093915000_380.0000000000\\\",\\\"557.5000000000_380.0000000000\\\",\\\"557.5000000000_545.0000000000\\\",\\\"407.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_0\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"767.5000000000_815.0000000000\\\",\\\"655.0000000000_815.0000000000\\\",\\\"655.0000000000_1205.0000000000\\\",\\\"-42.5000000000_1205.0000000000\\\",\\\"-42.5000000000_-130.0000000000\\\",\\\"278.5003105000_-130.0000000000\\\",\\\"278.5003105000_-70.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5\",\"endPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_5\",\"rawEndPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_26_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"781.4944090000_921.4738985000\\\",\\\"781.4944090000_1175.0000000000\\\",\\\"527.5000000000_1175.0000000000\\\",\\\"527.5000000000_1100.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4\",\"endPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_4\",\"rawEndPinId\":\"pin-type-power-rail_2622c028-5eeb-487e-a780-ae7d5e5671cc_0_25_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"795.8902765000_920.5741940000\\\",\\\"795.8902765000_1190.0000000000\\\",\\\"512.5000000000_1190.0000000000\\\",\\\"512.5000000000_1115.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_1\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_29\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"767.5000000000_829.4904140000\\\",\\\"670.0000000000_829.4904140000\\\",\\\"670.0000000000_1220.0000000000\\\",\\\"-57.5000000000_1220.0000000000\\\",\\\"-57.5000000000_-145.0000000000\\\",\\\"293.5002925000_-145.0000000000\\\",\\\"293.5002925000_-70.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_2\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_30\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"766.0509640000_842.5317920000\\\",\\\"685.0000000000_842.5317920000\\\",\\\"685.0000000000_1235.0000000000\\\",\\\"-72.5000000000_1235.0000000000\\\",\\\"-72.5000000000_-160.0000000000\\\",\\\"308.5002745000_-160.0000000000\\\",\\\"308.5002745000_-70.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3\",\"endPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_3\",\"rawEndPinId\":\"pin-type-component_802528b6-1c68-4132-8eb3-ef45339a8beb_31\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"766.0509640000_855.5731115000\\\",\\\"700.0000000000_855.5731115000\\\",\\\"700.0000000000_1250.0000000000\\\",\\\"-87.5000000000_1250.0000000000\\\",\\\"-87.5000000000_-175.0000000000\\\",\\\"323.5002565000_-175.0000000000\\\",\\\"323.5002565000_-70.0000000000\\\"]}\"}","{\"color\":\"#1642b2\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6\",\"endPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_6\",\"rawEndPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"844.4762800000_803.6079140000\\\",\\\"844.4762800000_800.0000000000\\\",\\\"917.5000000000_800.0000000000\\\"]}\"}","{\"color\":\"#ef9cdb\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7\",\"endPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_7\",\"rawEndPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"843.5765155000_816.2042525000\\\",\\\"843.5765155000_814.9979165000\\\",\\\"917.5000000000_814.9979165000\\\"]}\"}","{\"color\":\"#cc1212\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10\",\"endPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_10\",\"rawEndPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.6768110000_853.0936220000\\\",\\\"842.6768110000_860.0000000000\\\",\\\"947.5000000000_860.0000000000\\\",\\\"947.5000000000_859.9989590000\\\",\\\"917.5000000000_859.9989590000\\\"]}\"}","{\"color\":\"#f2681c\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9\",\"endPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_9\",\"rawEndPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"843.5765155000_839.5975205000\\\",\\\"917.5000000000_839.5975205000\\\",\\\"917.5000000000_844.9989590000\\\"]}\"}","{\"color\":\"#eed145\",\"startPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8\",\"endPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2\",\"rawStartPinId\":\"pin-type-component_59718622-87ae-47c5-ab64-77f43e28c079_8\",\"rawEndPinId\":\"pin-type-component_e5348ec8-9804-4ec3-98a4-c934e85c4b49_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"843.5765155000_827.9008865000\\\",\\\"843.5765155000_830.0000000000\\\",\\\"850.0000000000_830.0000000000\\\",\\\"850.0000000000_830.0020835000\\\",\\\"917.5000000000_830.0020835000\\\"]}\"}"],"projectDescription":""}PK
     �9s[               jsons/PK
     �9s[ζ�g{  g{     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"28BYJ-48 Stepper Motor","category":["Output"],"userDefined":true,"id":"de09217e-3b73-b82d-0145-70b2df9a4b72","subtypeDescription":"","subtypePic":"27b84e47-6648-4cee-a869-6ff1a6fc12fe.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"21.25000","numDisplayRows":"34.37500","pins":[{"uniquePinIdString":"0","positionMil":"862.48611,62.50694","isAnchorPin":true,"label":"BLUE"},{"uniquePinIdString":"1","positionMil":"962.47222,62.50694","isAnchorPin":false,"label":"PINK"},{"uniquePinIdString":"2","positionMil":"1062.50000,62.50694","isAnchorPin":false,"label":"YELLOW"},{"uniquePinIdString":"3","positionMil":"1162.47917,62.50694","isAnchorPin":false,"label":"ORANGE"},{"uniquePinIdString":"4","positionMil":"1262.47917,62.50694","isAnchorPin":false,"label":"RED"}],"pinType":"wired"},"properties":[],"iconPic":"50196d33-890c-4789-8115-a73c306e50dc.png","componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"28BYJ-48 Motor Driver","category":["User Defined"],"id":"ecbd5bee-2226-4f1c-8fdb-aaff666e8628","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"00941d67-c746-454a-b945-4fddefc776b2.png","iconPic":"ef87c5cc-d843-475d-a868-97060fb00c54.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"10.89860","pins":[{"uniquePinIdString":"0","positionMil":"841.32961,870.15945","isAnchorPin":true,"label":"IN1"},{"uniquePinIdString":"1","positionMil":"744.72685,870.15945","isAnchorPin":false,"label":"IN2"},{"uniquePinIdString":"2","positionMil":"657.78433,879.81969","isAnchorPin":false,"label":"IN3"},{"uniquePinIdString":"3","positionMil":"570.84220,879.81969","isAnchorPin":false,"label":"IN4"},{"uniquePinIdString":"4","positionMil":"137.50165,680.89094","isAnchorPin":false,"label":"Vcc"},{"uniquePinIdString":"5","positionMil":"131.50362,776.86339","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"917.27685,356.98425","isAnchorPin":false,"label":"blue"},{"uniquePinIdString":"7","positionMil":"833.30126,362.98268","isAnchorPin":false,"label":"pink"},{"uniquePinIdString":"8","positionMil":"755.32370,362.98268","isAnchorPin":false,"label":"yellow"},{"uniquePinIdString":"9","positionMil":"677.34614,362.98268","isAnchorPin":false,"label":"orange"},{"uniquePinIdString":"10","positionMil":"587.37213,368.98071","isAnchorPin":false,"label":"red"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"MB102 Breadboard Power Supply Module 3.3V/5V","category":["User Defined"],"userDefined":true,"id":"307d45d2-aa1f-05de-326e-55c453eb206e","subtypeDescription":"","subtypePic":"fd3ac6b5-800b-45c8-a4ce-2476671127d4.png","iconPic":"915d9337-ea3e-4fec-8caa-7acd53f715e1.png","imageLocation":"local_cache","componentVersion":4,"pinInfo":{"numDisplayCols":"12.59843","numDisplayRows":"20.86614","pins":[{"uniquePinIdString":"0","positionMil":"159.37736,1995.85039","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"159.37736,1895.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"559.37736,1995.85039","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"3","positionMil":"559.37736,1895.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"160.37736,203.85039","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"5","positionMil":"160.37736,101.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"558.58118,203.74848","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"7","positionMil":"558.47927,102.64657","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"8","positionMil":"263.37736,1397.85039","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"9","positionMil":"363.37736,1397.85039","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"10","positionMil":"463.37736,1397.85039","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"11","positionMil":"563.37736,1397.85039","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"12","positionMil":"263.37736,1297.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"13","positionMil":"363.37736,1297.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"463.37736,1297.85039","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"15","positionMil":"563.37736,1297.85039","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Arduino Mega 2560","category":["User Defined"],"userDefined":true,"id":"972688b5-e2a3-1d53-e820-bc24d2f5082a","subtypeDescription":"","subtypePic":"b949fd05-6e10-4256-9d1b-e11f1f9900de.png","fqbn":"arduino:avr:mega","iconPic":"01119c27-1bad-421a-afe4-dfb48490a906.png","imageLocation":"local_cache","componentVersion":15,"pinInfo":{"numDisplayCols":"42.49620","numDisplayRows":"20.99812","pins":[{"uniquePinIdString":"0","positionMil":"3149.60741,99.90612","isAnchorPin":true,"label":"A8"},{"uniquePinIdString":"1","positionMil":"3249.60729,99.90612","isAnchorPin":false,"label":"A9"},{"uniquePinIdString":"2","positionMil":"3349.59328,99.90612","isAnchorPin":false,"label":"A10"},{"uniquePinIdString":"3","positionMil":"3449.62094,99.90612","isAnchorPin":false,"label":"A11"},{"uniquePinIdString":"4","positionMil":"3549.62082,99.90612","isAnchorPin":false,"label":"A12"},{"uniquePinIdString":"5","positionMil":"3649.60682,99.90612","isAnchorPin":false,"label":"A13"},{"uniquePinIdString":"6","positionMil":"3749.60670,99.90612","isAnchorPin":false,"label":"A14"},{"uniquePinIdString":"7","positionMil":"3849.59269,99.90612","isAnchorPin":false,"label":"A15"},{"uniquePinIdString":"8","positionMil":"2249.60846,99.90612","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2349.59446,99.90612","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2449.62212,99.90612","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2549.62200,99.90612","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2649.60799,99.90612","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2749.60788,99.90612","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"2849.59387,99.90612","isAnchorPin":false,"label":"A6"},{"uniquePinIdString":"15","positionMil":"2949.62153,99.90612","isAnchorPin":false,"label":"A7"},{"uniquePinIdString":"16","positionMil":"3649.60682,1999.90612","isAnchorPin":false,"label":"D21"},{"uniquePinIdString":"17","positionMil":"3549.62082,1999.90612","isAnchorPin":false,"label":"D20"},{"uniquePinIdString":"18","positionMil":"3449.62094,1999.90612","isAnchorPin":false,"label":"D19"},{"uniquePinIdString":"19","positionMil":"3349.59328,1999.90612","isAnchorPin":false,"label":"D18"},{"uniquePinIdString":"20","positionMil":"3249.60729,1999.90612","isAnchorPin":false,"label":"D17"},{"uniquePinIdString":"21","positionMil":"3149.60741,1999.90612","isAnchorPin":false,"label":"D16"},{"uniquePinIdString":"22","positionMil":"3049.62141,1999.90612","isAnchorPin":false,"label":"D15"},{"uniquePinIdString":"23","positionMil":"2949.62153,1999.90612","isAnchorPin":false,"label":"D14"},{"uniquePinIdString":"24","positionMil":"989.59606,1999.90612","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"25","positionMil":"1089.60983,1999.90612","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"26","positionMil":"1189.60971,1999.90612","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"27","positionMil":"1289.60959,1999.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"28","positionMil":"1389.60948,1999.90612","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"29","positionMil":"1489.60936,1999.90612","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"30","positionMil":"1589.60924,1999.90612","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"31","positionMil":"1689.60912,1999.90612","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"32","positionMil":"1789.60901,1999.90612","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"33","positionMil":"1889.60889,1999.90612","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"34","positionMil":"1349.60952,99.90612","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"35","positionMil":"1449.60941,99.90612","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"36","positionMil":"1549.62318,99.90612","isAnchorPin":false,"label":"RESET"},{"uniquePinIdString":"37","positionMil":"1649.60917,99.90612","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"38","positionMil":"1749.60905,99.90612","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"39","positionMil":"1849.60893,99.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"40","positionMil":"1949.60882,99.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"41","positionMil":"2049.62259,99.90612","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"42","positionMil":"2749.60788,1999.90612","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"43","positionMil":"2649.60799,1999.90612","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"44","positionMil":"2549.62200,1999.90612","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"45","positionMil":"2449.62212,1999.90612","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"46","positionMil":"2349.59446,1999.90612","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"47","positionMil":"2249.60846,1999.90612","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"48","positionMil":"2149.60858,1999.90612","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"49","positionMil":"2049.62259,1999.90612","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"50","positionMil":"3949.62035,1999.90612","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"51","positionMil":"4049.62024,1999.90612","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"52","positionMil":"3949.62035,1899.90612","isAnchorPin":false,"label":"D22"},{"uniquePinIdString":"53","positionMil":"4049.62024,1899.90612","isAnchorPin":false,"label":"D23"},{"uniquePinIdString":"54","positionMil":"3949.62035,1799.90612","isAnchorPin":false,"label":"D24"},{"uniquePinIdString":"55","positionMil":"4049.62024,1799.90612","isAnchorPin":false,"label":"D25"},{"uniquePinIdString":"56","positionMil":"3949.62035,1699.90612","isAnchorPin":false,"label":"D26"},{"uniquePinIdString":"57","positionMil":"4049.62024,1699.90612","isAnchorPin":false,"label":"D27"},{"uniquePinIdString":"58","positionMil":"3949.62035,1599.90612","isAnchorPin":false,"label":"D28"},{"uniquePinIdString":"59","positionMil":"4049.62024,1599.90612","isAnchorPin":false,"label":"D29"},{"uniquePinIdString":"60","positionMil":"3949.62035,1499.90612","isAnchorPin":false,"label":"D30"},{"uniquePinIdString":"61","positionMil":"4049.62024,1499.90612","isAnchorPin":false,"label":"D31"},{"uniquePinIdString":"62","positionMil":"3949.62035,1399.90612","isAnchorPin":false,"label":"D32"},{"uniquePinIdString":"63","positionMil":"4049.62024,1399.90612","isAnchorPin":false,"label":"D33"},{"uniquePinIdString":"64","positionMil":"3949.62035,1299.90612","isAnchorPin":false,"label":"D34"},{"uniquePinIdString":"65","positionMil":"4049.62024,1299.90612","isAnchorPin":false,"label":"D35"},{"uniquePinIdString":"66","positionMil":"3949.62035,1199.90612","isAnchorPin":false,"label":"D36"},{"uniquePinIdString":"67","positionMil":"4049.62024,1199.90612","isAnchorPin":false,"label":"D37"},{"uniquePinIdString":"68","positionMil":"3949.62035,1099.90612","isAnchorPin":false,"label":"D38"},{"uniquePinIdString":"69","positionMil":"4049.62024,1099.90612","isAnchorPin":false,"label":"D39"},{"uniquePinIdString":"70","positionMil":"3949.62035,999.90612","isAnchorPin":false,"label":"D40"},{"uniquePinIdString":"71","positionMil":"4049.62024,999.90612","isAnchorPin":false,"label":"D41"},{"uniquePinIdString":"72","positionMil":"3949.62035,899.90612","isAnchorPin":false,"label":"D42"},{"uniquePinIdString":"73","positionMil":"4049.62024,899.90612","isAnchorPin":false,"label":"D43"},{"uniquePinIdString":"74","positionMil":"3949.62035,799.90612","isAnchorPin":false,"label":"D44"},{"uniquePinIdString":"75","positionMil":"4049.62024,799.90612","isAnchorPin":false,"label":"D45"},{"uniquePinIdString":"76","positionMil":"3949.62035,699.90612","isAnchorPin":false,"label":"D46"},{"uniquePinIdString":"77","positionMil":"4049.62024,699.90612","isAnchorPin":false,"label":"D47"},{"uniquePinIdString":"78","positionMil":"3949.62035,599.90612","isAnchorPin":false,"label":"D48"},{"uniquePinIdString":"79","positionMil":"4049.62024,599.90612","isAnchorPin":false,"label":"D49"},{"uniquePinIdString":"80","positionMil":"3949.62035,499.90612","isAnchorPin":false,"label":"D50"},{"uniquePinIdString":"81","positionMil":"4049.62024,499.90612","isAnchorPin":false,"label":"D51"},{"uniquePinIdString":"82","positionMil":"3949.62035,399.90612","isAnchorPin":false,"label":"D52"},{"uniquePinIdString":"83","positionMil":"4049.62024,399.90612","isAnchorPin":false,"label":"D53"},{"uniquePinIdString":"84","positionMil":"3949.62035,299.90612","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"85","positionMil":"4049.62024,299.90612","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/05e0cc9a-68eb-4905-ae12-aaf8623b6ed7.svg","propertiesV2":[]},{"subtypeName":"LED Two Pin (Red)","category":["User Defined"],"id":"5f0a7f7f-5908-4e39-94d8-2714a0462581","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"3d0a314b-f708-4b2c-819f-35c414b123ec.png","iconPic":"6608fa58-7afa-4488-b64c-2b761d69d6bd.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/a9e23d57-c0ac-465e-ae7a-a15cecbcb7b3.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"4.24452","numDisplayRows":"5.30565","pins":[{"uniquePinIdString":"0","positionMil":"161.90689,79.96916","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"261.90689,79.96916","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"LED Two Pin (Blue) ","category":["User Defined"],"id":"117aab52-1b06-40f5-98b6-df63a601b0e6","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"2c98734f-75db-43ce-800c-ea69461525e8.png","iconPic":"d4c851cf-9fb5-43cd-809f-e1699313b4d2.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/1f9f88e9-950f-4940-ab85-21b1c84421ad.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33334","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33371","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18643","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"LED Two Pin (Green)","category":["User Defined"],"id":"a70bb5a8-99ed-4f1b-882e-eac0873b75ef","componentVersion":5,"userDefined":true,"subtypeDescription":"","subtypePic":"f9728bc6-2422-4ead-9082-90351081a874.png","iconPic":"9ba3df0f-d630-43f7-8169-617793654d93.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/3749fe76-cef7-4b42-9f27-525b8a44301e.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33333","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33333","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18606","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"LED Two Pin (Yellow) ","category":["User Defined"],"id":"1310de1e-180e-4aed-a1c6-f80032a2bfde","componentVersion":4,"userDefined":true,"subtypeDescription":"","subtypePic":"42e39361-2f02-4030-a678-a3271aadd3f6.png","iconPic":"a4af1710-95e2-4b5e-9600-8e4d90487313.png","hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/e51a5bd5-4abe-4a22-abdb-307c464150b2.svg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"8.33334","pins":[{"uniquePinIdString":"0","positionMil":"266.66667,133.33359","isAnchorPin":true,"label":"Cathode"},{"uniquePinIdString":"1","positionMil":"421.74257,134.18631","isAnchorPin":false,"label":"Anode"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"DC Gear Motor (3-6V)","category":["User Defined"],"userDefined":true,"id":"7115dd0c-9076-1603-96e1-f4f66aa483df","subtypeDescription":"","subtypePic":"e2e2c934-b375-45fc-834c-534243cbf361.png","iconPic":"6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png","imageLocation":"local_cache","componentVersion":7,"pinInfo":{"numDisplayCols":"26.87010","numDisplayRows":"12.94650","pins":[{"uniquePinIdString":"0","positionMil":"119.68733,976.07429","isAnchorPin":true,"label":"V+"},{"uniquePinIdString":"1","positionMil":"119.68733,317.15429","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/7f9ce5f4-cc5c-40e6-be98-a947128d0a84.svg","propertiesV2":[]},{"subtypeName":"Rotary Potentiometer","category":["Input"],"userDefined":false,"id":"7013093c-3557-9fba-53d2-85a05ece47f1","subtypeDescription":"","subtypePic":"028dc4b4-5e34-49e4-81aa-ecc68ea503ed.png","pinInfo":{"numDisplayCols":"4.05403","numDisplayRows":"8.29847","pins":[{"uniquePinIdString":"0","positionMil":"103.01395,7.75694","isAnchorPin":true,"label":"leg1"},{"uniquePinIdString":"1","positionMil":"202.98622,7.72916","isAnchorPin":false,"label":"wiper"},{"uniquePinIdString":"2","positionMil":"303.07656,7.75694","isAnchorPin":false,"label":"leg2"}],"pinType":"wired"},"properties":[{"type":"dropdown","name":"Resistance","value":"10000","options":["1000","10000","50000","100000"],"showOnComp":false,"required":true}],"iconPic":"06c5fde6-b2c8-47bb-9830-971f0c5559bd.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"LCD Display (16 pin)","category":["User Defined"],"userDefined":true,"id":"23598c1c-7607-4538-b177-9ab948fb1937","subtypeDescription":"","subtypePic":"31959ea2-aec5-42cb-a646-ec7cb3b6e41e.png","pinInfo":{"numDisplayCols":"31.57611","numDisplayRows":"14.25319","pins":[{"uniquePinIdString":"0","positionMil":"318.95833,1322.88889","isAnchorPin":true,"label":"VSS"},{"uniquePinIdString":"1","positionMil":"418.97222,1322.88889","isAnchorPin":false,"label":"VDD"},{"uniquePinIdString":"2","positionMil":"518.95833,1322.88889","isAnchorPin":false,"label":"VO"},{"uniquePinIdString":"3","positionMil":"618.95833,1322.88889","isAnchorPin":false,"label":"RS"},{"uniquePinIdString":"4","positionMil":"718.97222,1322.88889","isAnchorPin":false,"label":"R_W"},{"uniquePinIdString":"5","positionMil":"818.95833,1322.88889","isAnchorPin":false,"label":"E"},{"uniquePinIdString":"6","positionMil":"918.97222,1322.88889","isAnchorPin":false,"label":"DB0"},{"uniquePinIdString":"7","positionMil":"1018.95833,1322.88889","isAnchorPin":false,"label":"DB1"},{"uniquePinIdString":"8","positionMil":"1118.95833,1322.88889","isAnchorPin":false,"label":"DB2"},{"uniquePinIdString":"9","positionMil":"1218.95833,1322.88889","isAnchorPin":false,"label":"DB3"},{"uniquePinIdString":"10","positionMil":"1318.95833,1322.88889","isAnchorPin":false,"label":"DB4"},{"uniquePinIdString":"11","positionMil":"1418.97222,1322.88889","isAnchorPin":false,"label":"DB5"},{"uniquePinIdString":"12","positionMil":"1518.95833,1322.88889","isAnchorPin":false,"label":"DB6"},{"uniquePinIdString":"13","positionMil":"1618.95833,1322.88889","isAnchorPin":false,"label":"DB7"},{"uniquePinIdString":"14","positionMil":"1718.97222,1322.88889","isAnchorPin":false,"label":"A"},{"uniquePinIdString":"15","positionMil":"1818.95833,1322.88889","isAnchorPin":false,"label":"K"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"181","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"ce527fa2-4558-4370-a5e7-21077342728a.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Pushbutton","category":["User Defined"],"userDefined":true,"id":"232ac546-6e45-4194-9a27-0fa614949a21","subtypeDescription":"","subtypePic":"e2a053a3-24a6-43e1-ac97-395cbc045e87.png","pinInfo":{"numDisplayCols":"2.45180","numDisplayRows":"3.30020","pins":[{"uniquePinIdString":"0","positionMil":"221.06000,315.00000","isAnchorPin":true,"label":"Pin 3 (out)"},{"uniquePinIdString":"1","positionMil":"221.06000,15.00000","isAnchorPin":false,"label":"Pin 4 (out)"},{"uniquePinIdString":"2","positionMil":"21.06000,315.00000","isAnchorPin":false,"label":"Pin 1 (in)"},{"uniquePinIdString":"3","positionMil":"21.06000,15.00000","isAnchorPin":false,"label":"Pin 2 (in)"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"PTS645SL50-2 LFS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"C&K Components","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"6b551873-9f16-48c5-b1b9-2fc6ab10f815.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Pushbutton","category":["User Defined"],"userDefined":true,"id":"232ac546-6e45-4194-9a27-0fa614949a21","subtypeDescription":"","subtypePic":"e2a053a3-24a6-43e1-ac97-395cbc045e87.png","pinInfo":{"numDisplayCols":"2.45180","numDisplayRows":"3.30020","pins":[{"uniquePinIdString":"0","positionMil":"221.06000,315.00000","isAnchorPin":true,"label":"Pin 3 (out)"},{"uniquePinIdString":"1","positionMil":"221.06000,15.00000","isAnchorPin":false,"label":"Pin 4 (out)"},{"uniquePinIdString":"2","positionMil":"21.06000,315.00000","isAnchorPin":false,"label":"Pin 1 (in)"},{"uniquePinIdString":"3","positionMil":"21.06000,15.00000","isAnchorPin":false,"label":"Pin 2 (in)"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"PTS645SL50-2 LFS","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"C&K Components","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"6b551873-9f16-48c5-b1b9-2fc6ab10f815.png","componentVersion":3,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Water Level Sensor","category":["Input"],"userDefined":false,"id":"97784b10-4dcd-a3be-9167-75f1272c8490","subtypeDescription":"","subtypePic":"0657d52a-d145-430e-bb7e-5d1be0618b5b.png","pinInfo":{"numDisplayCols":"7.873610000","numDisplayRows":"24.409700000","pins":[{"uniquePinIdString":"0","positionMil":"278.9027,2373.2617","isAnchorPin":true,"label":"SIG"},{"uniquePinIdString":"1","positionMil":"378.9027,2373.2617","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"478.9027,2373.2617","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"iconPic":"8ade0660-1c92-4b58-a3e7-adda420d3982.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"L293D H-Bridge","category":["User Defined"],"userDefined":true,"id":"155f7657-2d2d-eaf2-280f-5c76a41d0679","subtypeDescription":"","subtypePic":"022fab5a-d187-48c2-96d7-20ad2a5d1671.png","iconPic":"39d025b2-988a-45cd-b457-87e73cc458ec.png","imageLocation":"local_cache","componentVersion":1,"pinInfo":{"numDisplayCols":"8.00000","numDisplayRows":"3.30000","pins":[{"uniquePinIdString":"0","positionMil":"50.00000,21.69999","isAnchorPin":true,"label":"Enable 1"},{"uniquePinIdString":"1","positionMil":"50.00000,308.30001","isAnchorPin":false,"label":"+V"},{"uniquePinIdString":"2","positionMil":"750.00001,21.69999","isAnchorPin":false,"label":"+Vmotor"},{"uniquePinIdString":"3","positionMil":"750.00001,308.30001","isAnchorPin":false,"label":"Enable 2"},{"uniquePinIdString":"4","positionMil":"150.00000,21.69999","isAnchorPin":false,"label":"In 1"},{"uniquePinIdString":"5","positionMil":"150.00000,308.30001","isAnchorPin":false,"label":"In 4"},{"uniquePinIdString":"6","positionMil":"250.00000,21.69999","isAnchorPin":false,"label":"Out 1 ( Controlled by Enable 1 )"},{"uniquePinIdString":"7","positionMil":"250.00000,308.30001","isAnchorPin":false,"label":"Out 4 ( Controlled by Enable 2 )"},{"uniquePinIdString":"8","positionMil":"350.00000,21.69999","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"9","positionMil":"350.00000,308.30001","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"10","positionMil":"450.00001,21.69999","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"11","positionMil":"450.00001,308.30001","isAnchorPin":false,"label":"0V"},{"uniquePinIdString":"12","positionMil":"550.00001,21.69999","isAnchorPin":false,"label":"Out 2 ( Controlled by Enable 1 )"},{"uniquePinIdString":"13","positionMil":"550.00001,308.30001","isAnchorPin":false,"label":"Out 3 ( Controlled by Enable 2 )"},{"uniquePinIdString":"14","positionMil":"650.00001,21.69999","isAnchorPin":false,"label":"In 2"},{"uniquePinIdString":"15","positionMil":"650.00001,308.30001","isAnchorPin":false,"label":"In 3"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"DHT11 Humitidy and Temperature Sensor","category":["User Defined"],"userDefined":true,"id":"a76bb123-3d3c-417d-b1f3-c8417efb7bc7","subtypeDescription":"","subtypePic":"779eddd4-9cc6-4216-b155-89a4f50be07b.png","iconPic":"44e1934a-57d6-434e-9b76-9cc9cf9f98cc.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"7.00000","numDisplayRows":"10.00000","pins":[{"uniquePinIdString":"0","positionMil":"200.00001,100.00056","isAnchorPin":true,"label":"VDD"},{"uniquePinIdString":"1","positionMil":"300.00001,100.00056","isAnchorPin":false,"label":"DATA"},{"uniquePinIdString":"2","positionMil":"400.00001,100.00056","isAnchorPin":false,"label":"NULL"},{"uniquePinIdString":"3","positionMil":"500.00001,100.00056","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"componentVersion":1,"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Resistor","category":["User Defined"],"id":"1c569fa1-772b-452c-b113-493dd976b9c0","subtypeDescription":"","subtypePic":"b01488b3-8551-4b4c-b09f-2812c4acc168.png","userDefined":true,"componentClass":"resistor","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[],"iconPic":"d3b73945-fe79-451b-b309-b64aab767520.png","componentVersion":7,"imageLocation":"local_cache","propertiesV2":[{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"200","displayFormat":"input","showOnComp":true},{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.1%","value":"0.1%"},{"label":"0.25%","value":"0.25%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false},{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"integer","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false}],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �9s[               images/PK
     �9s[������  ��  /   images/27b84e47-6648-4cee-a869-6ff1a6fc12fe.png�PNG

   IHDR  �  R   ���P   	pHYs  H_  H_#�
{   tEXtSoftware www.inkscape.org��<    IDATx���yx�y&�������7 ���)�(j�6[�6Ӣe��H^�ǎ3��s�L�sg�vnf�8�d2I�+�"�Z���H�i9�lI�H�%�;A�@��ݵtm�	��H�]]������1��h6��s��	�낈������*K�t DDDDDDD���������*0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
0A'""""""�LЉ������� t""""""�*���������
�* Q#۴i�"BD��� !˲� "�PHq'!B�q��(������+��A� 
������EQ4]�5EQ�[��0B�P�u]˶����ի�`��DDD�a�u+Q�{���'��8�u�	��LEq��M��6	���I���}���q_B�u�!A�Ar]w����s�(�'A�w���U��+4Q�c�NDDt�>�l�$Im��L���s�;�q�ɂ L0ܕf�w]��(�']�=��c��p�u�c��{o��aU/&�DD��^z饴asA�#�\�ug�$� f �W8�zS p�Q�u��`�$I��ٷjժ�ʆGDDT9LЉ���;�P�� �ug� s����o�� ����_�}���$��������Z��#""
t""�===r*����"�q���b �H��w�u�] zEQ��7�n���������LЉ��&���SLӼV�� ���{� 3���Ƙ��� �%I�[�(�u�]w��t`DDD�b�NDDU��g��-I�
 #��r �*U�S� ��- oٶ���{�=P須��.�	:U�g�y&)��2�qV�p���X鸨.d]�}�+� l�e��;�c��A�`�NDD�$����\׽�uݕ n� �XḨ18 v��_����=��Ӌ��扈��t""3===R*�Zp.!��� ��t\D�v]�uA^�	&�jŊf��""�������y�搦i�����V �J�ET�! �.�ˎ�\(�loo�+�'&�DD�^xa��8w���������<� �o~8������.i�uݟxQ�W�Z���Q�`�NDDey�Z��8��\׽K�Y���.�yz��j������b	�H�߀���u_��?���{3����jt""*�s�=w� �X�z R�C
̥�l~~^���H�mA~�8�&Q���'>���Qma�NDD���'�L&?�� ����1�e�s����:?iYy������
��)�����o�+U7&�DDtQ�<�̤p8|ή��	@�pHe9?I�X�.��^�	|A����
�����OW: ""�>LЉ�h���??M�ϸ�� �����$��M�����M�m � �m�O�^��x�""�������=��s3 �/B;���L��d���8���n��O~�{*Ut"����x��8�AX��J�s%�O���EW�FWڷ�h�v��ի�T:""[LЉ�ĳ�>�,��\��� w��W���=?���O֫=ia��8?�B�<�ND���ձ͛7't]��u�� ��tL��q��Ye7]��7 �P��ﾻP逈�(LЉ���7���ꫯ��eY_N$נʪ����8?��ڌ$�U��\�}R�G��_���_����C���V0A'"�O?��"�0�a��b��&M�(���+�T�ޟ�WSҞ��2�㼒L&���{��Y�x���|LЉ�j��͛�gΜ�=�0~�0���OO�ӈ���m$)��՛jXaw]}}}p]�  ���D"��?���~����FDDea�NDT��zꩻu]��b�x�i���U.�2Ə?&11!�FT�d]�4d2�|_�$'��
��졇�ɘEDDec�NDT#6mڤ
����/��9�J߿'N��P���p�oY�g	х��N�`�e�L4̈́��d2��U�V��	:Q�{�'�/����i�9�S��d2�d2�K,#��@#��ju�q���]�$�	�ÿ�D"��C��k0DD�+&�DDUh��͡����d���>���jI�0i�$��u��|~&�\�\���H$rZ��oO�8�oo��v��`���WLЉ���/�В�f�i���bԯyǏY����3)'
�H�����ӧaY����p،D"�&�����'?y���DD(&�DDU����V۶��0�,����j<G:���g4��(ue�X,�̙3�]_�$W��-�X�wx���|����<a�NDT9��?���}�0���^H�����$�+�D���D�R	���TU�ڑH�t$���z�; ��@DTLЉ��XOO�,�_��[��'����͈�bLʉj��V�]�ũS�/�(�rA��E�����@/FDD`�ND4FzzzҎ���akMӼ��>E�dѨo�ډh���n��ڡPȌF�=�ƍ��w�ygv�.LD����lӦMS��w���i��X^[�e(�Y���LD��,�B����uC���F�L&���O~��^����0A'"
ȳ�>�$���O]�o�m{̲�P(�X,�h4�J4U/�u��:4M�i�cv�s��H$�~�}���5&�DD>{���o�u�_�X2Vﱂ �&��pxL�ID�gY4M��끟M!���.I���v��_��E��t""�<��S+
��w�X6Vﭲ,#�!�p;Qs�b���٪���{B�Я����E�����'��V���u}�X���k��x<�P(��������k�6&�έ���(������ Qc�ND�ѦM�������i���Z*�"EA,��r"�P���0
ض��έ����֭{3��!&�DD%z������k�v�X��r;��0���b1���#g�����O��o~A"�:����
=��S3UU��a�8�h�,��h�7nc'"�ضMӠ�j����%�[EY{�����bDDu�	:чx��'���C]�?t�4Q���"���8t]����oEэD"?7n�g���@/FDT㘠]���?��r��4틖eIA^+
AQD�Qnc'�1�.��"��<,�
�Z�PȎ�b��d�˫V�2�Q�b�NDt7n�C]���4�h��	�B�+�DD�4RP.�6m�p��(��=��C_�Q"��0A'":Ϗ~��v]���0��A^G�e��qȲ�e��Jf�&TU���^'�b��noo�a�""�!LЉ� ����0M�S��yA�/F�Q(��p8�5���`�6
�t]��ܹBr�#�Ⱥ|��و��1A'����3�L)
ݚ���(��Qͱ,k��{PA��(�(���}��w*�U9&�DԐ��o�.��B���	,k�F�H&�L̉��9��B� M�[Q�$ɎF�������׿�u'��U1&�D�p���?S,�[,���F4E<gs"�;c�����\$�͵k�n�DDU�	:5�'�xb�aOh��,������hW6"��9��iZ ���H$��������r"�*������͛C�O���B�𥠶���5*۶�����.I��(ʏ�����?���t"�k���_6�ۦi*A��s"���N���p!��փ>��@.@DT��Q]���iYֳ�a,
b~Y��H$�bND�>�e!�ˡX,�>���� ���>����*�	:����������Alg�$	��@QY�'"��a ����m��E�Q�׮]�;�ONDTALЉ�n����T,��u}��s���x<�X,A�����.��]ב���8�wM�ey �L>t���o�}r"�
`�ND5���WޱcG����	�=-�#�31'"��q��
UU}o�&E��$I�joo��<�a�ND5����aM���4͘�s�b1$	�b �߉|%IA��8��T��u]��y������pX���_|��7�>9�a�ND5���'mY�&M�n��},
!�N#
�:/�刢�H$Y�!�2"���0dY�$I�B��=8�m��², @�X�eY0M�i�~mt]�i�c��$\!9A��~�8��Gyd��ɉ�� t"�96l��i~۶m��yEQD"�@,��b<ѨH$�X,EQ��FU�#�m��u�a@Ӵ��Ț�qE�c���}��B�b4�Ok׮�G_'&"
t"�O>��B��c�0��s�s+.�����N�iǗH$�J���!IR��*�뺣�z�P@.�C>���15.�qP(����v477߹jժ~�''"
 t"�	7n�u]׿c�����,#�J�\�D�)����	�t�d���˵j8��|>���a�r9�J�KP��%I2E��5k�����	:U��}�{�X,�cUUo�s^I��L&�D���L8M���tþ�\�E.�C&����
�B�C���:r�����A@4}�����U�V�l:U-&�DT���5�|���eE��S��q(�¶i�I4EKKZZZ�L&�:��4��d088�L&���T����|��yeY�B���֯_�����	:U�-[�������w_�p8�T*���T�X,�q��aܸq�����ض���A`hh��$�eaxx��.����lٲ{-Z��~z"�21A'�����u�a�۲��_s
��D"EQ����$I?~<&N��d2Y�p�eYD?��l�á�ir����1dY�F������ܷI������������M�qǷ=ÑH�d�E����d2�	&`	�� ]���ߏӧO�0�J�C5�u]C�u����D"y���6)Q��Q�����2��aL�kN�4�RH��I�&���Ѩo%�
���L&���>U:�A��e�x8�uݺu�|����&�DTQ===_QU�X�����h4�d2��O�P�h�&M¤I�X��
躎�'O�ԩS<�N�D�tI��X,�;k׮���MJDT"&�DT�7o�<y�9M����}(
!�J!�2կT*�)S�����Uث�i����C__�������Eöm_��,�\Uջ����GDc�	:�����kt]�I�Xl�kNEQXȋ>T*����ӑJ�*
]�q��ׇ�Ǐ3Q�Kr]�B�B��9eY�B_�~��&%"�LЉhLmܸ�
�?wǗ��("�J!��1թt:�����O�]ׅa�u}�u]�i��,���gY\�E(� ���("
!�@��~)��X,V��A��ɓ'q��	&�tI~�����(��k���/]&�D4&}��h8~I��[��3�"���աj]1w�|~tկP( ��C�4_�H]�H$2��'	$�I$	Ȳ<�\�mۣ���P��M�D"ۛ��n^�z��]t"
\GG��e�d��/{йjN&�bƌ7n\�C��PU�l�l��þ�s�H��t:���&���hYhY�9�S�N����4��@6����
���d����g��2!�%0A'�@uww�����կ-�H�t����$I´i�0y��n�VU���`ݬ���ojjBKKZZZ*��k��C�!��T,�^�� ����7]E'�}uݺu��eB"��`�NDA;;;��4�S~�ό$�kN#&M������T�wgΜA?}K��(�hjj¸q�0~�x$���144��BӴ�\����i����S�P(���v���	:����k�eY�4c���a455U}!+�EQ0gΜ1��oY���q��i�9s�}��b1���b�ĉc~��q?~Ǐ�}�m�F�X�e>Y�O���׭[wԗ	���a�ND����y@U�n˲|Yƌ��[���&�"���0eʔ1;��8p��q0�EQ0i�$�����ϰ�iؿ?�����TF�A��y_�$�L&�k|���|���LЉ�G������:�Sv�$IR�T�U���N�1g�D��1�^.�É'�����
\#I�Ә:u*Z[[�����S�p���9�O��� P��׭[�{>�FD�������#�ş��Bm�rt5T���"�"fΜ�������8�h�����^#�$	���hkk�#	�b{��E6��ZT[����0��e�h4�KY�?����'xDT&�DT���������4Ͳ�Y	��x<�x<�GhTgE��y�}�E?~ǎk�bo���Ԅ�ӧc�ĉ�Q8u�<�#	������P��3�$�����!4"jPLЉȳ���{u]Ҷ�ϛK��t:]�
�T�A��)S���h�@UUq��A���1�C��`���:uj����B{���]�j�i��f��ly�$ɌF��[��YB#����<����sM��o?ΛG"�R)Vi��Ø?~��UUŁ�����*y#�2f͚�iӦ�^���C����3]E7�������ChD�`��Q�:::�4�3�����t9�T
���lWE�PM��YX=dY����1cƌ����~�߿�;%����.b��s�ׯ�קЈ�A0A'�+����G��u}i�s�J;]��ɓ1s��@�&�E�۷'N�`b^Ţ�(�Ν����@^���w�a�� ˲044�˖�h4�N:�^�z�j�� �+����HOO�t]׷�Ų��ɲ�T*�*���$aΜ9?~��s;��Ç�СCl�UC��$�ϟ���f��m��������sSms�l֗���pxP���֭;T~dDTчڸq㝚�=kYV��݊��I{%�=�H.��(��}��I�۷���5lҤI�7o^ Gb�9�cǎ�>/�6�uQ(P(ʞ+
c�ؽk֬yɇЈ��1A'������MUU��8NY�AA@*�B4�+4�#�x.�����6f���Q1k�,̜9����gΜ�޽{y�>�0d�ٲ_�(��D�?���ۧЈ�1A'�K����UU�\�<�$���	�Pȏ���455a����ypǎþ}�|9GJ�%�Lb�H�Ӿ�;<<�w�}�i�:/�>۶��d�~?����u����O�Q�a�ND��������;[���Q.�͢���|޷9������6̝;�ׇ;��a���<A�.��,�({�H$���~�����&�Dt���+���0�%���ǑH$���Ќ30u�T��s��C��M��(��%K����n�&v��Ue�m��|>�˹�H$�}����}��_g�J"���F=��M�Ph�aegM�t����fϞ���V���4;w���АosR�3g���ٳ}ۭcYv�ލ\.��|T_t]G6�-{�H$r<�H,������ED ���9�ڨm/�M��#�"�����
�� �;w.&L��ۜǎÞ={x֜�N��d��:ض�ݻwcxxؗ��������!8�S�<�px8
-����0&�D����|>�s˲"��#I����ߜ.JE̛7�ƍ�e>۶��ۋ��>_�� I/^�I�&�2��8سg}���m��e��K]�$#�����u�B#�����uww߭����e�Ub=� �N�Z��(��?>���}�OUUl۶͗s�T�f͚�9s����8�}�]d2"�z��f�.,(I��(�k֬��>�ED5�	:Q��������+�ǹ�(H$L��A��y�0~�x_�����Ν;�^�����܌����,�=��8����vw�(�uQ(�~h(����~cݺu��ShDTc��5����?�4�o�y�d�X��Ȩ�̛7Ϸ3�{��šC�|��C4�5�\�d2Y�\#�*X8�.EӴ����*��׭[�w>�ED5�	:Q�����B����!���|Y���5s�LL�2��yFV/O�<�CT�h$I�ҥK}yPd�6v����tI�b�l���q�  �s�ڵe}VQ�a�N�`�������o���J�t%��s^,�}�v�P����`ڴie�e�&v��	M�|���eY*����(��~��_��/    IDAT�),"�LЉHgg�UU�l9s�R;]���V̞=��yTU�֭[��of̘������yt]��o��4}����8�#I߰~���>���v0A'j���O���@9s��a455A˪)Gu���,(�h`>��֭[a�O��5y�d,^�ؗ��Ν;��M��u]d2���(������W�U1&�D����9M�V�3ۨѕPK�.-{����0�n���I
̄	p��W���qpp��.x?E��.��l�c��O~��;|
�������\WW�K�&��hMMML��dY��N�3��l�����ߏ�۷�����҂3f�գ����v<�4��=��/|
���WЉꗰaÆWu]_Y�$�x�D¯��N����K�"��5��� �m��-�4f���q�ז����~�:uʧ��^����; D���y�}
���WЉꓰaÆ7�MΓ�$�s�"s��);9�eE���Lo��Vٯ�Y�f���>T"�@2�,k]�oذa��B"�*�����=��[���(g�t:EQ����Xkkk���s��z뭲�y188�;v�u�\E̟?��'�C)�R��1]ׯ}�Ƕ�U	&�Du����U�0��3G:�F4�+$�c�D3g�,k�|>�-[���,�"򠿿o��vYIz$�UW]�z���(�j�򎎎7}��� t�:�aÆW4M+k[{SS�s�"�p���/�쮦i,GU�ԩSx�wʚ#�N���ͧ������k������U�"�
c�NT':::~����^�����D"?â:6o޼�^/�ib�֭(�>FET�cǎ�СCe�1m�4��i���D���T���������B"�
c�NT:;;�i�G��ió�t�&O�\�M��8رcTU�1*"�ݻ'O�,k�y���=���,�hnn.k%]UՏwtt���aQ�0A'�qO��z��� ����,��1EQ�����ۋ��A�""�_oo/���<��es���1"�g#Iz�G�����x�ǰ����հ���nM�>�u�(�hii�*]1Q1o޼�n"���_��$Q�����ۡi��9ZZZ��p@�#���������cXD4Ƙ�ը�����P(��:^�$��� 
�չ������������>FD�b���۷��#}���,�IW,
�����$�����Q��"�����uvv�wM�~��xI����I�|���]2�Ĕ)S<��4;w��1"���r9�޽��xI�0w�\#�z7� ��$]U�/tvv���a�a�NTc����HӴ��:^E&�T2A0{�l�E�F�±�9բ'N�رc�ǧR)L�8�ǈ������AWW�W}��� t�����EUU�庮��#�ڙ�S��N�Z�����^��m�0M�_�mW:�������1c�}PI�H�5M�����/�L�z�ODc�����B���m۞>�EQd+5�$�b���W�O�8�]�v�U��m�\�\�B��B�uh��4Q,/{6:C�eD"D"����_MMM�����(X�r�燜���ػw��QQ��,�L�s-Q�x<��5k�<�shD &�D5�G?����|�e۶=�
���p���ŋ�N�=��4���/���C���\.���d2�P( ���D���MMMH��|�w�N��E�y_n�6jL�i"��x~OEщ�bw�[�n����ߘ�U�'�|ra6��n۶�;�>��&/&L��y��y�.�|�M&#�`�&���p��i�>}�a�4^���, �pg�^tḀf���.ƍ���VL�2���4��,[���r]ױm۶�*�Sc*��f��_;�P��J��>��{|��|����=������b���2��9�CE,_��H���`���>GU�L�ĉ'p��q���_v5,*��,��E��f-)鸈椈X�×?r�@^sP�\d.���qj����6
��?�S�&O��ɓ'�����߷^ɲ��+Wz��8|�0�?�sT�������dr�<p��Ј�'LЉ�ԦM�����æi��2~� ϙ�Wmmmhkk�4vxxo��W	qv'A?�=�'N\��۸����$�laz��I�<��"����q䔅c�m>eúD}�T*�ٳg����E&�?~<�/_�i�m�غu+L��9*j�bCCC�������X,6���]�94"��U'1���`rN�"�2�N��i�����m��ܶm=z�h�oI�Na�0�ja\jl��K��qͼ�;l���a�Z�=dB=o�}xx۶mî]���ֆY�f!�L�i���̙3���Ckkk�c%IB[[8@dT�dYF:��||�4�	�(n0��Ȉ�\A'�B6l�w]�o�:>�N#��5�y��a	��>|{�4�G�4q��A�۷�b��&���!\�@��Y!�".���v\<ac�A[���.�W�Ǐ����R�(+O�e�t�M������۷CU� "�F`FY5>b��O~��;|��|����tuu�s�P�u���$�;QY��.]ꩭ��ix����m�طo������<��X�D���h��rY��m�L�����}V����X�hQî��S�=��`���>GD�DUU�r9��E�����{�� "�1A'�"���R(��?��D�x�稨�,X����[o��3g��Q�;|�0v��]�/����>zM��!$U�jy)���xeGo�5aZ�O	���ӧc��{��Css���;w���+���Q(<�O&��f͚��1$"*t�*����|>���8���c�R���aQ����X�l������ضm��U�L&�m۶!��^��i$�}C�f�-�V)9�ŋo�xmW��$	s������!���S��D+W����$��b׮]DE�dxx���(���(��]�v��a�LЉ���O>�pxxx�eY�
7F�Q�R)O7�D�[�p���@�q��k�5�yZ�4�{�����,�ޛ"X<�>���:x��:��3q��D<�5�\㹎A-Z�`��\E'?�0OcC���(ʲ���^��"�1A'��6�l�>j����oY�������V��y#�;s��n�z��%*��#�ui�p<j�O��!��p��̙3�x�b�B��4F�e�r�-���\E'�d2����R�p8
�f<�����"���'&Qu���59�BH��L��ӧO�4�X,����>GS}���ݻ�w����b���n�"k���#�l�l�����C��	�p����uq��A�����CSSS��T�XġC�0w�ܒǦ�i�R)��S���42�,���?�>�i&A�`���ITA\A'������k��/c%IBKKKC�����z��;���ѣ>GT]4M�믿�L潅�椈���0z�=�>x��O��=d"p��2n�:%*@7\<�_���^E,]��fͪ`��E7�|3b�X�c��������T>۶��d<wӈF��y䑏�]!&�D�aÆ��u�w���ƍ�$I~�Ej�ܹ�8qb��t]�+��ǩ�Ŗ��~�����\~���n�!Zz��������GO�hI��m����d����u��Ɵj�Pokkòe��z���ɓ�d�Oc�m��0u(X�e!��x~o����Y�n��{"*t�
����\.���ן���&D"���F�q�u�y:*�{�n;v,�������c�����a~4��4Nfn��[{��ɖ"Ngl����,�*I��k&��x��T�;��v���f�x�uێM�|��P�䱧N�������Q�X�`�O�����֬Y�!�`�N4ƞ~��E�Lf�m۞���ɤ�?�K�1c�N�Z�8M��ꫯ����Ν;�o߾ѯ�7I��U1L�;W����w��.fM��+"X8#TR�z��M���2F+�+���+W�mkH����`˖-0M���0��4�sm�P(dE�ѫ׮]��簈�2���������i'L��T-)�#�H�50Q�b�
�����������DUY��`�֭��?=��"�[�s��Wwxy����̜\ރ���Lt������w��a�t�Mhii�#�R�*��#G�zW
��\.���,�YMӦ|�+_���1R�����P�X|�kr�F����&L��)9�u'O� ��ro��&N�81���h�=V�����b��_�2a;.��'�c+d����c`��0��"��l9Յi�x�W�r�ʺ�>R�~���%�mmm������K2���8�u���b1�H$^���Ȉ�b��N4F���-
_�26�������wW_}��?{��šC����l��믿�S�N�~��"���<+=�x�����uO᐀�q����<��:�_O00|�h�(�X�r��"��L�z뭞���ݻ���DE��u]d2��'E������ߨ��b�������/
��y�y�$	��ͬ�N�S�\sM��l���/���n�r]o����}A >uK��~����*-p���Z�-���_Opr�l�P(��+Wb���_{,͜9���+y[�Q�i�&��W֬Y�/�FD�a�N����\.��KQ8Q���\�-��rf͚�ɓ'�<����سgO U��x뭷p�� g���o��֫�SB��҂��\���|/I���[����PU
�B��G>R�V�u�u��Z����mx:B!I��D�]�~�� B#�s��DQe���?������S��s
�(��V+]׭�V�w�M���7�_rn�.�|�����㻛
�,`��1��g�ȲȘ'� ��	�����|��Ѳ,���k�4m�c	�eY�j5�Pw��:H��t:�i�m�R�X|yӦMl%C &�D�b�詏P2�d�s
LKK���pgΜ�\��7���E��k���N/�xy����A�/i�G|iu�.�����<hIE�W�S�>w��0���ku�f���?���3�T="��碳�e����f#"��1A'
HGG�3c����h���)P^���S[���l۶m������č�Q.��x�u��0��w�&��%��Ʊhfi}̃֜���qD�Ac˖-��?�B%��F�u�'�*/�{^�u�����o����( 6l��0���26
!�L��(I�<��5gΜ	 ����:^���s�s����㱪J\��:x�������Kf����	|i����[hr�x��G]�����;�S��s~۾Rp�;�����1:�0�h�ƍw��	:��}��&۶�q��[}A�N�!�{�e����O��z��<��|� WsRį�RPˍ����|Q�7���^7-����%����o}̃�pF�V�����;�\�򮖝>}�S׃���פ@555y�<�m[�u�駞z�~�:U	V�"�Y8~M�uO����4��Q�no�R��ٳgt'@H��Uʘ���[��y}d�Z����=mc���gзlق;��q8����>L�6��q�p�T
�l6�Ȩ�I��T*�����ǚ��������GFԸ�LG�����u}���,
Gc!
y����d�8\&���(���E�6�6V�G�.�{�·{����y����mQ��瓸�h�&���wk>����ۓb�xA��Z�u���q�|���B���4mAWW�w|���1A'�Iww�ݪ�~���H$¢p4&���=mg���Ǝ�`˖-p �xV7-�+Օi���9|wSf�JBT����G?y�$>\�ʗ�fQ(J���@4D����b��j�������9$�����===i]ן�r�<{�IJT����Ǹ�[	��ﾋ|>�l{�5�v3:���*-��UZ�O�p�u�=<ٵk��b#򇗟#Y�=�n�"�Jy:f�8�`�S�>�(ϣ���]�|P,�ݲ����G�±�A<Uo�d25��r9�ݻw���|4�D���r��Wwxy�����U2f�6�G��E����6��"�~�m�X���a����Ә={v��ZZZF.)�N{jh�f,�np��A5�������ot]_�el*��T˥���$�IO�#}}}D3�v��1��}�����pD�v�Vi4�*�1�s �D��0�A��ѣ5��/��y������^� ���˺����琈t�2<���k��'^��b1D�Q�C"�$/7��뢿�?�h���ӧG�rX���W���ci��g�Ka�]1L��Vi~k�$����ܹsg�񇗟�x<�p�z*Q}�F��G�Ӟ�����BTaLЉ<ڲeKXU���;�BH&�A�EtI^Ο�r�����.z{{G���2M����;x��w7�����x爉;���k_H���bH'�{�X�č﵍#G*QyN�>]�A�J������rG�u��͛77�v"��ȣ�{�n2��g�0ϝ�X
�B�:�����Ǐ����Eܾ�:Z�.������q䔍q)��-������p�XD�]�G��/4 ��ݻ1m�4O��A6�E�X�,��A���`"/F�U�nIc��bs__ߓ >LtD��6?݈*�����B�੥ϝS%�R)O�j9Aw]�w����룈E*����U�e�m����Z�19��[��w�7��i5���.2�L��x�ƚ$I�w��������a�C"jLЉJ���Ӣ������F�<wN�M�i� ��q�СѾ�M	�,�\��Vi��[��_k�U��D�s�{����3Z��yY	�F��D�c5�X,��<��0�{/��BK a�5nq'*�i�?�,��$I�x��*��kopp�䭍��u]�߿��{n� T��+ê��v���"��{�U�u��*�O+���Y����ѣ�1cF���dpp�Ӹd2	�0|�����$LӄeY%��,+200�o �&2���t�lܸ�5M������f�;��E��6E/�p�ř3gF�F�"V,�
�g�l<�����Vi3��*�O�(����@:�L��4�S��x<@4D�'�鴧{M�Vtuu�q a�-&�DW���c�����2��Ω�����l6@4c������i��m!i���y�������b~I�����pM�H���T)�P��Q) �u��;::f�Q��c|�+�8�Om�.�;�x�'J�/�n�e!��M�TUE__��g�W.�����6~��@�!���;���#�"/JWoB���x�ͳۼ��ߏ���W8*o��,�M�VҘ��m�z�j��((�%��m[r�g j�L
��
:�����{�0J�`񺵘�O^�����M:4�����W��.�{��ߘ�w��Ԡ�O��׾��=7T�b|��e�{;"N�:U�g��`E�S�D"���iO-Ø����_���0A'�O?��"M�~��Xnm�j�%A��������ã_�r��U�GZ�}󱳭�l����R*.��g�W���c�*�7�B�m�<��6c"?��୪�����}��!�nq'��|�Ƕm��0+��%U� �V�ju{������	s����L/�x}w?�b ���59�O���!���غa��݇�V�>r��̙S�J�.������\�8��J9��iZI��M�|��NtYLЉ.����[����:.
qk;U�X,�@�H�Zs�����/���G��Z��u}�'qwL�,����.��,
�BMV8�f�%'���N��k�5�0�wvv�����PhD5�[܉.���g��i�e��v$D~�r3o�f�+#�b�8 ,�S^k���J��'��
��
�$`�����8q���x��AWЩ���]��?}�'X՝���Nt	�b�%/U��B!�hQu�r3_���#+� Д1u��$�X��_l+b�"䰀�������	>Ӯ&Kg���;&��;'�͛W�J��g-�@�$O�׉���H$J~;�#��<���DFTۘE]�ƍ���z�OwC�PMn����FKS�����޾xV���k�U���83d"�:�,@<W��q]�u��hJ��,C��/~?̟�P4]d2���p��]cMUU��[�h4:�0���E�a0M��q��]����g���PhD5�	:�����LUU�/J'������3/�
UU �����}��+K�\�}���*�    IDAT��q��Ƹ��O��M�媫�nZ.�4�W�T*�	��cV2v.9���e\��BUu����Ɣ�2&4�~,�CfM����뢿�S�L�tX%�m�����EQ&�TA@:����@ɭ9��7~��<����x@��$&�D�cY֏�lm���l�FU���Z<nY�h_i9̝z��7�v�m���0p&�`�x��a�U�����q\�?f��d̝�M)��J9l�q���(1J�SZ�������a̚Es�~����x���"U���gۭ��s�!TM$IB</y��m�R(z��`"#�MLЉ�������.)u\8fe]�:�(z��[�+��l�s6Q�:A�x���#��~���aթ�ViC9N�X�p	��Ӏk��UQ1c�8̘҄=���D��!V�_�D�w300P�H����&���ꃢ(�u�KU�������nݺ�Q�a�Nt��øm��.u�H%SVm�j������u=�h�5444���I�h�x����~�T���M�\N��G�O\5k<�s��:�%W%����%Zǉ���ٞ�e�\�N�0J�t�6�ou/U�X��͛7o����k�Ç( ��)F I��(�%�����!���e�M��ѕ�Z��dF~�}f�ƿ�]�k;M�p�|��;��`bsuWd?t�D(6�,�����r��\�h2�����	Ģ����0m����Ϯ�a�����4^�q���H��R�#������p0�Ֆ�C!#]]]7�~w��X�������z\���M�p��F���!�7v��iI��$�������iR�W-X�5dY��ŭص/Ӫ�2�6��l6[�H�a�N��뢅������)���j��� X������d2�h����&��V9��4��s������T<i#����(nZ"#*���Ἅ��ĵW/)��y��a��O��=g�|Q:�ki��v �b�@/[���0DQ���.T߼nuw]�b�G �Q��e�1����-�0&�:NQ�bPU�����,TZ.�=�m�.�����/$�k#5��;����m\��1�f,B��8����#Z[/A��!T���.�u}�ƍ�2���j
tjh�<��$]����q�$!�H�o�lq����`/��?����2BRm$�#�4q���c�xM�����	�����pޑ�ZL��)��5�����ֳ������??!���jtjh�B�i˲J�a�v�^�b�@$�:� ���RU�K�0��"�G0�urE�?wF+��S������t�4a����c,NJ�l��M�L�=@HD5�	:5����5M���q�h�[۩&��j~����i�����v씉��W���x�f�)��[���g��]��?��{x�y/��}���@	�`c��'���[����69��wڤ�i�&=mOJ��Mz���yzڜ��\��� L쐘�Nm'����K ik�ٳgf����X3ڳמ�����S;�5�I[��z׻.�~�7+�LЩ؅�aW�}���[6o�|�!��?�d�� ������pB6�#�p���q�q��ḋ�� ΍h�={��f���7�

 ����u��ILЩT%�IW��L�{�C�LЩ,=����fg:�L&]%=D*�K�>�,�"�ݴ$"�J jc��C߀��@"z��ΏU ܃N��m��0f>���_� $���L���Ν;�����:�ż��n����ON����Z8�C�������<�l���"�N�����e1�E<wU��f?�u��jB"*j�t��s���-�e9�\***��|����U��܄|X�;��1�qA�'���6t�'�N�[�C���큦i�2����CTԘ�SYټy�M�L�V�������%?��O.���-��Hɱ��h i�y��j�����K&7��$��B�f�w>��c�=��h1A����fr��g�S�����,���j�hʕ�A͗�k�rU?~���	:���>>�e	]׹�Ne�8��
`˖-��f���~�***،��F�$�NLNT�xLXQE,�,�)�&e�LЉ���i�<t]_�y��{QQ�ߓ��6m�2���v���p�g������BJKZlY����L��ߟ߿��JY,C(r4FJ�L&��>ꂨ@��SY��k�&��V:WY�xQ�(�}r�������@&�Q @�-D���������\:���Q��#���5*LЩ䵷�'���g��s󖗨����׍���d���Q��!�a  r�}I�5��M�k���M����M�'
!�:�����?��	�<&�T�,���i��2m!��W!-?�A��"-��_�RS������R��9��'}�ݜ�����;?��@4.�L:��2M3��QHDE�ObD<��c2���N�%	_��M6�����c���,��=b�\��0p~�@u���[ I_,��㑘n~߰ĝ�, �;��d�iooo� $����JZ6��l۶�W������ATl�<��q�qr����t ��sM���p�'��z6�L���nJgU�t*G�D����m��4��{QQ`�N%���)�ɬr:���������
���'-����4�k8��^e󛦄e����X0����G"����r�%��wBWǮe2��nݺƃ����?M�m��vs���.�����s)��ǣA�s�u]���Nc�VY��3~�wS���Q���b��H)�N���QHD�1A���e˖꺾��87MK��U��A��б��W����_(�����Ce�_�]��c���2~ܞ�i��c�\΃h�
�ͱk��/ݼy��C����J��@��s�z�F}��B�N�$�~l�5�D��?K� 	 ����<o^A津ěG�|��dU��<i�'/gq��D<r�O�p�RLJ�t*�p�H�lv�c��0�_��.2"5��N%����׳��\����`Gt%nV���`+�N�@��0r�,s�yt�~�2���`n�`�?H	8a��S���Q�l�{k�,��R���G$�-o�9�TJ\���lٲ�W=�H����L�P6���.�xܗ{o���0�c���!&3)����]E��#ؿ��t�7�`F����⮚0-���4�����:Fa��=�/|"�����gR�DUU��H�qS���s*5�@���)%t]�'�B"R�	:������d��:'c�v%*vnt�n󨩩���S=�݇ �X�(�}��������nK��7{��4��ݐ��kY|�;#xhWq�nK��?Z�떄��J�O�^�z�1A���p����J��g1]��l���x�2\2����f���x<��pT����
�|� ̘1G� ��6���	�]�����3K�^�||J���8ԍ�s��.ҕ�ᴍ����k�����B�cmͳo�v(ecpxl=��I��]U�"/�b1d2G����_�o�"*<&�T2}��?�f��N�!|�@G4�\RJ�/��Ѩ/�qGϚ���{7M,����A<�󟣥eM0G�����X\�`���r��[x�u���ABbUk�.���w.�;�}q�|�̙�|���wt*U�u�Q��0�7o����|�#��ahD��JF6��_N�$	hwzP��f����%�I���x�7b���$R�R����o_q����ą����'��f��mlD<q���Җ�L�lW?`[�?7�d��������2		�xm�[AU��?����"i�̙^��7+�n�c��`|�dtt�ѸL&�% LЩ$0A����#�|�0G�{�zN� ��8N��z�A]]R� ��i�dt  �Ί`�,`85�cG�gh!D" �e"����LacfUWϏ"(����]~�'�'rH��X�{VD�L-V)�7N\\A����*T�!X�N��D�L�=����aT?��#���G?�C#*&�T����1�dҗ�DNd2�K�M����Ǐ ��0��U�lx�n*�AT&/��6-����mK¡0�(���Ro�4�ԋ:��Y�Y���[��qi!�e��z,�����/�X��b��Hb�N�l|e���T��	 t�=&��{�7o��a�Z�j��jՂ�o�6�������#��,�4��H$c��.�H�
�0��g�W���X��c�ǰzq��/���.��766�)��rӵڲ,��� r*�#�N;]E�����[7n����y�	:�ޅ}G�p��ʅ�=�C�4GF� �����ݰ%����믹�>m�֨.���,��k �K�o�C�ᚖ�?~8q�,�ٳgO�~*TTT8�N�=����!�H$�C1�+ �����;�ږ-[��a�:q��ʉ��y!��ġL^I�s��9��Fll}6�/{?�e-�����$>��D^���6z���G"�K������3�ͳ��*�9n��z�c�=��DDT\A'_�d2_v:Ư���i"��!r��\UU���!���Ncc#����4q��������|](]v�l��������¨��o	�/\|�2{�l�VDq�蝹]E�d2_�mO�"* >��o����o������!)��QD��͊�nce� ����&����.��H��Na��n^Ɵ<P����{rnZ�������޿P��� 8n�E�g.W�6o޼ѣ��<�t�-�0�^J�h��S9Auu��1N�/&MMM8}�4���d�����{���xG�����x�����Qi�]E��&��aT�쯪�����NOW  )���D~�v=��~@�7Qy�	:���͛o�u���M�\�V����X,�P(��n�uuuH&�H�R�x�h��b��|�m��C�y9��A{ZG����׳�>�|��󊛗`��ò�w�����b1���:j\�����{�}�Ї��04"O0A'_2��8�ǹzNe�mIluu5�������X�p!^{�5 ���e����[�J�S��QiN��p�g,A�Bhjj*��p���t���==���#���DE��A'�y��ǯ�u}��1Bvn�������q~-������p��.#蝌�O�B�_~{O<��:���m	��G��nI�s xn������f|�w!�:}xx؃h��_,s�Ȓ�f�m۶m�G!y�+��;�L�N�����LT�FFFo����U�X������СC ����u�󄨜����W�xq���\=/�;�F�4KMR�{��+�.n�X�`��8򡦦�UEWЩ\i��x<�驔�t��|��Ȉ��ʶm�f�q��1\='r�`�H$|ݷ������{裝���*�Tt�x�G|�{#x~_���G��ħ��ʒs ����»ٹs�"�H(�e�jkk���rlGe-�H8~����m=���8"���N���d�ɲ,G���xܷe�D�r��yW�jjj��Օ�h
#c���8|�0 `��Y|��A�����=Y�q2�HH��ea�u�	���,�rh�h5!�,Y�8��q��s�����^t'��ei���=����(����%��ݻw���Nƌ��;]ב�f��·p�H�ɫ�'�M�z�x��EJ��	��%�olI�t��;�F�g�Q��n�Er O<�O��755�ڿ],�񸫪.�?'r��7��~t���\�$��7+�F���r9G��F�Q�='�`hh��������A�4G���H$�ŋc��� �Vѯ]*�q`��mG�U��vӵ�����	�/4�����G4=n_z�;w.ϑ�����N�{�r�p���w��3�l6�Y�c�zNt��А�1�@����`�+��Fl��S���	��,���<�+�@@�c����OT�=+�/97r[v�A�����=E�����u��ω.p�l��f���y�	:���͛��u�QK�p8<Q�JD���;]u/6��a�ҋ'3�d���V�ULG�9��u�}���8Z[[G4=�p����nv�JQ0D8쨠���>���yQ^1{!_�f�_s:��~�����J��߭���N�7,&hhh@WWlx�'i|��	�53͓����3%���k#hV؍}�N�Xxn��cՖ/_���������Wc�Nt�x<�pV����
�Vo""�������޾8��.v2&8~�JT'�P555�(��X�b������p��_���u�=F�J�l<�r��A`ek�������sFN�?ve`]�7g�̞=[qT�7k�,�cl�v�=���E"�A��ԏ��f�K:::������ahD�����i��p�r��s����y��kll�}��F�t�R��� ���^2/���z�Qi7-�QiN<��s���+V(�h�ܖ���,""�x<��t)%R���X�]TD����Tv���oG��������IDo��:���q�����ȶ����� `��*�����}�?G�Mի�sxa����U�V�DE��ٳ]��x���9��0�;������B%�_����D��?�,�QV��\=�7��@�Uyn1Z�r%"� ``���(?n��m�7��C)|�c#i�{o��O?Y���"��GОA���b�����Di;0V��m۾�\!����\.(��#�B"�&�T�L������|X���n�b�D�v�ډ��7N���/�����lN�g�e�����>*m�2Y�o�L#�{[R]]�e˖)�*?���PQQ�x�����%*7ne����!�&�T�6o�|�a�N�D�ђ(�%���訫2�����yV[[�k��f����_�Q�磧2cG�}�;#x�Y5�8*m*l����=7v�Z(��%��͙3��8��]Y ����*�0f?���xѴ�I-�4��9\�$D^���EKK��qMMM8t�P�R���CCC8}�4�}&�꤆EM���qp���^��QiS!%о;�C��V��X�vm�4������,o'��X,]ק|�����{���Ƚ�x5M%���=���:'cB�B��W!����>W�ϙ3���TV�Z��ڱB����8�U��l<�����)<�/��B���+��x�$� ��y�8p�za��娯�WQ~566������g�v�)�Î�����������%*&�T���iY���O��M].�ùs���%�;�aݺu���V�(:�me1��4����;��M�B��OV�cw�|s��T��Eϼ|q���E�0�|��_SS��q===y���t9}�,K�4�yѴ��oz*�a����y��s�����577��I	�p7�t��^&+�/[S8�W�������汣���ZcG�}���CE�t����|1���br���rI_�RPWW�T_�uG�;��h4������
t*:�=���aT;�惙�ܝ?�\��x<>Q^*b�n�喉}������}��e]zTڨ�{k�Ɋ���"���&%���:v���Ѧ�&�\���>��͛�j�ۗgD�J�x�&���x�'n�($"ט�S��f���pD޳m�u"�6�(f�D��r��牞���)8��c�ƏJ���ƎJ^8*�O����wcY��?�৯\\9ojj��իF半�
���8'�dy;��x���RJ�����7��'�4	"��Ν;#�����iN��4
aƌ^�ET���0֬Y�j��^r����e2���?G*� h���(޿��Q>���H���,��k �K�o��k"����:�{a���#g.��hii�ʕ+F�+V�jv700��zQ�tT�u��ů���>g��
WЩ�����p�Ɣ�.2�����.\�0����r���* �-������L��K��a[���+���~�E�� >��I|�É�Hλm�c{������+F坊�
ם�;;;�Q�p�,.�o߾�y�+��T@�b�槜\�i"��j����N���9WSS�����\E�F����[��K/��� ��~gz-<xW3+��~�k����r8!���!ܱ.�ڪ�y?��X�8=;�rL�	    IDATC�4,[��亵O������FFF�Q��F�H�R��đ��~�׽�����S�زeˢ���CN�'�����HD�޲e�\�,bϞ=DTl�ƾ}�p�ر��-����/|�sw�wY�ɞ,�8�C$$���>�&Z���߉aO<���/V���a\w�u%u��[UTT��np5�����sDD�%�Jattt��k��������w�	�"�:��S�0M�+lG�FWW��}ƌ%���=�-_�555x��WaYҺ�wv����0�5�hx,�x㤉]/�8�m�2�Ꮅ�wE�$��_��?�Q}�/�bUWW���/��m��纮cpp0����h4�(A�m�l�/ <�]TDS����a�\
��[�(��d\%O�/Ƌ/��R��jjjBUU^z饉����C�s���2Y�ݯ�=ga�� >v{��
A+�Jv c��������/|;!��҂e˖A+񿐚�W�E���d��3DT(�`�`�9�8����S�`�;���mppp��1���%�CTHuuuX�h������/��V�ea���8~��ے��uܹ.�kZB(�㼧��c9<�s#W�#�V�^�Y�f)��0�����]U��r9�ٳ�ѾY"zg�t�Q?!fΜ�+��{�S�E4%��*�|C��/8�^��pDy��ߏL&�jlkk+�=�{�@ ��˗��o|�	݃Nv[�������>��X
�~2}Ir>w�\|�(�� ]�D9}�4�s�<�F����R"����G�9�tR���=��d�\.7�z�h4:q��tVя;��G��9��e�&<��G�^�\%c�������KxN���]/x���ɏ�X+W�,��{qs��7�zq��s"o�?�lv���A3�G7n�hyѻ*�G�`0�)'�9���(MM?���\��͛7����W��&b�ҥhjj¾}���� He$:�S��W��uy�/��T���}�y9�W��.I�� -Z�E��E5�d,p]�u��&�D�F��t�4��m�7�����1A'�t]�]'׳���;RJ�>}��*z ��%K��+�xY񪬬�M7݄��^�߿CCC ���/f��KY�X���"hi�g�j����xn���g/m��i���p��W����d2���fWc��,zzz�c=0���/���0A'�X�NJutt����Fl۞r?�X,���J/�"*{˗/G2�t5���_Gwww�#�)%�����oNt{�lN] 7]��!ģſ��=h�ox�`��KWy��;w.�,Y�D"�(B�����P]]�j��Ç��ח稈h��𰣪.M��%K�$o����(���tR*�J}�Ir�����?�e˖��x�b ���9��'�@cc#��ۋcǎ]��l���g2x�:�7�t~K�1��xz�vX�{4��Gs�x{�u0DSSZ[[�617w�\��y*�B�#"�ɢѨ�ݶm��ٳ��u�"�2&褔m�8�> {]022���A̘1���p8�E����D����������(N�8��'O�0 c%�GΘ8r���3X:?���4nu}(%q��ġ�&��a(u�ʺd2���̛7�P�`��h4���V��O�8�sω<�ݜ��)0A'�X�N��ر����o���)?�&	�e�D�L4�ʕ+�i�Vw_y��Nb�6Μ9��gϢ����i�5#�9ug�P��*�I���>q7-�％�s6z-��p�����;?��a466�����˚R�j�*��ֺ;00���9""����Q�R�)_�Y���뮷�S"* ���2������`y;Q!麎��n466��5���^�X5.w��������0M������BOO�%G�+3�� �&�j�*���dL �A�`��@��I������1����X,�ٳg�������_Д���f�ɹm�8y�d�#"�w�F%�e�t:�Y _�.*�w���1�ל\�[���N�>���ZW[K"����j���kD�o�`pb��m�D__p���˖c�600lc` �wLo,CMMjkkQ__�*�w�L&]�r0������1""��@ �P(�/�a�	:)�wR�駟Ntvv�8YA���D,�2,"��3f`ɒ%���߿���y���ٶ�T*���!add�t����:/;#����������@uu5?W�4�֭CEE����W^��s�sS����Ry�m�M}Q�p9��8���9-ogs8"5]7��%K�����H��y��4i����JTVV�����_6�E6��a�f�0MRʉ����m�+F�P�H�h�Hy����:9�#G�09'R �8.s���� _�.*���okR²,G��C���W�ѻ8v����\��\�/��",+���(� ���,���a޼y�����`x�=��T�&餛{.��$�����B�s�ΈaW9�R"����S�\�O$��k�Q���q\{���r�i����9m4���<����D��
.�N��i����������=��ٳg��d��؍W�Lg���c�5�"��s�,iY�8{���(�w��
.������ٽ��8H)q�ȑi��_u�U����cTD�Z�t)���񽽽�cDD䆛��e�D��
���=���չr���x躎cǎ��iV�X����.ĬY�\��uǏ�cDD4.�ܯݴi�%*(~�Q�}�4MG]��~����������z|8ƪU�&:��ٳgc����K)q��Q6F$*"N}r�\pٲem�CtYLЩ�L������ �ۉ�бcǐ�f]�O$X�b4��������`�ҥӺ�ٳg144����(ܔ�g�Y�C����i��\��s��d�&><�3�kjj�ٝ�N<��ˣ��a�>}:�QQ���aG�[�u�G�]t*����kr�\���?'*^����>:����/�SDD��F�z��im���r8t�д^^�w�.�d���-[�,�(��a�N#����MӸG��ȝ={v������p��<ED�N8ƚ5k���PJ�C��0�<FFD�
� �p4�4��z��0A��1M�W�\��s"8r�2�̴�`�̟??O93�����i���ɓ�wN�.�D��Q(Do��
�駟N�1���{��H˲p��Aض=��������)OQMM(��ի�L:ځ�6����STD�%�	�a�O?�t£p�.��
"�J}ʲ,G�DLЉ�#�N�e��%K��ܜ����l|弢�bZ���Ç�y�E�81<<�)��!�t*�0~����P��/���� N�<9��,^����y����+97o��ƴ+H��p��9��r��e��bDa�J'�s�9�?uvv���{���?>-Z�����.�bݺu�.k�,o�������gM�4Wx
�%����x�kL�t�y���D�u��q�;wn��iii��%Kw�%��D"��k�N�[;p�c���h�"#�Br��iFb۶m,�"�1A'����FT>��T*5�{555aŊy���݌3�n�:�� _N�^D��P���t:��<
�ht�i�w8����D�7^��N��}���:�]�6/I����F�Z�
�`p��:u�T^�r�ZNWѥ�wy
�&��M�6i�i::ܘ	:Qi��r8p� t]���***�nݺi7���p�B,]�4/�GϜ9�3g��!*"R�i�����}W�)&��U�V}�4�)�	!�������䥉V$�ڵkQ__��Ȩ�A�X�,������p�ԩ�܋��s��=�y��[<
� t�����`0ȆPD%F�u�۷�\n��
X�b-Z��
��D"�u����NOO�?��{Qq���X��_<
� t�i���2����4麎����%I�:��Y��7tY�f����_�D"�������رcy���GL�|�G�`�Nڽ{w�0�9N��y�t:��_�l6/�����7܀����܏�O�4,^�˗/�[����N=zNN#!"�p������G��g���g���n�,k��c�NT�t]�޽{��������x��4 #�J&�X�n����vϳg��ĉy����-��4M��G�1A'�ض����C�����\.����ctt4o�lnn���_�.�eʋ���ӧq��ɼݏ����in��}£p����wr�����N?�ȿƓ�����s�
*_���X,�5k�䵂BJ��G�����y�?�=�LӼɣP����g�eY��������������/o�߃����&�@ss3n��F̘1#o��,o��&zzz�vO"*~.���硓G���'6o�|�������#۶q��ἯVVTT�����ŋ��,��CEE֭[����aؿ?Ν;��{�?8}5M3��c�q�<����	˲>���p8̒T�2v��i躎��Ty|����D^�Kj�A,X���-���x�7`F^�KD�0ި��g�a� �sr��<aY����,o'���>d�Y,^�8�5�x�V���� :�T*��{����;w.,X�����~9r�m���D�Nt۶��a8TƘ��'L�tt��ۉ �����k�᪫�Beee^�=s�L�p����ơC��Z�3f���ŋ�L&�~o)%N�:��g����D�?.��x
�9!�T��;v,���>:�����c�;MB`����={�'�7M�N��ɓ'a��'s�{UUUX�p!fΜ���s�<��S��ߤ������B̜9���{���W\A���5'��A&�Dt	)%�;������K7�����	�N�©S������*,X� �����1<<��"��y6���`pʿ��0�� ����Q�a�NygY��N���s"z'}}}H�R�ꪫ�H$�~�P(�����'O�ę3g��)P]]�x�b�=L�9sgΜ���rB������e}L�)Ϙ�S�Y�u���y]I&��޽{1w�\̝;ד��P(���V,X� ===8~�8FGG�>]$�@mm-����z���躎#G������(
!��L�z�4�y�)�A��joo����,˚�tmm-�t"����J���"�z:�����8u�=��܄B���-^���'N��eY��ED�fY��#9��L$��7���+�W�`��N�s!�s"���.����G}}�g�7����C&��ٳg��ىl6�ٜ����s����Y���S�r��ѣGq��9��"���iڔ�]�,Kh�v;������	t�+�0>��z�?'"�,�#G���[���X,���V,\����8{�,xn��b1444����X� sJ)��Ӄ�'Or՜��B�^��r�����	:�eY78����[���x�W��Ԅ9s�x~��Uu�4��ׇ��&�o�FQ__���zTWW���t:��G�bdd�`sQi	�Ît۶�y�!&�W�e-pr=t"�)%N�:���~,X� ����7����z?ʲ|"�@]]f͚U���d�m�̙3�����"��`�Yzd��B�B�2�&q�7;w�tuu�N�����y:��xW�B4�)%���'�����<�+cƌ��|�r���p��)� ���R���w�������ۦ~>�p��fdd�N'��`��9��xb<g�̙3��M(����BUU.\˲0<<�s������rt�n�������jTTT�	���8q�R���P����70�j˲D�- v{�&�7R�;�\ﴄ��h*��8s�zzz��ԄY�f){PSS������2�FFF022�T*���躮$��
���H&�H&����@UUUQ}^뺎�'Ob``@u(DT�B���&��e��	:�I���%߳,�Q�vp'"/�r9;v����;w.���W�!����1k֬��ݶm��id2�����:Ø�'�� "�"���(��("�b����R�w��:Ξ=���ޒ�6@D�#
9zqj����Ce�	:�eY��dӊ�.]�q���9sMMM���U�����i���Ķmd�YX�)%Lӄ��t��]R�
�
�|����9��gT˲y
�!fH��6m�ZZZj��)��P"*o������8}�4�̙�&����
w�11'"U�>���9� �+�6vq��ضm۪�����z��i����2$"�+
�B���GCC�����atuuapp��9)��������������_�0$*\A���d2�\��ωH�\.��gϢ������={6���ʒm����CWW���p��
��hY� L�iژ�S^H)opr=��Q��R���===H&��5kjkk�� ��4������{�^z""ծ��!
�&�{�A�B!��!R�b�DyaY�'�s���Q*�B*�'P[[�Y�f]�q9g�&�������3̉�h�7��4�r��ۮB�*�Jt�˲�\ϕ)"*f�eM��G�Q̜9���,�wɶm�?�����r"*z�p�gϞr3Q)�R�C�2�&qy���K&�3-˚	�V��4G ���9!D����?���$�@}}��Q�_4Emm-fΜ�d�]X����A�ܹs��-�JY)僲<��4��m۶b �R���7fTV
��;�m۶VM�V
!�]xS�r៙JSH!Lӄi���r�,�\�i���`0��3�����JD8FMM���Q]]��  �LCCC8w��������i���8N˲<�����'�'�l��_�뮻���O����m۶5��m۾]�+ �U�Tl���\��r"Q�'r剈J����Fee%���;~.��\.����chhCCC�:�+=�^�m���sy= ~&��`׆����1A�����< ��KJ٢:�b�/"�K	!�H$PYY���J$	D"�aM�m�H��H�RA*�B&�jF"*]NWХ����� ��R~���~Au0ņ	�O<�DS0�u)� \�:?a�ND��ƫ������?ŸҞ�f��d�N���d0::�t:�O"*+N�q���rRJ�p0��,�S�	�رc�z)�x���"�	N�]r�E�P�X�H�h�h�p�`p��:Y�y7�[���,Àa���d��:?������$�� ����m��.Ke��oڴI[�f� `��x��	:������4�@ B��������mO< J)/�bY?����s�{�]&���ƍ��/���M�6i�]w�R�/X�:�R�.""""*E���Rʿz���/}�lJ�&A߶m�*M����c)%,�!"""�R��(��i�o�_��EՁB�'�[�n��� � R�glGDDDD��i��g]�� ~��������?�:/�t��}����^u,��	:�*V�� ����Ձx�$����d,� WK��[E""""*ULЋ���������7�Tǒo%��?����G,UK9`�NDDDD��ICd&�u�G���^SH>M�u�ttt<~	&���l^&�DDDDT��>Ӵ,�BGG��$�Jb���=p����������"�2)����d>S
��>A߹sgĲ�����X�t""""*e<j��O���mܸ1�:���u�{{{{Ҷ��`r�Kx�����.�gd5����b���v�R�t�v��'��m���PK�bWK""""*u<V�w^�4����w��_���ڵ��ɹzlGDDDDDEf�mۻ�z��q�w	z{{{L��09'""""�"����4��=���O'T┯��� �ձ�s\A'""""���0��w��T�~J�E,�&��UBDDDDD���"WЋJ���ȿ���7	��;���T�A�Ç���������:���E��۷� �����X�"��NDDDD�g���i��m��s��U�n�~�����!�xLΉ�����ȹ��iwttԪ��{�.r�ܿ��:��ۉ����.���Ei.�����u��}��? p��8���������o߾�s�����݃�����  ߝ]W�д��߱m�Ǭ{VCn    IDAT�/�ٷ��M�\z�}��P���
�7�䜈������'�Nu�(��۷��n�q�;s���o�����\pzqB|hǎT�q9EW����B�R���Ł. �8�M!�))��< ���4-�iZ��r��*)�J k ���� """�rQf%�&����ٶ}PӴC�m�ڶ=u �RV!k�DJ��� ����d2y�m�ݦ�d�bL��'���B����?jkk{������s��J�4ߣi�}Rʏ ���DDDDD4N�m!���! �B���e��{���g'�ǎ;��R��c n�w�y�0�J}��U2YQ���ڵ�J�� �U��R �UӴo�_��P>o����F��	!>`u>��@ ��z����9y��R¶m�ɛ=B��M$[󽒼m۶Ś��������hж�/$<WT	zGG����8.cT�w�`�?��z=م=�!�����b�NDDDD����_ڰa�S^O�����B��� �^�����ھ�:�qE��wtt�P�:����4�3�ׯ?Y�yEGG� �@m��~W܃NDDDD�D��ؔ�d��q�Ƃ���1�_x���NAO&���q�ƌ�@��J��?��c�!!�ݰaC�� �m�6KӴ��]eoUbo�������*H���r����*�رcǯI)�@��8&B���Iu@���{�� �ϫ�c������9 �s�=={��� �?�,�����H�bY�t��?��ٳ^ur 6lx�u ^U�8)�^�I�+���۷�	!����۶}15
���q�� DU��t""""*'NK܋�5CJ���w����@��駟Nd���B�_Q H)��}��;U�Q+蚦�>�G2���bL����m+�6 �*�p��DDDDDDJ���wcr w�y種��P^� B�U� �
���պ Ĕt$���o��6Sq�j����B<	 �b~!4m��v���!�k>{�i�v�����*��ڳgO���k+���C�M�l���ΫB�
���
������s ����S |��rŝ�����`��A?$� �f͚\8�U /*%
�>�8�	: ե��molkkK+�Ñ���� ����c*�zNDDDD~�E���Ј�7���QM��Э2)���J��;w��Ya6���N�1�����E�����|���L&�g��pc���ݚ��&Ԟ\�����Z��M�m۾��WQ���������e͚5����B�룷�DDDDD�B�m��7n4T�օ��o*AB�G��jt)��N�c��/�.M�~��C �FuDDDDD��_�s�=GT1]B��	@�y�R����P�]�^J�E���%��|�i�qјBV�
!N$�ɯlBmذ��?Q5�B�"������j �X���***��h�۸qc��U��N|�_�����ȗ��_���t�q�KCC�w�'T�-����'���bn@a����T���/G�MU&��
���	7��"~�J&��VD>�Y�&u�BJy�������V4��U4�g.����B��&qDDDDDE㛥�z>NJ� Ê�V��*M�W(����lɱm�� �����S����� 6��[J�Lż��}��I5M+���ou�k㋪� """""�	!���:�:)y� �(����=@������џ+��`��;U�@DDDDT�
�-��BL�J2�|j��w��U0��=��b#�O7n�h)��`�?QQ�+DS9)�3�O�Ѕ���*�Z�S0��=
5���O�[0/(�=�DDDDD~Q��ц�����D5)�n�j�V>	�m��*��OѼs�H�C�� """""O���_��+��NŤ���ժ�TӴ�*�-4!DY�9������U�<�+����*&P�`N㗿��i��m�GT�@DDDDDޑR�r��	�t�$ S��5
�T����7��/}�V0o�	!Ϋ��������y�$�\��/4�)��R���� \�	��BϩP����I!�W�4�+�g�Pq�ZD��jt!DH��is*!�Uø��HDDDDTT�^��m�lNnB<��4���ʀ�]JY�n�R�X��T(�:�q\A'""""�?M��&��R&
=�m�F��ԕ����V(�S	!D�����Z"""""�)eRu�"��*�SY��+��rӦM���%�����\'""""��,T�8��.�pO�5M+�]JyN���5k��U0o�I)[U�@DDDDT�
�����	���ի�(x3)�@���5�S�m{��y(�?'QQ*�
zY<�U��IХ�}*�B\�b�BڳgO�U�� """""O-ٽ{wPu^�R.U1��_ż��d�R1��=*�-����(�.�DDDDD� %�t:���IT�R�WѼ'U̫$A�D"'T��������BJ�~�1��B�fd�vI?�_��nU0���Ee%	��w�9
�[��ՑH���]� """"*w:��������Pӭ����-�`^e%� �OŤ��}Bż��u�� 7���x:�'nٱc��AxŶ�M���y�&�{��ѝ;wF��`0�I ̆�����ʃ �q�Axa���Q Q1���t!�+���1M��V�/|���8������p���U�����BMy;���rUu	�eY?Q5��K�H����OhT��h�Q9�kYփ��ȧ��������SU+K���N �M�pdd�c��λݻwG�T���p]Y����XJ��X�A ����������A���Us!��k׮*U��S*���y���M߈�����8}.�3��4?_�	��s��J _Q5�BY�7�8AW�����d�\��y�s�΅ ��:�+aBODDDD�-!ğl߾}��8�˲�� hP5��Ed@q������!�J!~wǎ����v���,�� ��c!"""""�bB�����֎;��+Aحp~�	�������!hR��?�䓳�����ȗ�R�y���
:�E}�n�sO׶m�fI)  �0������ί6A�໊�e����)�;vlB��l8el*GDDDDTR�?ޱcǇT��D{{{LӴ�PX�~��ϯ>AB< �8���R�G�R���q���(��MJ�жm��P�T���b�����2�-t�4�Ǡ>�۰a�9 �� pO*���bO�;::n�|��%�DDDD�w>{�k�־m۶�Ur%�w��b��aձ �~�}��W�������O�R�����c�������<�Re,Y'""""��"xf��4���Z����O�R[<�: �P��\Q$�L�I ]����X,�LGGG��@&�q E���J|��������TD���ttt�>��y(ߺuk��� 6������ƧT ���  �o��y!�ߨ�c�A!�onذa�� :::���<J���������gF��ۀ���B~��f`dF�Im�H�\���B!�/$Q��KNn�/�&��bd��l�%�vX�06���w�I���VU�����xF�����~���9�Q=��������Yֈ��%?_�""b���\Qk-a�X   ��(Ͽ""A�TIlWض��s�=w<�"���?""���,�Ok���6m�����I]D�u�O�H�[�/�Zk}���������O���W������Tr�   ,-/M��k4�8p���$�n�5�\s����/��H�¹��V��κ���t�ED���ʿPJ]�u��VJ��a�<444��v���7k��ZD�N�ϊ��A   ��˞�����M�6ݘ�t��ׯ�V��?�������Rݸq�ǲ��)W����Z��%�MЎaRD�YD>=<<�`�7�����6��J��y�a�֖��
   8�.]�����'�|`�ڵ�$o����T��ok�? "+��w�&��i�s�Tօ4�*���8p௵�ͺ��E�F������7o�?�M.��2��Ed����Ț�JLW���   ,I)%�����Лi����ת��M�R��&W^y��J�sDd���Ar��z	�e�E̗��~�������D$�u�q�RD�+"wi����R��a�h�ka��Z��y���%J�3�֯�׊��i�1E�a�׵8   �qui}1U��R�Ga��0��� 8���1cR)�a8��^��:U)uf�/SJ�NDNϺ��RJݯ�~����\ֵ̗��."r�WnUJ})�:�4:   zE�:Ͼ���:?����)�6m���Ⱥ,�   `qQYh?���y�"9�""�i~H��^    �fV�U���Y�������{E䯲�    � ���_nܸ�Y���t�[n��oE�ڬ���E}�a�   :U�gY�}s뛷�r��g]ı�r�����կ>׶����G록,  �ân��ù��a�ذa�cYr,�����<���!"|�    �
��;��E: ���lڴ�F�Yׁ���  �Nųlg�Z�ŦM���u��]Ddxx��D䢬��3�<   h7��sgﭷ��7Y�\�ED�|����Z_�u!    z����J���ݻww�fX��e�ڵ��V�)�Z/n    ���J���T*ճ.$��
�""���s"r���,�Zz�w    ��=�Fc�T*�f]HT�ED���A�^)ugֵ    �^Qg���ʖR�N�4�<22�Dֵ�ё]D����HD^���nֵ`y��  �NC��(?�Z�ihh����c���ƍ'���E�@ֵ�"^�   ���w��"�����CY�
�_@��r��裏~FDޙu-��4�H�A�R%   @�È�y��Ŀ����oݺu~օ��+zӁާ��'q���W��  �nFC*�j"������("]l�*���8p`���R9#�Zz/X   �VJ)1��
�ZKv̑۝����M���u!I��5�ٸq�-�i�RD.ͺ�^�6�   Т�)�^�m�\�;���߿��"�"�:�Z�U�)�a�q   :B�:Ϻ�;�����7~.�B��u�����?c���暤�:   ��i��i�/��p.�������W)�>��zUֵt�(��Y�  �N�l�\�M)���7~/�Bڡg���7�`����W�����Y��-�   �Fl���_��������O[��
�M^x��W�j���ByY��t:^�   Ѝx��ĽJ�������^
�M=Л��?��d]O�b�   �3E�����n��֯�޽�g�"{:�Ϸ����Ȩ��S��	   ݆������|nxx������^x���W�r�a��Z�]DNʺ����   ݆&Tj��D���r��r�|1��8p���D���9"�9!�r'j@g�   򎀞�9���^D�߸q��ԱiX=�/��x��_�r��oj���5yj:��"R̶�l�>   ݄�ٜ��'O�~���n��7�|�O�/=!�\s�� քax�R�Ok�JE���`�)�����	�   Ȼ�����K�H��Zk�Ԥֺl�a�4�{��Y���H�UW]u���r��s   �,�k�:+�Z�;��p8��O#^�V)   @Kb<�ޙF�=t$"û��   HY!�#�a�A  @�"�#V��;�ax�rBw����4)
m�   �����b��ض-�e��8�<Vز���X���!1W]u�aY��8�}_|ߗz�.�FC|�?r��5k�n�   �*9t�г>��۶�q�#�ݶmQJ=144tb���AGb*���Fcu�ѐF�qܣԂ  �   W�:mHk-�z]�����)���vՆ�G@Gb��j�R�,�z���q�+   �i4˾Vk-Z�S,=�M���MQ����   ���%��a�wS*=����X�uE��	�   ț�Sؗ�4�+S*=���$}�0�e�:�qש   ��a��S�4��w�y0Œ�c�HL�T
,˚�2&�"    -QgxZ�5�{�n:NH��,�(�3�   y�yd�f�g_�x�H�al  ��u�9�!it$ʶ�/E�>�    ��;�_�R)�Qt$j˖-�6Ms��p��A�%   ���~��R�ts�%�Б4m��Q0�   Y��=�,�1Y�	F�rБ8˲n�r=   Y�q���S*=�����qm��Y�  ���8b��JA#�#q�m�SJ-����}   �$�ay����AG@G�l��eY�(c��  ��D}�m{�T*=�R9�at�²�_F���  ��D]ri��=)��G@G*LӼ!���C  @V�>��q}J���Б
˲.�r����5�T   ���?w'ҳ.�\t�b�֭-�Z�+�֚i�   h���7FFF"+,��,��(��  �n16��7�R :�cƷ�\�:t   �[�gP˲nH�������}!���F���  �6q�Y������Ԝw�y7��,�z�u�:   ��bt��m۶ݔR9 �Ҏ�<e@�VK�   �(Q�=m۾OD8z�!�#U�e}+��l  �v����7R*:Rf����\�:t   �C��ϕR�I�@D�H����M�mGZ��n�   H[�gN۶k�R閔�D���60M��(��  �����-˺3�R�#�H�m��\�Fq   H��:�3�aW�Tp�SJ}R)����0d�8   ���}�z���+�dpp�_S,	:ڠT*=hY�L�1Ls  @Zb�?�<��sM��:�¶�F���  ��T��H�[�u0�R�������r}�^�5   $.��j��^�R9�Q�h�0���)q�   I��9�i�ᩧ�zYJ� G!��-J�R�q�����:�   8��K)ǹg�ڵt��t��Rj����z��5  �c�s��eY_K��Y�h���7ǭ   +�F#��j��bI�Q�h�͛7�o��d�1Q��   �u	�mۇ���N��Y�h+۶o�r=��  �����u��R)���h+˲"Mb�;   ��_�0�1�r�E��V۶m��mۑ޺d�;   Zc��ڶm۾�R9���h;�q~�z:   Zc��S*XmgY���r�����~Z�   ��5	� ��ԧR*Xm����4�H��t�  W�gI۶}�0.I�`It�]�T
\׽#ʘJ��V9   �r1���V*���܁Б	�0>�� ��  ���Lo7��)��x�_�/�iF:�3�  U���e'�xb�f�:2�v�چ�wE�:t   D���8��֭c�&2A@Gfl���(׳�;   ��3�ݲ�ϤTp\tdFk�I˲"Msg�8   ,W�gG�4���~֟#3td�T*Ulێ4ͽZ���:��   �%�֑�H��{����*�:2�8οF�>Ci4i�  �.Q��%#M��q�9�r�e!�#Sk֬��eY����;   �'���~��K�`Y��Ժu�|�qn�2�V�1�   K�ZGn긮{�T*E�QH�3��Q�Ð#�   ��8�ٶ��)�,�۾}��lێ����  ��D}V�m��u���S*X6:�@;�sc��Z-�   �~AH�^�4�u�o�k(�9:r�0�����4�i�   X(j�\)%�B��T	�p����8SQ�T*���  @�����8��������"!�#7l۾,����s&:   ���둗Aڶ}IJ� �Бn�f��?t�  �uz�i��0��)�DF@Gnlذ�1۶�2�R�H�i�  ���s۶V*��L�$ 2:rŶ��u��   �����R9@,t��]w��)˲"-,���K�   t��τ�m���ϦT��{���u����}_|�O�"   �]�^��<h����w�f�$r����q�Q�D��  л�l����JZB@G�lٲ�f�u�2�Z��Y  @
�0�D��>2::���Jb#�#�l��T�����	  ��gs8�q�)�r��БKg�q��,ˊ��hnn.�3   :[���g�q���R9@K�%��H    IDATȥ�k�6��V�1AH�^O�$   �L�Z� "�q]���k�F:5h:r�P(�>��  `)q6�+
�B)@"�ȭ���;\�}8ʘz�.�o�  t;��#Ϟ,
���?I�$�et�Z�P���c�  t�8�s˲>�B)@b�ȵ;��ǉ�={�V��	   �#��ݶ���~��O�T�:rm��ݡ�_�2�#�   �[���
�v���T�:r�X,~�4�H���  Н�֑�4������T�:roxx���y7E�!]t  �.T��#/gt��y��xJ%�!��#x��!�\  @�\�t�RJ��HJ� �"��#�w�y?�<�(c|���5  �.�h4"?߹���m۾�RI@����m_uL�wX  �_q����)��B��:�ڳg�T�V�2h͚5b�fZ5  �� �C�E���]�V���::�.
��:hvv6�Z   �F1���9:eŊ�8�eL�Zߏ4   9���T*�Hcl��O9唏�T�
::����ˮ��:��  :W�����:�h��g�ʕ�7#�T�j���L   d/C�V��Ƙ����H�$ 5tt�s�=��B�pS�1Zk��   (�~B��������)������T(ޫ��4�R��E  � AD^{���B��JRE@GG��P(�e]t  ���٭P(�222rw
� �#��c����/N=Ô*  @R�v�]����JRG@G�:���z���(c�  t���9�:���ݵu���T�:::�m���0�}����E  ȱ0�=�PJ%mA@GG۶m�7
���Q��E  ȷ8��B�p����u)���u��g\�E  ȧ�͔b���S(h+::ޖ-[x��P�1t�  �\.�Y{~��͛�M�$�m��
���n�1�r�s�  r$�XM�uY{��@@GWغu��
��#Q��E  ȏ�k�غu�)��]����CQ�E�����  �q��O���{)��]c���_v�Ѩ�fff�(   ����c\�}x�֭_K� tt�q>��^�դ�h�T   ����X瞳�݆���r�|9��""���)T  ���,�8ν۶m�J
� �!���8���]�z�.�Z-��   ��F��9����M�$ 3tt�m۶�P(~u���l�]C  К8�����m۶ݐ|5@���J}}}��iFJ۾��E  h�j�y/ ������;���L�ѕ�?��;]��n�q333t�  �@kk�y�P�i��ͷ�P�9:������i�a�1aF>   �U*	� ��4�i��H�$ stt����G<ϻ2�8gp  `��0��s��۷o�7���\ ����X�❖eEZ�w�   ��\.G^VhYV`����Jr����6444�y޿DW.�#oX  ��k4��
�-�J�)��]O)�a�q"����  �c�3SѶ�O<�C)��
]�T*��~4�F�!�j5��   zR�V�z�y��8�n�:?���\Q)�^�gϞGk��IQ��!k֬�TZe  �C�E޹�u�Gw�����Jr�:z�mۿ5h��a   G+�ˑùRJ\�}OJ%�C@G�ؾ}�~��n�:�R���3�
   � be�R��Jr����bYֈi�a�1Zk6�  h���l�c��=�+�T�Kt��R�t_�P�8�z�Άq   1�}�*
{�l���Jr����s�I'��u�XǮ��"  ��i�ezz:�8۶��<����P�kt��u�����}(Άqsss)U  �}���"o'"R(>�v��F
%��1k�Y{�R�����֬Y#�i�Q  @��}_>y\�P��Ν;�H�$ �蠣gy�w�i��ߡ�3M  ����d�4Mm���:=kdd�b������0  ��*�������<ϻ|tt�G)�t:z�)����q�J�q333��Nk  �	a��l��xŶ�j__��J:=�Ϊx���8�q6:  ���md
�?fG^�46�$��q����8N%  t�z�.��
���ܹ�)�t:耈��9l�  ���LMMEg�.��P�q耈l߾��B����� ���
  �����ƚ��yާGFF�N�$��Ё�Y��۶'��+�˱v)  ��FC*�����8�����BI@G"�O+�JA�X�g������  �EZ�XSەR�yި��<��̳m۶����Q�A �r9��   �mvvV� �<���m�vm
%��,P�Tγ,�uS� @����27�d4˲��emI�$��Ё���̸���8c9  �
�u�m�R�����R��N����,a�޽�V*�WDW,e`` ��   rcff&V��P(�`�Ν��BI@ǣ�,A)��4�F�qsssR�E�!  �1j�Zܩ�b��!����@@�066v�X,~8�����X�  �]���������ᑑ��	�t��Ǳw���*��oD�8��Q  @f����Z�FW(nݹs��J�t�8<�{�eY��g���)  @^U��X��4�F�XJ�$��Ё�9\(�(����Yi4"/c  ȝ bOm�<��GFF�H�$��0�X����۶-�����J�,  ����x�<��;v�&����CX&۶�lYV�9]�FCfg9�  t���-˪�ȹ�Wt':�L�Ri�X,�#�X�^  ��^�K�\�<N)%��{ǎ)�t%:A�T�R�X�z���  :M�255k��y_ۗpI@W#��y晛]׍�Np+g�  daff&V��q�陙��)�t5:�ڵk���4��;,�j5�^  ann.֑j�ah˲�{����Q6@Dt �R��b��Oq����J��Xu  ��ie�[��>366vc�%=�cր�ݻ��J�̨�Ð5k�p�  ȝ0e||\� �<�u�v��uZ�U��:���mێ��P&''�7�  @�����
�e5����S(	�t�ccc�۶��8c�Y  ����ΕRR(޿e˖�S(�t�Eccc������3�\.s>:  ȅF�!333��
��o߾�3	��:� �479�s8�����X��   �A���m�����H5 t �R)(
����P֣ �,i�ejj*V��0��uݷp��:��R��㾾�?��3���2==�BU   �6;;+�F�|],?�}���.	�Y�$l߾}ߜ��{s��+V���.	  `Q�ZM&''c��<�;v�xk�%=�:�0˲��8�q���̈��I�  �,����m�۶=�pI@�#�	{z=��,ˊ����299)ay);  ��5����4���K�R=ᲀ�G@RP*�����w����]TY~  ��ʦpJ)�<R��)��<:���[������gl�^�})  �����J����y�W�o����K�46�ҥ.���{����q�i  HR�R�}r���ڵ�ԄK0t ]�q�Wٶ=g���t�w�  �k4�g虦Y[�z�o%\��@�J�Ҹ�yÈ5]err��� @K� ����X{������6<�Bi �!�mP*�n,�gls#vv  q4wl�����GGG��pY �t��.������[�uGV�Z%qv�  �kbb"��9�u�۵k���K�:�@�ܹs��8�����   �V���m�W��%\�c ���\�r�eY�8�+�����k  ]�\.K�R�5ֲ�����+J�R����F@����{�X,��4�X��ggg�V�%]  �"�ZMfggc�5#,�C###O$\�� �(�J7:���'''��h$Y  ��z]&''c�UJI�P��R�tc�eX6�2t�%�|�\.��8c�R�z�j�,+�  @��}_���[ٱ�;v�xg�eX&:��={��R��^g�i��z�j1&�  ���0���q	�x��]�=�k׮�&\�x�2677�Z�q�36�t   �ùmۏ��ͽ!� DDȁ+���ĉ���|��⌷m[9# ���Y�i�����V*��L�, �Ar����6#��ލFC���b�7  �Ik-SSS�����7΁| �9Q*�~\(�aF����q*  �3���J�Z�5�0���?�}��[.@Lt G����y��q��������L�U �<���������]�ݽm۶�,	@�X��о}�>;77����������/ɒ  @����f������ t ����{C�RyS��R,�,	  �@�Z������=ϻ~ǎoK�$ 	!������sW�V{I��X�B</���   �j��LNN��v�zy�%HkЁ�����t���i��jI�  2�j8w��N8�	� atЁ�ۿ�������F��J)Y�r����ti  �M���LNN�>Rղ�Y�qN;�pi Dȹ���C}}}��,+V+\k-�����G  ٪�j211;���Y+
��p�� [�n���o2Ï{���Ii4I�  RV��[��0��7l߾����:�!FGGz��v�Tg��Z���� �!�FK�ڕR��C۷o�9�� ���t����o���a��<�N:  ��h4Z��n��<�;v\�pi RD@:���襮��vܐ�����	B:  9��pJ))
�r¥H�@;v��l__ߟ(�b�o�t�� �/��y�Z�&""�b�����>�`Y ڄcրv饗��r����|��8	V  �H�s^,�vtt�O.@�Ё�o߾�W*��'� йZ�""}}}��@�eh3��nll�#��4��s� �N�^oiC8����!���:�%�����J���V�r�J)
I�  ��Z����tK�X,����ػ��
@V�@ٷo������K+��b��TI  `	�jU���Z���y��رc,�� d��t�K.����ryK+� � ��r�,���-ݣX,~ill��PI r�5�@�����wY+����i��  ,�R���s��΁�C@������Ba_+�H�}  p���Y���n��b�;v�ؚPI r�)�@ۻw�W*�w�r�ue�ʕ��J�,  z����T*���Q,�����#�� �t���ر���ϵr�Z���  �2��LNN��=����ntЁp���c�V�`+��e����� �\a���4�����9��-�� �O�@عs��z��Z����211!a&U  ]-Co9��ŏ΁�@@z�����y��׭�%�}_&''Y� �q(��V�I-�g``�/���� �� �S܁��/~�wggg���:r�6C֬Y#�eI��K `J�#K¦���\.G��a�X,������.�� ��A�^z�;���>�a���f�q���Zk�� 0��p�4>>.�ju��0C
�w����{���7:У.����J�� ��\?88(��=��t� x�b��СCR�׏{�0B�uK;v��J���?:�������Z�v]���[�r�����^��� �S)�����0�СC�����������[*���F� ���K/��׫��|�v{\D���eŊ˺! Ћ�X��AȓO>���0˲*��vll��4j�� 䢋.z�R�'�z}p��=ϓ�����-�)� �^q�)�Ki4r�С�~Vڶ=����[�ly8�t: ����k���Z�T�ue��ձ�T#� �]�p�T�VebbB���8�#��y��ɄKЁ� �����F�q��h�}�s���y�t @�j%�7��e�V������R��1 "B@����a���>8� �m����8���6l���$j�=� u��W��Z_�D��_�4����  �dɄs��:ܵaÆ/&R����� ]��o�W���uY�1�KjNL��  @&�Rb�f�?˪ڔ[���p`)V� ȯk��y�B�f=(+U��{���t @�Ib���ȴv�:��2-�]	��K�ApL�ڑ���.�|/�0� :F��V��}rE�t��-��� ���M��q��"X��Rt @�%�<��p�\�*�.�� �%%��/��O��X�>It%  HRR�\�ȏ���w��I��. ��t ��� s�#o�K���|�i�M  kI�7�Ő����@U�%�� Dv8 �JY�-�+��!  Z��̮Ym���i�s ��T ��ړ���ca��q  +I�&"�hX�+�ɸ.$P�^D@[U,��?Unִ|/B: �ݒ����`P�	N��f38 �@KBQ���2�y������N8�a�֚u� ��$�Qr����J�~ z@"�WɌ��[̇�����՜n��h�ַ ��$��%��O�'���� �)� �D����{P�(6 @�����.���$�'_ ��[4N���Չ܏�� �V%��D��O��r��T��
 a�� H\(Jn�O�_}��qTk�ɕR��bm:  �$��7Đ��'�}��D� ���p@&���-��2��-߯����fm: �L3�է�+��_ ��M� �S��jJ;rE��v�e�; �x���&��p�\�8�p ut��.C��?O3��:�11��i�� XL�o���f��rgxB"���!�h�{�U2�(�:�aY��-ߏ��  MI�5yjJ����8]s m�w muH䫍�O�dvyy����@oJ�X��v�9�v����1�`p�<���z�Qq$h��͝��@�H�k�C��,�d�v !�����
9��d���<ר$r��A �W�M�$gN=�=����h'�{@TLq��Ym����� �x��� ȇ�O�Pr{�F4N#��O� 2��'�/�	b$�Iz�#  ;���$_���^=(?��+���	����
 7��+}�)v�_͝ޓ�
	 h���"�R�g�2+l ?� rE��gRVE�j3����; t�4��u1eF�h����@.�Œ�6ΐ�������3� �/�#4���+�IUXk ���@nUĒ��ʯ���*�	1%L�͠�N� �?i�x�Ő���g��� �� rM��O���`�/�7%'s���0�Z� ��4�NyB����d��t :��0���?M�4'�5��b���J)�ZK&sO ���}1����=8A��� :@��"��`P~����_��rb�f�; �_Z�a>�;��2�� :@ǙѶ\�*/1&����b'�6]�i� �iu������w��5Й� :������P�_^g�J^�p7�9흠 �J��ˇ�~�^p�������]� :ZYl��?U^h����cR�Fb�f}: $#����S'~��?W�	W%~o h7:���`8 �Ջ�
�Iy�9!������t�: D��:s-"�W���D�j3��@� �F]L9�$��+�l�1T�D��Fr �|iv�ǵ+��'Oh/�{@�� ���(�7N����|2�#ٚ�� �: <[��<CnN�ۂ5rt�.D@ЕBQrgx�<����r�1���AP�g��ED��}�$�e8 ]�����hG��O��ey����T����f�����ڑ��I�P؟�� O� z�#a�|-|���8,��:$V�g��p4�ޓv0ohCn���	Lg�3� zF Jn��=�U�j�	y�1��#A@/H�,��������� z@ϙӖ��?O�6V�k��w{!��Ni�á+Ó屰�ڟ yF@г����ty�1%g��%�ۻ��A�3�t���y]rsx����tv =�Ⱥ  Ȗ�{�Ur{�:� �<C���; �RJ��4S�a���j�y0H8�������.w�v��A��� �*��ߚ��,b8 x
 �0�T֨țvs^� `qt XD��]A]�7x`�nYt� �#��1��i�o޿� KX��v����1�(� ������45�y���vu˛� �� �vM}a�;��3���" �G@���iC�ƕ    IDAT��DW@��.�� $�� -h��."myf�w �Ѯ7E� �$: ���P��ܭ�A}����1����-!�@� ���Cjs3�v=(ϟ��F@oi���xc ���Ws ű������5w}og`VJ�i�m��
 �����0� ��w��?[`Qt K�3��i�+�M�ܘu-�j~Po��l�{OX�����v���M��x���Og]��"�8��֟X�
�����4���{
:a�|�.y�����[�D�,�qғ�EG�i~X'����^����E0��u�K�,��ғ�ugjaW��do~0�"�g�b#����`����rӥ���)�@{5Cx��P�w�9"q�s ��DBHO����,�W�;����<�7Ƙƞ*�9�X� "k�t%�?����a��bk`ē�Pޜ���o�#���� ��֟X.x�Bzz�?Hg��j�,6�:�³ʳ��Y8��`�*�9����FHo�<u��w�Y�<c�2�,�*_(�qz�@�� ZBHo��u֭�.y^ް�[��9�D������fP��x�g�[�CX���.y��ny֯=�p 1�����ҳ5��</v�	��47w��Oyڧ���$�� 1���i��<���}���t����N������� �H@���0�8�<>�/�����C>���!�H@������>O�����tIk~--���uF(�-�9�������O������>�/RySȗ��|�t���s�p Ut �!��['ǴX�3��[l���@�w��A8��������a~@���˱Ԕ兛��;����Ra����	��p�-� RGH�<�֛qC{���^3��h���bo�t��3V��p�m� ڂ�޹��N�C�������:�b�������Ŗ�t��O#�h+:��!�w�n� .��3}�؎��^lZz7�.�=�M�'=�p��� ڊ��=[CۍAd��Ŧ�/��.�n�=:ͱ����/�������b�7t��A"�Ȅ�u z�E�O,����7T+��k�o̺�na(��@v<�u֏������Q��?�p�r�b���R�r��k���F8�:� 2A'��-�*vs�=	�C�bk���|9�-6n��~��4�n����8
�@�� 2CH�7�"� ��#�k�g�d�� S�����Hr��`��!��{�@.�d��'����U��Yׂ����w��%A	I9�C|��.W�Km$��:�\�3�����'���p� E�±,�:��o8����/�Ⱥ aw 9�JXͺ��b�j�glt�{�|O�FTT�� �� ��5z�B�P�}�{� ݆� �J��/�<�5�����q  z �3��q_�׋}�x����� �^G@ @��5e��C�bgLE  :  �%p�_߼�X]��Y����?�n  �G@  ��ظ�6�0�j�&� �.:  9G0 �7Y      �     �    � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     ���.  ��W2 umf] ��CR̺ �: �ȸ.ȸ.d]   zS�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     �     �     � �    �t     r��    @�    �:     9@@     � rCk���:�B  ]2�� @�� rCi]m��R</ �a�g~m(5�]% p4:��0���/	�� ��	��Z��t�� �Q� �#��"� ��������W@{��y���~��Jt @hY��>�3, �B@�SA�����  H�
�7�uݶ�ɲ ��� 7���j"�@���Z��  ��U?�k-�Ⱥu�f3, �B@�+Z��_�bV�, ЅN1�ٴ]i}0�R �Y� �E�o5���o  �z�����Է�q) �@����V���6�Ǻ �e[��G-�҆A@�+t ��Ʒ�����͏_jr<-  /�fD=���ox�[�̮ x6:��1�/4�kִ� h�-/����֟Ϭ X@�Ap���"O��~�5�qE �Nw�9++�#�wbgY ,�� w�p*�}͏_c���� �I�ȫ��y�P_z�9�<�YA �:�\2��	EDVu�u��� �x~͜�5�l�C�>�e= �:�\z�9�ܥE����l��T�eI �TP���9��'������ۗ �!��-���PDfED<ț�'2� �i�d?)�3o��)��H�� �����o=,Z�U��X3�rk*˒  �%֌��:j���>�-oy �� ��� r��8� "�m~�f�	9ѨfX �<Ǩ�ۜ���`��>�z `9� rmݺu����"rHD�RZF�GdP�3� �W+TCF܇�zj�Q��@뱵k�6�5 �F@�{�54��6�w��g�T #�G�g ����0|�RxD�Ϭ;���x����eY ,@Gx�[�z�h�.��D_���}P��̱9 ��ڨ��YVZD~�����ϰ, X6��κ X��\w�G�ȑ5�5m�u��䞠?˲  ;Ü���c��Oj���[��o��
 �!��8߻����ZJD���~�X%��#�VV h7S���9$�iMȼ� �����_����U ��t�o_{�fC�/�ȑ��Th����}A_�� ��TsN��<1J��HYi���ׯ�RVu@\t �W_�1�/�R�1��E9�8A~zY� H��FU^c�����ߺ�T�מs�]Y� �"��h7�t���|L����X������+�ޠ_�	 �RZ�0g�׭)9Ř[�ہ��W���k����� �)� ��w���7�0>�D�^�{u1�>�O��PP�imgQ"  ��!��y�Q�ӭ�8.v�����9�����@�� ������o�a�QQꬥ.�jS&�-��#�{w�i]p���̮�e�nfVb�ه�EE���D�DHt$t�IJ�P�AD�lV��a��b��k�����<���;�����N�{��f������>:/�#ci�\�dZ��9�Ǯ���{<>v/���Y���m�<_���P�-pJ��)��7���y�����1�g��{ ��y�ʘ�Ͽ���o=�� l7���~��z��]��1���1ƛ��� ؔ�4�2������߷o���T!Ё��~�g����-O�E�<�p��g���4����p����;:�y"���Ӂ�<oi��C��GO�li��l�M�:��v�#���V�����//>w;nZ����{y��mu����5+�:o;nZ����}������=�o~�wz���ᤅͻv=8_rɷO�3��y>2��1��y����y��k���d�p�t ���7�c��O�C������ꚿ�x����|���������꒿�|��1�۶�����W����.9t��4��{��M�����ƭ.�}Ϟ�Mc|p�ٌ��=x���L �|�   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t  �Tv  IDAT �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �   +'�  z����e����c��s�����}s�}��~�ɛ�G7�Y>:�̍�rdZ{��ii�F3����W�i<m�}�<��{��,?���fn<�yi��8�v�F3��s���K�Yd����}�>��l8�c��M�x�g�G?�6�v�F3w������Z8�����޽�Ȏ���&N<��ȑ��KK��h��k���ع���y>�c{�F3k�ˏo�F �: Op�ַ�q�ׯ�暥���{���{���;~�ջ��+^��'�yt���O_p��g��E'���^����lf�O��c��Ⱦ����K��-��g\�}c��6����������<x�uw�����C��cܿ������c���W=��	��S�?q  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      VN� ���������_��/��q;�0M�c��������|�f}a��������}�&�4Mӹ�>r\/٤i��<Ƹc��y�׏�9 ���y�O�   ��O�   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �      :   t   �    �   @�  @�@  � �   �oO�=�     IEND�B`�PK
     �9s[�����  �  /   images/50196d33-890c-4789-8115-a73c306e50dc.png�PNG

   IHDR   d   �   1�S   	pHYs  H_  H_#�
{   tEXtSoftware www.inkscape.org��<  6IDATx��]	tTU��߫Je��!$�!�g��6=Ҩ(.���ʸ�8�L�����l=����Q���s��TPQ��i!�;�RI*��7�w��QVBR[.�snR�������/w{�Ig!V�X!���wEQ��ɓ'���	Y�|y���{G�_}��$+�#�#!2\��p��4�S?N�8p�6��sj�t�S�}��r:�)���#!�/���6��ʢ��zr�\TZZ
�3�����Fs�)�Lb�0]m�p���jNk�>;N�8A---���S0���|�6m�4z��7�|�|>y�^
�����!��n�t�r?炄��|�k$����B��_TU]��|����I������/Snn.�z��S�BV�^M���'��!�BX+.b!=�?���
5M�&H�i��Ʉ�p��Z1���_��]>�[.�_��ЪW^y�***zĜe�����Ӟ={Dś��A�(n����n���V�����aw�\$��M|�B&bV ��˰��o���-��Ç��W_�;３2�����R|��%����A���E��@xH �
� 9�����"���l�nf�y�_h��d����L!#����k�q��,�k����	5FK�u�h�~qq1���B `����yp�0�@GĘ�CC@^��\�����s=��L���//���8�;�t#��D�YC3X�N�l~ɇ�����yB���d���'O���ǉ(� �ȷ���(H9p� ������q=�%k� N��5Oq�ebC��2k�,J'�J*��@,�J�ϯs�����(�'�B��۷/4HwӦM��{=Fk.++�_p�"��������} h-�ǚ6��h.�L��H&HI!(8BZ�<BN5��-p�0��� ����Bv��I{��%�K��Q�����444M>|�gw����{�}!&�J��Ϲ�S�~[Q�t��B�X�Ͷ�H�誉`�����O�>�a���Ӊ�o�����I:":t:G�-|��ݻ;5_&p-�())!��al�V��k�N���������|�r�Õ��������Q[[+�8��BP��������9��t��$��ѣ�̍5
¥cǎu��({�����;N�0��k�}J	Aag!�p6ˬdt�`�]�0=<�����Dy�^�)n��ܐP�V���7�	���K��P�s�k:$L������[Lu�dR�q�.�su}뭷RڳO)!f%��y�%9$������oX����}t~�TS�Z�:ı s����c���Hێ���R�)��+D`�u� u�bs���v%׷av*�2B`S���t��g$�w���)����EQ�|�]�o��&��שūS����U�0?�*ˈ
rw��̢���bX�~ɑ#GD�мD�:�������a�宻�T %�`��O7���E��	�9QY�E�}~ꗿ��P	-�p�y܇p���$��O��6���^���u��' H4��j	ꄺqg6[�/�����7�x�n��6J)!�6�Qͅ{
�3��5Q8�S�W�@{#UV�Q}#n�n�\�+9��0\d�7�)T��Ow#��#B���@���Cc�Kʇ����}���|�sڇ@&H���p��>��{*��(-4y��- tA	���,��n�D�񚮑檢��

�7��{���z�����s�Q�)�#� y"��5���aʸ1>��݂����N� iB�a&�Ӡ��k���ؚF�s]!*+R�Y���ߙSN*GQP$��8�F������H>
E˅ԕ��3 /ԕM�t���l�>46�AR��E �*//W�I�;�~���
T�n��Ǡ������k�{���J�F�[uD��t򴅩͗ł�3;{�;Yᙦ������o%�'-Y-I�S;� 7rEǂ�TL(��'C�☪�TJ�d�~�(!Uk�l�@s3��9�Q�S��Dda*X'�X"R*l>�:s<�;�7����Z�H�L��Rk׮��c�>'ם1�� ��H�,�8�H���2�q��z����6K�"��;�ueq�J
T������ɕWN @�З0C��:�x@٠%,<��W_-7n-Z�(����	�v@�/�䒉�u
�
퀐�7 �g���.���m����)l�t��ag_����S�i_v�7�{�Y�LUUU"��X[*1�B&x��_<��Zs&$L̉1L2�abRA�|Ё1b��8�PG�O�Qaqmo�kj�n��bk������: L�uY��3��J+�d@���{��%F}�~I*��ct�-�,��+���w���mq	;���~C� �cr	-C��ׯ?%@v�E%���c�����
����{�]t�[ʡ� *.u�5�7�6l��̥$e�2`B��L��6%j�"�r�yMdZ��E	]���Fh�B۷o�0����D揠&��y��1�뢜�����:x�`��5��T��?�,8o��e��q%D����&#bId��L@��#0/h��\��x!r�0���-�9�p4�2�5���z���ư4p2�s�fA�����&e<ZF��J�?HA$MA��Sb�C� ��C�R���ŸFx�A�	Ȃ	�`>�<���{�uz�;���C̥;���)�~����ǋ��5W<Z��j.t i[�lI�߈�!�!�P��=�����k�s�4B�-[7����;����{�	����o�H-Z<�4���������B�t�`"���퉕��8���u�]=%��&�:�3��?����3�7�J������A�LU�x&�2��
!,BbhLʁ^=��.��ݘ��Hq/L;3�eA?J��4��Y���巔˥��~ʔ)�x&����l�;�9bo�h*Ժ
ӡ�h�y�jj&��-#c0�ep�L�t��C����돂�v 4���s�wqk�nS�:Z&�)mMVY��C�?��3�Db�ΡSd ���8ab�aN7[s�)BdF# �9=����N?�_YC�O�'
B��'�������ZN�8M1��	��B`~�]����rz��~;���n�d�>��"�ŀ��ގs�ߓA��.��q�A��I�my�Ld/V]X	�m3�)A��]��l͎#d��VB�Q�#�v���$NKc2J~YŹ�죘c�m���Ed/`u�`���o/prsZ�)��?p�����Gǈ��`a��sـ�������Y���ԁ�)Ia�$��p��(F�-� B��"۶���RD�QB0�`?�ɩ�re����C;��.:�����[N�)"s2��!�&M�vwP$>�M��D�Ctp����d�4��8<I��9i��E�&�����	Q��^����#��f<t�Pߖ-[n��oc��,�!g,;ǜѣG/޼ys��!����.� W̰�w2��*��UU�eee��2�s��x<~M�6�[�N+..�t��)o+�J2މVO<������B��Xw���d����ۇ��3�1j�0Smmm������T/r8[�imn�b���L"H��ọ�`B�Ҍ�c�2 c��Csn&$�!�l��l7����q�\5[��>Ȃ�g8��E�S�E�^��(�cV��,��> �n�+�q6�\�r�-	�pxf��z�[���s���y{���p�	!���pbڭ:~���>�o��5�e.gR�.--]�9�d�	_9c�z�����1̅z��2������I���N�<)�,�� �T����r��d2���Xr�h��l�j���&d��:���9s��6W~֌�q�ކ��+����Pw� �z|���A���~ayy�=�����^���%�^��Gl�b!w*�u҄�E`(OG`<�-e"kJ^�6���Tq]�l�bq�e�xx@JF�%X;�v���>Α�Ӱ����#�1+DS�e"6�<G%H	!x�/444<Å������TR&����x�,����L�e��@��͡�x6!
ȶ�^:z<���<|FV�OR�mc��
��!�)�Ȁ�¶n=�l[�s���)�>�� f���il�q<�CF)%jk>M����tS[[����fR̈��Ҋ:1�憠d��X�|��?��1�۽�+3�+�9�����fpZ�tnTk@B�t<d9-s��' ,G��*�i��e-r�JUH;��ĉ�8�z��4���۸q#�3&e�����(M0Ii=q�<�/\�5�r���hG�?��m.�a�Mrk�WБu���J���	���7nXz������8��h�<\RVJd��6����$/9�������+��<3���"Ӗ��� ]���/B}Hw�4@�P��% YgqjS��VHk��u%�4��(�e���U<�R��z!},��T�6�blc�I��n�N��և*�\��f�$D�K��9�ݵ�.Z��3L�Y[��n�$^ܒ���]����$ܟ˨So
��8�w��$�N��=���x����v��Q07j��s���6Y���â,f�,�|�*�2B*l�:�����NJT[�	�O=&ܺ��JL��K���EM"N۹k-O�\�>�B�� �t#�,���n^��[�Bx	G0�r�6����b^OtZ���yM���y�$t.�/K�f:teI��uI72�!��"����n�9L�z.\�����ƕNk��-=�X<$��|%�n������B_Z<��2����ES�#D'�9��QB!U����wk	d�@�7cd {��Ӕ��qf�ʜ)��$C�����MO����Ä�䫄!�0��;�B�=kP{����+������+�)�L�C������&�'D���PH���R��N=����)b�{Z?�A�+�C�'�o�K�<$9\J�s��x��QB��s�P�|m_8���ZN瑍�G=�\��q� 4{�⛘�0M���o�)j4KE�_��{�>�q�-��˚��+��@���˛�x����?�*�I���C
��%��x�~w��Vs���+�+P�թ�r�JP��Y>$W�ݭjaQ��3��	ӝ>���RtEՂ9y��3_	5�t�<��wؒ�JVӗ��.��(!���V�	��>���ϋ׾��߯�|�y�;��Mu������!��
�]v~�ҟ���4�aԘ���ի��ʇ�EU��u��~z��'�0f�^�<�����C;ʎk�>\ê�V�=����*ǰ!~��nU �SC��N��3��Eɧ�&Ћ����$2�C��
�]��-�3}�>���UolSݰ1L��9��]�+!�Z��Z�~�|�Ps�x��<���:Ԥ��NGsS?�m�Y�z?)��������{����`4��]�����c.<�W�w(=�����e�Q�L`M�W.������r�vD�cq���a���12Uu�A�Ug������E�tjϊ����Y��_.2�j*�� ؈�&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!��&D2؄H��`"lB$�M�d�	�6!�AvB�F�7^�c}em���cx��f�-������bRU�9d�2/z�G��(d���Q������lRH9���E2���i	i�T	L�_�=e���ƽ4����;JS�v�\�H��7wDs�9�@_V6o�[��5��ѼuPq~ۃ[G����|���yb�纮O����F�νt��=+W�++#!-!�K4�!eǶ:�G�Юk��z�ӷO����˟�y߆����Z<����^�վ�R����zޮ�:��}'���y�-j�5k��Ңy��K�������O���~�j���6��R��P;ɩ����ͭ��IΓ��@oR�P �@����'������.&�&r45�F�fo���].��m���X �]����ǜ���{<�:��C�z����d섄9�9�5��o���9揓�t���)S�й��Ǵt���	    IEND�B`�PK
     �9s[���HT T /   images/00941d67-c746-454a-b945-4fddefc776b2.png�PNG

   IHDR  Y  x   ��H   gAMA  ���a   	pHYs  %  %IR$�  ��IDATx��w�%�y'�;�}��oބ70�0D"�D��DR�"�i����z�ZU��r��Z����Uk��Ү�Z��%
L	 9q�3�	��_~7v�����{�(�5�>�77t���~_<��o]o]o]o]o]������������uٮ�@������2^��{O<��ߍ�c���ҋ��X�'MS���#?��E��d������5����]�g�]	B I���z� @B�N��R�R	ˋKԌT���O�D��o����r�,��?=�����C���^^^�r����k���R��
�����#�{��-�0�{�a(��z���鿹�����ȵ����I�.��2F�)�N�#��P����#���^1�E/���<�2�i*�lnO>�2�<�2����A�}�^�-m�~����/0�F6��L�<c\�铟w��;��+����<�>?g�'+c)����X�WJ4�ܟ��'��D��朗����?�m�&���ٺ��hx�Y?��f6n}�)�t}|66�MK��>4�|_}]ǃ��Z;{�+Vג��7�����j_ܼ��G�ͷ�x��=^�����+t%�wk�J{�}җl�i^]���)�K���{_d��}�x|#��kL�>�9�Zly��s�1J��UyT���䳡�7��%Yǲ�P{Sjr�}skO������_�v�����g
3���~��R�G7�������o��\��/����=�9a�� e�`�a�K�n�@�>�:�a��a�t�J[�+B'��9[t0��n��[�I�:��h#v�]zF,����o8�@?��u�<�p�H���������H�b��.}.� �g��d���=3q��ZY�Obdq�M��N�bl�H=(�QYz�#������L��<��NG6�f�o62�yȽ�F��c������0���O�j�B�E�w����a�7�����}�	�l��\�x,���_��+���&�#���I����P'�V��/m��>����LH(�o��[H ���\vV@��u�}�}_U�)(��:��f��d�Ʌ��������8�|�8���}��L�`1ֵ�	����ݫ�Д�@�	u�'��p��Y�����T���>�<���^�	�^ڕ�%3�"jK,c$�r���L�%�}�pB��L�$ ��w�݄7m�d<��;C�$܂#{�pM�Ix�vd���D������zAI�醹�k�Y1�8l���������SO�������쁥��g��9f�s�A),I�z��܄?����闲Ƅ�����kP����I��C#�"�i�0pk�;���L��ɗ�H�E���7�mHӞ��5�!�,2�lS���\�`��y��$��I`�y�s��H
�"SvhS��L��
���6�I	�L��
��¿�='���הIXG�l��� Ne���5d&M��:�i�5�_����S�~`���I�=�m�'�l+�> �>{�
:��`3u���A����m�g�b�$�S�߳�\`f��t�9�rڇU�$;�n?S��b�:�i
�3g��s��tN]t��D�;��︬[���|%�@���$d���o.����q����<j��[\�~/z,,O?,c�ڎl�<�=�6�$�
�P�[X6s\�� =�+p*1��,<B�?#r�WCH m�H��g�H�b���W���ҩ~�����`��-U6z~�����J*� %���%�@�'@wz���H��H�^�!H��C�{$І3s�&�����|�<$�����j��/�gЏe9{s�L��Y��&F�-�-
���/�S� \�o����|f��8�jK������~P�*�og��bQ�ʚQ�`�����|�]0������p�4�A��gRx6�5\�#o.)�D?ÛP���{i���Uty�׃�5m���m�&)��Y����Z��f��W�$t�RGX<h) e{� ����l-ًLB����/�@���X��
�<f��$�F_k=sQ�j�x1��U��0�E�:!( J*��9$��k[��:?gNc@���&�*P ��b��2P��ʾ{r����p�y^�x411G���11�&\�:V�#~��5k��j���,�$��I#��AY�n�Ma^2�qLC��UI�ZU5��'h8��6�c��>3��L����Ŗ/�d����t`	��	o��XB6>�îk�J��c�L�,�S�L$���i����b�>s�-�����d��9��=�'}m�螅Ϻ���.R3�����+�^?��d���L�X����c��IVbg��+���h^(ڊ��-f$���%g��5�K��B�黇ߠ�oʰ���T���ڮ���5(8��������̙®�͂7Cr��^���\�=���2?̈́㌷��F���2YƲ�i�D#��0c�b�6�j�b�L3S&�^�AI�l� ^�?���$���{�� ���B��0b�z���)?��<��Ξ=��R;_H�jx�F!�:�
JN�Y���Aԉ��:XU���6��Sv�
Ӕ-��d�W*c�TSπx@;���@�4V+�[�͙_`�rس�oq\0艱KEGjs�	�~����g���$SoC6~����2����ĉ�����Y��tQdRn0���f��t�~g�G�_^������	A���� ��A(:i=�,���g�< Yx��dU���K���|\��U 6P�.�[����Y���z[+��M1}߿x�]�s���f��M7�\��5����XRy�
�@}�p!3='(SS�l4c��.�y{��8��q�5k�lŏ��75�^Nx�����W�����0� N����/�{��#�Z<'���N#�j�J�TBA��/(��lH�M�C�VXMH�j"�� &j��n�Ƀ�_0}����`C�S�z�J'�h�rO�UGJ��f�����]���bs�v�7��?�7�pf���[|�_E嘃1�Q�/e�
�"勎\�e��ſ���8X�y4�S?/��:͝z�~;w���#�Ȩz�c�Ne k�l�'�3!�rWZ�G�2T�����
֙t�G��9�&�q��l��ɭ�Af�~b���`à�YO��'�E�q�x��� 9��Ƥ6s�2�J�Ӵ�<�r���o����$��ǥx��F�@���|�_��+!0���mx����@oIN=��j��h6D%����F�^F 6ߒ':�|_1+Su��Q�	/&�ٔ��%��Z���X��3�B��2G.��s�;�2�]�]�⮆Mx���Vf�z%v�&E�bɏeVL�ժ�CXRb�}٦nc�0���;�8Js��xM�}$vw1x�v��p���6-�>�l�
8��=� ��5: �?S�p���}-g����@Ș�
O�����N޽(tG�)k^��>�����9��*��T�a�S�p�o���[is��l`)��c`�l�^܏�o���0Ꙁ+2:������en�,�p�)^�T�XX�B?qB�����ڢYH�<�5�~�3�Ǫ�%I
�z�bS���p�K��%�_����W&�ݚfU_C�rpO3�Q��n�e�q�8����&,�����(�J��w�ơ7yX�?��'1��OKo^	kĠ9�0�;���)bƓ�d8�W����P��h8�Q/9��8�6����U�8t�� l��d��$FD�^戅 %v	��"�Y
Xz=!�cCU�S1/�����qI#d�bd��l��s��F3�h=�F��0	�q,"c�^�{�ڵh��XZ\�XI�%VV�"
���D�������C�u�n�V�(d�⿷��Xl�9�ɕ��m~��0�8��~�:�˰������M�~/�
|@��"9��b?��rG��ץ.��gk��X[K�B
}�Y��$�� ��>�H������9��!�q���(b_�#;�,Y�_�,/��8�5߭���͑�-�
&��������1�]�-�PG��D�/�T�©��wD�m����R���P��y4�.i�jf�dS(v������N�+�8?~]�X1c���ygFy���H,�,P�QX*���;r�V���#B���q���� ������0�\±�fI��q�:�r���L�q(��D"���Aq7�񯜅y��X�/u좨�ɪ�1waF���N�2	���'�O&���u��m���~��M�����f��Q��B�
�(����,N�3�$o��Uë虇߁��f���N8)�v�wN�F��	#	�	\�2r�x�uL����k���>�1n�9�������[W�Ⱥ.��[�4�;�Y�$?6|�T�S�oh�9h=P��×��%ոo�����Hx�h`����{'�P����B[uLP���=#��	���r��8��
���͜�^���Z�-2��s!�����u���{;!���`���Ee�k�zp� kY	����}K��|f���!�����]��>\&��S�a]e�&�vhCQE�B��|���N�KM��l���&aQ9�*iL;�*��6MLa�6�o��}��˞�,?����i%�2u�Xbޙs��Pn��H� �tFsb4��J��ë�FXV��Z�hT�z�Ȏ�:�7F���3i�v	���Ҡ��plaG��X\�Y����,Q��-��F��X��G @W�<q;S���Κ��9q�Y���I��y�ۭV���^�mI��y�~ �e���6����'p�����D7|��@h�A�Q�1��j�62G��sD[[#C�ω
��Jh�J�$��j���f�cU0�{�CehTcK��㨓fG@�PM���#
��u��S)�#	��P��	4N�%�9[/�ą����0Q�Ӱ?U�u�B��4���>�<�@��gp&!*���zG�)����%�F˲�Y����c���̅�V7t'B��]�D�玧C, ��T\Щu4ih�qBS��{/��?����p�\�q)Q&����ҿi9V��E�)�'�$�\e�6�B�8;�X&i�}���.a3`�X�Th4�N��������ve������2���P4I��ơx�v}��B�m���	x�gY��
S��aD�WX��4�>`�G�~@7����W��bd�L����*§Q����Yab;.E��Хuݦv�_�Ǒ�sXUo�xo'ZsX4]Y�B*��KI��a"d>"Z�aa��L=cs���gXZ#-�VF�ZuX�l�e�$�L�*F���S����5c밾>�ut����}�����Ή�f�$�nK��+�G17�G��g�4�-��=�k;�l	�K]�0%	.IhW,�`�$ˊT[�ʛ�JG�s���
���K�H��+I�L]�o/௞Kd*�u�W�Ձ |uRyA��K��m�b�M!�5�9qq{lJ�EyfÿK
�(��O�Fw���L(�a����P����{-�<�ޞ����.8ƪ0I��i>/y6�[N8��X7)���:�ui����ת��	UM�U�� f�l#?/��MYiO"a�u6]�y�W�l�K!�AC�!�f:����~�{3��ܘ|��y%���}��2_ �T�ؿt�j�L��i�t����:�B�w�G�P�ב,�رbq�}^�M�F)�P,H8V��c��G�S��nf��4?�P������&.nO�*TUq7)�#~'�ᗲqh�t3�k���J�|� �b�b��?b˘6ul��;6]��S�I�b�T'l*��*�EYRM%�aUu��Q\՛Ʊ�^�p{�O�|Bk��\ԯ.��CX��J��,�P�B���#�#2�N	7J�%���p��f:y�y9-a"�ccT�-6���75��!�IZT@��Z�C/�;d��$��Y��6Q/�09QƎ�I�����ϡ4cq&�`��$	��h�4b�XS��ifL��Zr9ۜ���Ev ��2k�nvi�����;U���y������}|�o1�#�a)�f�c�6j�*B�"3fI�����g�ϔh����	�н��,L�&�];��j$�XJԞI���g�Oʴĉ��r�نŠyP����)*��a��Q�X����l�L���a�=�����_PV��%�3�x�8��C6Ѱ��4a6Dmh��n����|��ʬ���)q)��s+�7�
����S땷�+��q����x>8+1,�M��|��Q-)uc�����5�2�������Z���HB�b��ȍ�xL�Ar�zs�@�^{ڢ@�Vn5(��<�ٷ��u�j^�cӂ���	�'a�b�9Ml3MG��e�H��K5'��H��/P.UQ��`�eߡ��f�wM���SW����h�j����&lT�K��Y�2=�N�=JZ������1�i�c݅q�v���a�f�><��C�W���4��]� C��N�$�B�p��'+Ɔ]S*��_�%��+��>�;�]�-$1*4���j�Q���N �U���B�J4;q��Y��gp���o^��pϜ}��bnV����{]Z��V�[��y�z>�n��j�6f?���^��M��q෷��\���u���^��2��#*ԛ��u�a����9��.�]V�̀��[����XW��4gU>g��s=o��$|����xV;	�]VQcM,�Fhq��gb�n	��m��l";KBhؤ�����d��:'`��v�	b�J:1qH�;�,��/�Za�:&N��V�	B�v�ռ����Mng��S�X��
�pTg��yZ��P�R"�OU�g�F`���
v�m��=RWKhF=Ǿ\ё\=R��@1���uz^��Q��|�ۢ{������$J|�+uR{Kb�Y�[hQ��pf4��i�����-�MeR���ch�14�ϟB�qV�M]�U=g������o�;���r�������]f]�=���@����lF�Y1��"5_d�1��5é6��c�N�xsJ�XH��@�\�P�r�R�Ѡ>_Al���W㎍Wc�6�0��="���V�-d{��>+�\D=2�U"�Ul��c��:<t�U�8wH-�ؔ4��0�E2"yt��H+�X
�iW&˦��`�$�ڼ���L�
��X�o�S+�{ltu޸JXrf`ctO5v���V)�2U�x������û������&N�d�[L�tmiNp�J��IX�	jZ�.�4u�6똅�}2��a�T�X��͐���=����K�Ь;ي󋰨^�7*f�֙���8�N���[�����=/������W���P�j%�~�g�����'���O�{����D*;�
s�'x�PHQg����mۯ�:�P����C��f���ZE�j�Z���$�W7l݉����^�3���$j�8�T��ڎ�>֕m���n^�/~��X5��~?��O�y'w�vא��B#n7^���Ч�n��W_Ʒ��X�J�z�c�kO@�����z�����غL���#�}� ���;��;p� }�]x�5o����{�Q�>��6p"�n�֘u�p�τ3�p�!M����4��ۊŹe|�[_���Ӱ��cW���u�>;AL�7?�_��Q������)^:~ I�mS�5�D�J���l�.wR|�ӟŮM���3~�̣��w�	ӈ�RW�D�X��~��{���Ƨ�?��w�G�^��e�QJ.��簃���yx5>������a��=x��~�]�\2ˣq*�hL�ٲW]q%!J	{N�����t�U�t� �Q}�snC�D�-*ב�,Q���q�����-��M�bUi��MB�3�_	(��0(@k�
\��;ilF�@=	1�Q�Z�=�*�k�`���B2��-1� 	Ϥ]0U��L	<�&��&�ъ6�	&��\Żhq2��Ҭ�5V3��}�5�"]j^OD&<���D!=��Re��;�8v��xwnފN��Gg�@�u��]�L���sꆳ�|T�asN���,�g4d#��?t����_�u�m�����&X;�[˰47	x �oc�Ċ��ۭ��o�@j�M4����[�µ�qd��{�Y�4$0�]W���0Vg�U�6M�fm�m�v�*�w�R��;�=\7���?����f�Y����+��(j����t�� �c�&���|	��:�kx��$��Fj������P�nHر��-x�U7Q�G0��q���8�<+Ql��,X8�}�m���ke�*$����ô����:�l>�����{1o�׬ߌ��x�6���N;�E�䡕�s.�VKh�O��g��e�]-	63�=<��%BC�8�-�3<�Φ�κ�z�4o�U޸~;��=<?��@DL������z�.ܲn'FH]��Օ1�$Z��������1���)�vSHC�<��GV�=���ľ�_�Lk��G%(�����'p�밺>I K$j�5x��g�xE�ئ�o�Ud��Y�YPr(��v�w�z�Է����?��s'�L@+fF�x�X�h���ny?��I�=�g7^>x���Ʈ$"k�c��� [�u��dJ" ���� v��Fe�ܐh'6}h�<��aX/���r*"���Z-�ar: �۴��^A�=C�#��^Y��M�&-e��-�N|�<��Ӌ�B�;�j�Jx��\��
5��ư0��F)���D(�� �Y�_yy��� U��7l�^Z�g����o��e<t� �s�`c��lӲb����o�����gC�#|}Sv�y��������9���_�iܹ�~�6cEY+�!�&Z4Uv����L�����X �G�X��P�T�vY��]a�+�>��l�����`/3��ՍQRoiA�ʴ���g��v��ZKs2�aCF ��M�Q	��U�T��{������X�ٲ�(|�_bK��E�&fU���k�}�F����?�bkmfA�.F���v;�y	�6l���)s�8�{��0�E��<���s�+0���K��ǾAj��7܆�k6�p Qé������Y)U1N������Ĥ8n{<�>�m`<��Ȝ@��5��i|���0�1GRs���/���n�I��fg�m)�_��e�i(f���I�޳��^x�_N��L��9������qb�z	����m���#Z-��8)��#�F��	���Z��o/v�aO $���BsR�uS��[]ç��%?�>ӑ��%Ly���\�][�VbDkz��,+�RF��$(B���"591q�hڀ�X���L��y�.�ad�B/�R�xg��Y�i��e�q]]6�0ь�5�����pۺ�X8�@!�B�N�����9�u'���*fI��v�)j�*[���r�$���U�q�vl�M!�Lh�;���A�<��-�Flk1p�n�:�m�;o@���1A��{�^K�}�;�"���}F�V&C�m���q�b��A">�+u`�+��9d���g���ŊW�<3�o8&���-�� ��{���Y������ ���<o^|Õ
	:����=X�҈��F=��c���jb:۫�"����X�D�)�Q%l�\6�������w�p;ݣ��+���6D���v�^K�\���8���y�Ώ�N6V�9�̠�=7�� ��w;,�����T�2���!�\���)8~NcqS�ý�����(6n�@L�4�R5�w�NC��6�~�q��A�bK&P��#�	�l��s��%�O�Ƿ����M�o#Cc�qE��u��*%������=2<���zH��hE���!�Si,y͔YO��a'��:��ʂ%�~N���OȼqV���A3�l�kY^x�]=����(��.�ûn�]<�e���u[��d�>56Id��4�I?�(4�X"1�%M0���L6軫	n_�;6\�1;&�Ĉ�N4'��Ma׮��[`H�����^��q"Ji�_Mk���4��IK�.�h�-"�Ȋ�;�5ལ�%����OT��1�&Ӥ�ݺn;1�����DC�oL���&�ę�t�%�Q$��hc��n�rg�Ԟ.n_�O�}g�hF�,$�xv���kq1�ƃ��8o��m2�i�54���m$α��
l��]���q����3�<�-�*Y�9����ׁ�U{��)�av�a+��,-��%����qU����^h�ToN	Er��{ZSxi�����"1�f{����j����9��&����
�7�i+{z���lm;��7۪�^b�u��1�v���X�3k艹J|!1Ł���VᰲJ��=��ĊΞ;C��I���TSre3}��/W��MF\���F�6%�{�\М�����+$����x����;߰v51g��vN$�ܹ�aX�+ ��R�	۲9|��T�׊�/�}�Ez"�F�=�u�^ZV3@�<��)���,I)^���N0���_\ą�XG�'Ǡ�����Q��e^Q�ƤIs��m��vq�!H4�ZD���-��V7�b��5V�U�&
ͻd|r|{�����9	
��uCX�qd��5@��q�\���LI��Yj׎�ոy�j�ZGMM�)�W,Ɖ�,t��ҥX�ɫϐ�V�$���7�Ds���n�求������V�+�4�	�^�@m�Fr[c
��h��K%	�?:,�j��^�3��0-8���F]j͑�RŖ��8��A+��ܖ0�x*�6o q`���Ϗ�AC&��\��c99'�QhH|��S<h^d�-��A�u����N���8�L�o/X��GZ�B���z�{�#�/D�>u� ?�$*��ĎV�I�҄-C�$�}J\F�X�$
�2�r	���j�!b�=U�͝�"���[򘇑T9Z\Z���]W�F���mW�B�&e�C�Z�9T��4���ʚJ��< �np6��B�J�����[��sq���ӷ�~�L�=�jJy�R���6`N �Z�,�bHԆ8b"HZcg�g5�6�u�í�4;wi���g/̢M�Î6�D<F6u	&����r6b����0��9&r�ըq$�E�V�H���9�,,/ӽ!��&�V��e��S���NzB$D���Ks�G	�i��.1DC��s�ª<iN��S���B*�>4��c�a��c����"Z�!`Dwj�j?�S+dO)�"d��i��h���*vMm���5�fNQ
Q*�L�	�7���t��(�Q�bM}�'����
�2��W�>��ׯ4�����ԌR�F�\$��	���W�u�N��`�����	�z{���ۯ���xa�1�4;h&]�ʂ����$��4����r�={4^��<�P�o��Û]E�6Ww�l��Ίb�����¥�_��N�%����������i�v��j�-��'����w�;7_)�!'�����,�N8Y�d]�u�K���)Q�����08z�JI6��0ݻB���1\v�*��%��f�W��:��
��1�,ժ��+��:}���=X�>41J�j�''�!�(�W�坸��a�굱�m��]�cc����s�T���Z��:y���\�$T�~q7���ӨՄIr�.�5�ۓ���������bs�DN�YʪZN�A���J8���PC�9ޛ���K/���q��KJ��0m�7o�֍[�X`��O��Ҟ�nj��[���l�~)������@cq��Y<���4�1i�ma�1�	����5s7i��7n@���۩�:l��g���������M�&�X�-�[˒��)��(�ʡ�q�5�fwͥEZ'5�8[�����z�	�P:��9i�Q��R�(�F�&l_������<�
#x9Y����Ah��lr&���)��Zb��b���:��	�J�쩫tR��c���B��A	�=Վ$���q����p��ڏ�s�}UR��4�P�<�,�J�������{:<�ey�@�=�������" 2�������<nE��F�4�W%Oz�xʷ�x �4	h�JY͇�S��b�Ө���xLNT�	<ς�3ȇ�1�<x������?�~��#�f�b�c�Nvr�ví��/��Z��殲㫅�o}t����Q1�4ڌ�	H9�'(a��cx���q����B��.�HsH�1LNOa�U�		�P/$õ-8�1��cG�d����u�V�c֙����#�iR��{�[�!�Q4��v3�Ekg�f՜a�Jٜ�s����Â� �t��}�\��e|��{����HI#k�-�eiU{�]{��o�6m䒌��7a�K�2�kK�2t�$t�GL%t����^�a�,E�}p���{�#�L̟�?GRԂk�a\�};6�-��	DiB��T��!6uf��i��E��ɺ��-������:^;}��C����4����_��}�W1�~�-}��i��˰�FguL���D�Xe�?�p��XEk�W�����$$��ơ	l#�_꜆���zw����Y�����~������S�(��X�p�����҇k׬��}�[C�*"�7+4�]W���慠�nC{{� 8k�N���w����Zs�,���`�oks��6h�,2��ݕ� 
G�܁��g�~���(��4�{MD�5D�2y���pxm�����H͟����ǎ��ד�?�Re�nm����60�+!�=�����U#\�,�O_z
seږ!m^�@���H"�rh�̝AB���G���2p���O��}�Tr�߄��������Y�15�O���b�#5a�l����j�����~$q�%b0����8q�4lU+k�}s��_y)p�@�_L����!,��YX¾So���Qm4��N=N��V�z_��"�fg�H����bgZ�yj��nRe�-Nߥ{,8w��Wp���h����eTR=#�l�Q{���/>����8q�v��
���sLf�����������R��[���o}/�z#�cx���P��Y�1�EX+	��˴����́3gqn���������qth�͑da!�bf^s��dS���O��m���-�c�����chV��s�iJ�KZpy�B�na�部S����G�� �\��x8�1JL�X�Y;4�u�1����N�����3��ҐN����a8J�&��`��Ԏ��^���O��y���E.���B�����m![�^��i�U11:�*-���HP���Q���oH�����XL�d���?݆!0bS����8h*�����]�,��?8����q5ˠr$���'�����	��_��]%i`�U 긓oy����_��&�/,�� �?5"vĲK;����R*�����y�����^U4JCZHE�Sqdɨ;��w�a����/Q�yj3`���2�M]1���)�r֒�[���j"���l���,u��t0:2�f����ԫ(�+�����9|��@���E���^w�rs蒜�[�)��ee
R)��$$��#?.�d�D�
"�E�.��pNv�pW�.�k_�z�T���Q[5J�~	���` �!�]9a�Ͼ�XP���?�G�牍�5�����#,��?���2CXXn��f)w�YzM�}ғ�eu���?�J��q��ګx��W4���r�,�7�쬁{x�&�ӏ㉧w���%yax���S�h��$p��lG�uʯKt��1���+��d�'5�Q�8Ҥ��g�u:m�=<v_��_s���ɑJ�8e3�QB�a�Y��b�%K�U'�vx�>^V��f�bF�e��g��܉h�'�9Ӎ�%���1��*��R+����8q���8��4Hm�Ip�@�2v��5#���:1Z<cURII"�����;���HX��Ͷ�uś�Ȥ<�/������������f`nm����|���h=�ꡕ�g��_����B���2{Z���7W<ͮ��W+59w��O�{�T�XO"f�u�������+�E|J@��Qi�Q�]�a��x�9�_l�Γ]&��iw�juHm���,�T�m����lj�Zi4=7&Uz�T��{Rb@e�5���V��z���gN
Sb���,�ʽ��!�v�C�9R��F��.�LӬΫ:S�&�����]ȃ�K��u6y�psxߪUS�Ukx��q�=��u�i�?hTl�&�1����!G+C��p�M�`�����b'�vZbC�)�%.���+��T	�,��=�'��B@� D��8�������VOye�>���.�}�M���ۨ�v���B�� &��.<v8���pav߿�8s�$V�߈s'���1h��)��~�p>��0�7���TX��M�I�	ŪTIT�*4�-Z�e���^f-��g������ձ�R�-j���IDLk~��ɱ�4�R�m���%Rs�u�a��x�'�RW�C��/�Z���X��e�6{5��`P���Е��"	d2/+/W,2��X�Z�,v2V?�d����H�4�[ꁶ ��� �v���M:�f��W/�9W&ﲹ2�
�	��}���Vk�
WU��w�_�įb(�S'�JơURFQ��դ��/^s�������޽8�p��'�t R�:%�Xq����2e|�3_��kn@���i%eչ�L��:r��3{_���I��E單;����t.9W�ޱ�m����e5.��e��@���n�E����j����~�����q�{A�����l�o&�t��,�:	>�������i�1ʲYw�<�[�s(�Цhcg������������N�sWX�c�at]��2VI�ү�#�ظ]��.j
Mɗ��C�8����<^���5f早��?�(0R��/)�)SH���$��~�c�e�;`\j�D��4��`����d�V��s~S���������5����u��\$�/���^�ݴ�iU����>���5�R�0"jl���r-i�^"5"w8ځH�}�?����["�$rå�g�D5S$��L�n��F�83�����\�K�N:g��V�B5%���!~��T�u�Z� ���R�3�6ԙR�ަ��0���|]�����J��LCw�:�J�/w���r�,�)�]��g�-�U\�I��41AJ�;�-���j|������L�Y�:n��7�הQ�;IA}/+�G�\52�*;�8��\�5����/���33�X���Ն��\�ջn�r���_�U�^���Y�b��|���PbeZBn8��:���w��3m�Z7�8'vŔ-35�0�Z��׻��GbZ;16Ѧ������Bu��x/W#�'seM:���GW��!`���Uڱl�v���
|�H#�HV[���� �$�Hc^9ӊ����o�8TQ����>r���+/�]R��f@���~`�GX���j���ɩ%9R��s/ՙ���m�AI��#��7L����p��.afZ��E�����t1��"PS!Q%a��r͕�T!ɠ+u�c��w���[U�g߹�<��&�|tIЄR���5�|"��8�7���*l]������hHk�)��5ؼ�HP�`�v�v�!��FU����4�@"#��}9</0�V��N��a���r�dE�h�)��l�V{zL|n.5#��:Q�ρ� M*:Il6�r@uY�Y3�)K*/u/��s,v��n"��z$-�����Nߓ��ĝ_����;���E�m��x�5c�����)�3b\L-����	��3�[?`R���Wu/ra!v��s���gl͒��wh��Z_�2�#��Z܆���*j'�[����lݥN�;!���|p6Zv��H�+���td���B�U��kCW�T6���DbG�F�+8�Y�-�l3&�oR^/p�$��1��34���ȎD�u{�����T_���d}q�ٛ�뀷!g��L�d�Ϭ�������Ie�K�k��z�C��n�\�P�fʺ��&�'V���éx�8�5�g��!�V�x�Y�g�N͞Ǳgp�UoC��a�Ǿd�������'�pv	�#$|x>Y���B�d�*�� ��R��ѦQ?z�4vP?z͖ؔϜ8�m[��Z.I������H��T�9Zg�G��OA�N�׺�Jp<�H5�J�d�}��z
]�L5P��؀h�Ky��r`�9�)g
r�D�S�9��a%�����ZeLĆ;$��\�qǡ�����y�f���m@���x��5�H��xƗ;��g&Jj���r_�Dj�҆�s�,2��%��[K1�e���L�vN�5�ƹG������$��4K�3�\^߇W�^����)�rd]$�+19�\c�|�����~�T���8�����Ý7݂��x-�D±x9����2-B�{y����Y�0���Φ�d'ká9j�=1����|'�+�3鶻��hcT6��7'?�ْ3�8K��k�N�V�䚂�+4�@��o~�(���arh1̲��V��#�j˕�4�5��]�7A�j4$Vz�����Z܉s��r�Q�䩛�;tQEO2��|/��*&:���M�뮼
��%�4,t�f��xdMs�ҁ�X�l�<:�G�
���	�Eu��p��Ɉ��0b_C�p���w]�5���ǝ���6uhM?sF@���WvZE2��V6Z/�'@b��ݯ��]���М_��NB�8V��_cz�FZ'e�6H�$#'!�u[8p�ޘ;;V�S4��aW�?0�v��.�ٳOa��i) #�Ks)�	���f51:�Jȉ���8m�M���4h%1�1e����	��!���e������m"��4��)��5Q2�e�A�����p��VTN��������q��7�r���$Fch�[�Xۮnh�\�"��d�Uf5
~��G��/n�Em�CV�p d�2�V �AP�U��V��2�jx>��%�0�,*j��� ��'"0s���A�rs�&vޏo��qli��A���8�_l�Q��
(�Q�O��1�������!S��56�߈w݀��C�j����'m��\�@��8��Z��[jX��ҧ�6L��`��<���2��ȷ�ۈ���AT�e�:���G�$��l�t�?��,���iHۙ7G�8������q����n�.�`���g��i)�Ȍ�b(	)!i1��:����R�����>hpa�  �@�^�� {Ͻ�}���Z�^ a�;�lí�ߌ�3`���H�O��=L㤅�95�ġv2�x����	�B��g�$����3A�mnǸi��0>>&��t9pZ�U��&����{$�UN�d;�����W*i�@u���Ş��k�n����q�2iQ�ܲ��{IK��f�&eZ#K$���U�BS9��́��	��Z"����v.�H�B�>���?�w$O��h�o-a>�	SJw�K�01�p*�x�� V%�m(�
�=wFy�š���rvJ	�� >�`~a�#�8�� G���a�
�J�����J��dW�2ֱ������X\1�R`�6��`2Bd�/2U��!�\5?���mg]V�i�bR�j���p#����[=��WX��Dm}��q���O����qӺ��hTEs)W4���J�-��9�\ȹQB�ӥE�E�����W�3�eܰ�F�K�- v<b!K�<^z�e�s��ؚ�3�b�����03��DM0��z�Ya��[o�}߇p�U���VĦ�����w�������ïR�"I�����ƍ�ื�bM=�H�}g��R\������'1�v�F�)p��B��G_ڍ?��c�Ǧ��T��3��|�u�B�je&9�ƈ��l�QGؖ������ۉ]�Hd;+و�6���"�{��������Xg�����XgI�%ͅ}$:;0�	�	� �E�y���/}\O��������}<=?�o�/~�؃8ݼ����Z�87�
%z���+%,�p��U$����;p������(�߲�j�g3�;y
���񣗟�9���R�U�Bk�X.�|[��s�eE�'L��.?��XoZLd��H�m5%���^|�j��]�,�4SQ� 'r`] F���R��0��3%�˞da4��Ǔq��I�?wB��+��z,��ک�B������So���Sce[8/S��l"˽�l��}��~o]��b(Z�5���#֭�N�T`N�s�A�m���Bb";�m���ހ�|��XC�u,�\	�*,��^�7��M<s�Et��v�*!��ZWp��p����l���,�#Y>�?12���s>���`��zb�U9���h�;{�{�><���h���̾���z�%�n��?!��q�|�/Z>VH���26Nm" �ϭ����D�u���Mq��1����x��Gq�;�N����u^���jYw�|��e|�fF"����ھk�|�?�������a�s��K�=L����&��U�i�#�ڒA"�E����f���8�J4���Ub��^�k�]�O����HM΢w2�E�X�s���?����s��I�q���Z�b����V���g�6;�	Ɉ����߆����u��²s.�\tI�����7�ґ��(I˩���E�f�&���3�8v��grۚ]1�]����EJ,��a�zx���!@�ş�G�?�CgN`���I�Rp��m֤�� �#�;m9!�S�g�mo,�`��TH+��B_�2]Y�y,�Is�F��K�h�91�5����g99��v�mx3s�
�r�� �8O���.c�F�#�\�̂�CS���KR����,���M�ы�XU�SH�q��A����(�I�g�����B��J����L��.o�l���z靤t}�H���x����{�/�:5��^Y�r������6��ߋ�~�?c��׉��p4��UQ����?ZH,����ԫѓ||.�`�0e������w} 7]�6ڜU�C�-7%��]\ăO>�>�8}�TY�P3��|TJ�	���ԟ�(������0���]�n�Wo�5v���b�!�g5i�=��3x�g���G� 9;;�����r覌�3~��p��D���J����~>��O`��F�ޘ1�h�4������ϟ�+�_C������yمv���Lf��Tߎ���|j�x��/|����wb�!����S�q>p�0������Obfim�7Iٝ
j��L�;��g9�>�vYn�A�(Q�b�:�O|����?����41jbp���>u���װ���m��za#��䀋vw�g+,�[R��Tz+-wq=�S��	�wc��@�\�ZL�:�R��?�{��~V�ʺ��#�A�RÖ�h��X��c�P�V3X"at`�n�V9�����)�L�$�9���8�<�nI�HĹ[)��)�馜Ke;����f9�8�SDͧ)�Q�YL��[Vrb����>LMO��{0����ФqT��ɡv��HL��9���hjŗ93�'��K���k0��\�v�v�a�jFj����TK����ɻ>�/~�����ŕY��S9��᫝�(�����Z�І�����c��V9*ÛHE���ԴmD�3�=�#��O|����1٘�c���r�-����ž��J� g�0�Ͷ�]ږD H-�D��H�.�Vk`��L3Qiu�[ߏ����c���1�r��Q2У9�U�V��0�iM��������A��̣r�$̫���oRk��_Oܾ�z��g~WL�������C^	��ҽ�F��e�z\w��]�N¶��/���2�ݮض�a�
7�.�V���]�7&�[�����I�/�D#5�>�NGsv��&�>�y������n�s��t�
T��"��O%���|��n�@��(�;!VνⱨV�[n��w܎�������S�����}s?�d���.~��1�����	vm�ZJr�q/u�%J��M�=�&'������eq�=�g7�v���\�H�I�p�٬��v����!�u�5�#K�I�i��
�_�K_�u%��Y��깓8����ôd}���V�x:��:�Q�:�����;����W_�@�A�<.�`]\��E�E?P��,� }N�����q/�x�Q"�{�=�I(�Xe�M�@�o΢Ľ������ ��Ѝ��rt]�9��w�>�G��Ϲ��o���`�yJ���J�5R�b��)���&��%	7��"�f;��؆�Uk+�����������N�u@��s˭nNf8�RbƧ�Y~��Ɛt4`\ ��}�;�n���[�@��i;U�?x�g����+N8.���51���@v�5{�����׏Nb���d��Tq���.�\p�Νk�5:2��:��_݃����,�9f1��o .Z��+u|�waz|�����g��SC�)�F��]����L�>�(N�=|�4�q�=��"��,X����Q��"��j�fܴ�ZX���A�\ە3-ݺ}�u7↫����Dly������ql����l��T������Y����d`�X�����C )x����o5�mtx��/�|p�۟/\8�cO���u1�p{�k.�KϮ�����u��m;I�KDJ��jM�1zֻo��0n$HH[�a���$U<qq�ƙ�x�p��mw$]�KZM��y��	6�'P��$�ݸ Mo���qlߵ�o�����]\���{��	�M���u��Q��u �Ҳ�8YhA��%%�M9�&���\STbgI�F%,�m�=R6��6:��ɡ%Ia4���[�d�>�:|�Vu�Hl!���)���~L�f���H��M̳�b,��������R"�:��E�j�C��sW��j�cι6.Pַ��8�~"�R.��.B�$e��pjI3�^����S�^<rⴄ�p�+>s��j<0�Ը�����R���<�MB�j���WY>V��'k0��]��z��4�>�O?��ԕ�����`�Ԥ��k\������R���V7�_�7)��
�s%�� �'G�k(l�8!)Բ�����,�Q�~����Ne=b���D�j��z\6����Lf�HA�D6j��Je'����j]�ŖK{d������l�'�8��%-��VX&��z�2�4���|w�T-�Ҩ���$���k��;�؉�/ϊm�ג�p�"$b������)�Iwf����#{T�9|9(u���$�ɉ1�D��p�&���d��|�ƮK}aç�r�m�lbzʹֽ�cs"�
	�����Q���|	Ov� ���{��z"o�
ڇ
�I�O�h�w�h5ak\���W��bÙè����r����eʾ�yd��: N�|�=-��nȼ�W�N��xLu�'���r�V�u.ZDԭ�� k�	y��M���: 顋yR<�Ν�4�sR,��FT�e�����r>Y��"0X���)����v��c�N����V�ݳ��
�l�X
\��MRa��xp��̋om
�'���7���
\|��^���F;���JŢ�Y���3���c簱Z��E�<G�ns�^oY�a���̋s��t ߟ���d�=.�w��i	\���&�<Ѯ�]3�p�83IN�d!��)�5Q䲛|�]�S�3v.
�S���Tö
9�1Β�c��и�8��L{���MR��}��vP%RH:��zb�"�\�o������X�Q�GU��
�������sg���Ú8jJ��S:R�&�q���uz�dG.�sj�'3[�����eRX:N��j�-
s�,&+)���T܄����Jzh���sܤ�V����L'�"��%���t �."V:Gc[F^�%�~����99��m������]���J�9u�A@��l}W���ƛ߂DR|;�Ox%�_ҕӬ�Cg�����E��ĵ�,5K2K�����J؜Dk&Nq�4��N�v�� 漆4"N�O�uk�?;X$�B۷>�6�,��8���!�+��//��l�+��M�_�c��J��.�P�$ug��L�&��bb�d�&�d����9���q���▬�1s)�$#�`�ã���=����,o>�w������x�ş��s3�j�S8u�HsY]=Q{�F�*^�FX���9��R�+��7Whr����������3���1�/
�������%I�C=jH�e��to��qMNNb�x�ˍ�djq����9�v��F|�����<Ԇ2�ä�?��nL����<�(�?�E��sf���fZ���w�1'^�k���V2�������ɇqvn[�_��<i,�fM�]��9���H��Dy�J췂g^܍�x�@�*�������"� ,R����X�8Nڨeγg�6W�/Wh�	\���-I?��Շ�pb�<�~�%��D�E��OYs��(>-Ey���o?�#l��O�/���;t���)���	gSBH�?v�^���G=(�pƖ�ĥ
N,t���M���=�M��p�*�'����&7�ٞ�*Y ��;33�=o�.�>IDp��D���E{6Ѣ.?z�a\��*]��.���IWg���(?d�3z�=ܤy~�ŧ`j�ד�d\�u9"K֨V�� [ZDB��I���{���~c�'��qN��ʊ+����7�T2��5��]/\�|��ɧ��x?=�
N���D��6��5[��B��*���b].��]�TV�B硁��2^�x���*հ~d5�*5Z,ee��r��Yj�l� W
�`SC�]I���gg.�g��έ���p(^�+u/˜e!e��V��bp�LNU���YS�L�wo�6����#����;���l^P9������݅���{\��υ`7�@*U�Z�����v,��.�4T�E��N�ڒ�q�6�Tpt�4���`��*L��)�2 us��Xw.�vj4�q��cRk@�zt&����y���:����!�Ā�|�i<���RCV*L�Bو�ђ���#d�!U�xk^�,�{�K�,�[0��X�/�>�̱�x���P녘�X;�JTlΒ;�4Gc�s�Ԃ8�G��Ϣj�Z�ͅ8
���Hj��s���5T11<�V=9�?T0KRV��Ӄ���$��S�����:MM����HU5v@��`玫���������� I�6��z��c�Lr�\O+tq�:�\�zm���0��e-�ޗB�%�=�����j|��%�Z�lחet�����A��t�Z��{֢�>���Hz�d��4FWKs���e�z�+|D���`����7Hq�R�&E���?��;�Wޞ�C~s[��TH�	H){}~?>���X�8��-�/P�#�7U
mu1d{�Gg'!��#�a�����זϢLz�U7c�'��J\	O(>�eə�V*l��VR�Vy3���m��p�-׌��/?��HV,��진+�s	|VG��D�tf;;��y�����6�-T�����2��O)V�S�� �qaa��R����2.����g�u�V�}���|�W5u�S��ha&��t�:!1����9�4���q��4��G���/�TgQJCv�*�R�Ff�e9	�J}�ER���s8t�$T�ܼM�`�8qɺSgIݦ���Ha�"��Q9�" .�&r�(ض@]I�H�rFN�߸j֍M�	q��a9K���c���/街|��R��Y8�ܢ 3�B`�-t'��17�?��O�0?>��B_���s��i٪a��}��'�߰����,l��F�s]b6և��z�Y]\�Z��ԾMS��;?�k�]�C�����sI��1�Zl�&�X���my��ɮh\��+�e��w�1�rD���z/f/�g%;ȆH��^��������	7b�-�b@��'�Yڸz�Ԯ]j7i�X6'�=;X�θ�2N�����%�h����%N8W��.�֨�b�f��O� b5����[�.�T�E �W��6���b��jGZs�s�65&��5q��il۾c�c��*�[_�Ɍ��8���q�VLf<�<״��?�{��{��Xc��Mri����O\���K芝���W_S���iMڮ G{�h�'X|-��ۯ��&6`��Ue=iV�����A�6�R�+�d�+�|F�k���9�\�����wg0S��m�:�J0�	���ߓ�;��IOOmR���)�9C�;�.s����	��fw�FX��y��t�t5Xmnv�;��l�6��IlN��C�-���<�_�¯�G��C�>��h]��l;��F�I�gzl
��_Ƶ��E_Ý�����������1E���Q���*���	F��c�g�y�	Vw�<o�f��	$H�Q)�V�-Y�Y��]�^�V��|����ݮ�k�ve�렓%�r:�DRLE0@ I� �30�������W�ׯ�t7�̼������W�WAʹ��{'��=t��[ct	��_;BGO��S�/HۧoYZ���%����]��4Ġ7e��ҿ�~��~K�P�������S���=�e�F��/c�YO�ʢ���~={���2N!�N�xc�*��e�ʽj�q�p�x��裇��^�q�6�%�6���o�L�_��Ν�Z�]��)�?�ܴ���s���l�5ф�d m���J����z�[ށ �X�I/|��>JaG �[*|vo��/?!��iFJ_y��t�����j�] ܰM�����Ѻ5k�ǿ+ �e����{��1p�e��_~F�kQE�+�6����aڰf#�X9�z�}��O��9q߽��F��&�N��媐T6��;�!��^1C��5TA"!�j�<��c҄��Q�~�,y
M�c��3H�3ct�T����\��Ϩ�_;Ɗ��Nb~ݶv���ĉc��JvE_?�cܐ�#Q\��*��_èÓ@��Ěsҫѫ�NсSG�t��}E�4C	9�*L`���jc�&����Թ����L�#	]�'nI%Ӥ
�y~�"]z}�6f�鮍7���!��2r�6���U�i���`]���r�؝9·�ڞ��"���K�y���mH7&�l�n�(�dzg���E��d�!@���\)T�c,k�2�8��;�Q�� {����b�o�},����C�I%�*�q�䔬0��Λ5+�ݷ�[w�A�Wo�G��-,,��m.���?�h���N@,ܑkg�n��ڂ���ۺ^�{J��J�6v�����7�=�)��0 et��:����{���"={�E����-+�%Q�HNz�FVK�|A��K aI�^ɾ�;i��G��0}ca3�t�o����.�2�_!sVN�*�gg������RfȄZ�J��<3O7o�E#�.�[������:��B����PMӔY_��b��Wtt�'>�+��'��b���u�biI�Gm&e˝�D\]��p�#0J��\�����%�u�pMN���Ԭv��
���v����=��D�,;q�J���sD�ĸ�:u�=�{ �T16#�7o���.¼៺�mB����_Q�#�
u��ǔ�vO��zڨ���^x�U=r@�U��X���;NH1�;�+��};}��E��S�_�ox�fjsl�RF���ܼ�>�s�b�S�}��G����7p���ǋ+�e؊A��⪐�W$��i+P�^��c����U�s�N�~�Fʔk4��A� ��[�貹�w/�"�1����uNO�Ӌ#����+�2Uxu�[�Ε��t|}|��*��]6ݩS+�l�яb7�'�����Q/���Y�$vB�B}�^}y�n[��n]������/NQ7��m� `OJ�<{<���4]�6J�g���e)*���<�4~�N^��ya���e�T���ls2#%V�:��9�*'�f�[�_�w[r���N���]�%&HV�h�l�'p���*�:^,���}�{���c�ܱ�?����7�R� �����(�}�]�×_�o=�ki��im\@�4��j���������E���fB�Jl�r�"jK�-7�#?�!���Y����d�<�P*-��c��}��)��O��2
�x�]�j�������Y�E�k��%Uͥ
�Xɲ��VVv�N��>9;Ac�R#��+�802�Y�,�dZ�3)g�g�k/>B�|�Ct��7�٧���חF���0���(�ţ�N�@�2���(�az�;�C������7tiq\&�!�i��S���R�U���+��`w/06	 �?���]����^�&J��ɋctmbR�[��m^�����L����]ȑ쒈��hI~�U�� �x����2�T!J���.�x�=���Q[GA�Ȏ��б�'i�ֽB���2��oP��E"� �lE���KJ9YIm߲���@`����ԗ�d��2��J�zyr5�2]��>@�{+=��F����|+�r���R}�#�Øo��ʍ�P�\>M�~h�����#ߧ�����ik�J�gr�/Ui��w|~\'Z��7�V��U��l�F��5������,�ח<`,
�+�G�<k4F!�ܴ���;V�!����W�
JkB^\ M���F.MXЏa1�����4h!]�Y�Fc�蕉˴�w�Z��6�;y���O�;Q���❺t�&������H/\�+����5YLר�.���9j��#V����X�B<�!+KJ�=9�̺��<�i��!�Z�\8_:�����eԸR�$�i���%H�-<i(!ֈ�b��Bh���P�2���6��D�.cp�M��&v���J-9��N>x�Wm��|����o����2�������~o>��L<j]|�O � ��&ck���n����o/+���b�A�wN�̛cC���b.K��~'|�(=z�����{��I���B.d�.$
م>�g��	w���:~Df9�X&i��Bsa?��w�'����Y�d��f�h6:��Ƈ޶�<�t�q@7��^��$�� �Rހb>MY���~�[�`�����g` d<�&uRd�s"2��GZD�?��@�n3����>V��Y��}�E��jҲ�+��������~�?ӡC/Ӧ�=�X����^��qyZC�-���R�|,����� {
��&���<�����?B����C�/��]��O��5y	����=�&�Z�h�'��װ	
�0���>�VҶ�U4\� /o�ۼ��2 ,����������)�h)ey�e��!�J�1�6[�mC
Ȣ��U��d�޳<�1�(����$]<�H+���5�NZ�(���B���!���4_^�k�t��<]f�[b�[´�	�Y#Ӕ�P�Y��葖�걷�j�->Y��DZ���5#Y{�z�h�Ә�J�wi�JH��TKSȂ^Gf7��[��g���ޠ5�vZQ�>vW�h��|c�<�^�B#%ZD��+�(�f��V�g��#	z�H��u�wd�)h�k9r]7r�U" �#�M��<�F��{�V�@X��(���"��^�J''$-{�}�(I2�][�Bܤ��B��(t�=��!��[h��z�w61�:E�9����(���#�|�f�]����Ƭ�j�,��0պ_߳鮞/��$"jh�������+h� +F�����h��aڽk�^�Q����0�e�Fz������k��Eʭ��'M�=m@�Do� ��dY�L����,��*��ZX�:�Y���|�6n�D����&s�a��h� Ґ���&ׇ�g��V�@�fY�z����K~���������,mX�N��;�?�/��>�W���x�ں
,�R ���1�A~�2g��( �:�����ӧ�������4��ïe�oG�\K�#���L���"���v@�X��4�j�Pc�������w�/��)N�^�eT�o~�7����ҡ�YѲ�,�����,������]��s=Q�� �j�i�J�m��dH"��(c�\(�9e$�vx�~�_���ct��̳��a���LF����� �/-�_}���u�E6��Z�\�^0���PٺЈ�i=Mj�6hCF��\����1�p�=���{0?.秅3"@��d����Ժ�k�)��!��EJ%e���Ы�	ܰ 'Jh/��ܙW��\���,(����RM­����Q�JTÀ8F>|��D��5�1���@��f!��k���	�`V�>��@���hk�{];�����ݟv/K$%�fou7j�<VkoP�,.�	E�i�����a�Y���]r-M$��ߎ#�]��ZZ�c�Q��K��w���c�e7��[��)�ۉ��#Ǉ��3tﭷ����4��Z!�qtatJV�e��K,�$ ]/�G11����$���}�o���_=O�6l�5k�So^��6v����+���0z����Iŭ%!cT!JG[�J��@��k��u�����K�p� ��ha~�^|�yZ��'F^���9���dZ�(,cia��>��"$τ��,K=�6z���hך-��wHbq��p�N6"����Ԩ�;�Y۶z���[��������3�/���d8����F�b북Э�X�g��蠛v�G� #p��$�ob3����׳��@)yZKe�l7P6�c`H+ ���T/U(���Qi���,ý�����'��_����+t��;hu�0e��I	�ذ�Ő��c������ O'�¨�hU�Y��b�m6���y�sę���2�lߺ���c��*2���eg:���L7\�
e�F�.�L�E�<�
�w�q� ����`|N��){��c@�$
�c��,G���L�H<�]oފ�eW}m�p�۸����N�:��ƅÞ&��:+}�̕������T��&#�Z�Q���P��Q<~B&3D:�B(�p����d*m(�/�h��ݨD�X�z�14��&u>{K�&�1hL���-HBѺ�IA�YӸ��NZt����N�^����D��2��7Q���*��o�]����Oѝ�n�w��A�g��2%.0@���������o��mbf�ʌ(�P���D�I�)�Λ��`���k�A�����h'�b� ��_:|X��޸�FF&9ڽe�ڸ��9v�E$\��A:AW��}��s���N�9E�~�Đ�y�o��:�󴆕����$�l1G�RM!���0`1Ӵ�o*�0�*\��*%�d)�Tw:K��s�H?u�OQ��KV���?�^E�W��*��yĠ��im�ݽw??s�*�T2��9F;k�p��1"M�̗c4�U,���g�+�A{n�)�g(�G��/��Ghӆ���jJ'��1~�*R-1G.��Eó2��:�K��c�-��=Vf�Scd�֦gr�������j,�mE�H \X��_�{s��k6�9�5� 	fP9��������f+����+#���
.}�K��������syofg�7�u
���r��"kj�`�I�g5ɬ'r�Im������<���؂擯WC�<�ؠU:�N�D?��h����P�8p0�J��D&WN��ۗ"l_�a�[�dm�$���YAq��o~���_�l퐀�萁������^�/�h�k��oq��֥%Έ�X�
ָ�bh$��j������%���,��6;�V�q&$������!�(�	���;Oԩ��	Q+�5���&?W{���h>y�7�BxSڸ��j[(�����+��s��D�;����غ��2ՠYW����p);�zɤ��M�-K-'#A}z�<mA:u�4-���EVm�۟�MZX���kWI|1yԥ.-.��L�j���^N�_�u��A|�N2����pj�Ɨ�,�^=> ��>I#׮��N���;�����6k(����8]��Fs��\��:AҺ؈Q��g5lt����C�-����U+�(�^/-5�u�v`���!P��!��c$�P�0��$n�T�j�j#��g�Έ�\h��J�cgN�2���6A�C�=�⮻��r(�m�-�`�q���\�s|�����Hs�뚒�L#�%�a�K����+/�W��5��_�5ڲv��C�P�(�#p佼�s��/��"ޙ1`	�h�����R6[���.��w�MF���-��s����xV��;��zo޷I���鰃�h ��F�ȵ��Y	T��%M�����J��Ɉ���
����ʫ~h�y	^g�զ�ֺ*(������f��r�؛>����F����(�	$DZa�$K�D1
�?���"� ��#�&6��3����R0��d�:�@=Ĉ�fv�)0�M�um��H��z�	eQ�P��zR�(��$�aD�⯾sY͵�°@�^���%��%��	����
mcEkS\]!�����d}a�B�')W�%��
ֺ=-��/|���<E?�S�aᾟ��b�j���\���'�Z^$����N92��b�p�`�QفQ%��\���ij��"+zzhhE�`cZ�=�e���u�]��i|fJ( ���%]��ӄ�)z�	��.�_������#��$�~�
��\��JIh9��?��
WZ���B������ZF�?{��=^�L{6�,h�Rf�^�W�-И��I��@��R=hҋ/dW�l�A��Wӕ�Q�!�)[K�`�3�������s���רoeY���&�u$�+��ӁM����k|��(+�%A�H<W���/�BC 1ho��l��� �1@̝e��W����ѯ��ݹq�z.�6�#/���ϟ��Wβ|U5A�@M|�=��n�r�b�D`'
��sdy��y��¤�������� ژ����<�(�%S��`�AjS���'@� R D))�� ��&��m��^�( c�J���Y%�g~�MI��X�d�ܟ��V3�,.I|�B�`V�[Ôm�R��P�$��#&%�����b] A�(Ϛ��+��*M%�Фp�-�F��nW�)��dE�2b�����XK:��0�I�	��I�����ގu*�H��M�&�+Y�e]=��@��
$�o�!��
��|k�P�ӧ�|g�f�%�ܗ�@�{�Yz�����z+#��,��Ԉ�$�h��Mj-�b(�2��m��T|��_�_z��������F.PJ���ʉ7���E���[X�(�g���Kt��el��YH���d�D0}eC��7�~����i��&ʁ׸\�Ӂ#������:M.̈���riAv�3��q�{Zw��$b�X�Ʌ%���������o��K�o����G���/�ң#�%6��������WDߴi�����w���+��Af�as
ɪ)��������_���;��FY�Q_�y��iz���t���[X�NI�*T�8}�>��K�ӓR9"��-�u�*'9S ����왥9	����:6&0��~���O?E���?H7�Zw��{�~p���w_�
][��z�)=�㌐ZU/�,�%�	W�{~��1���.��y��fW^d��G(�F�j�o�3�	!��l�sK"���)�tԚ.�	W_�I[��n�:ix�윊�R ��DFEJ�����նh�$X��J�Pa�z뱒My~L��m	Uن*p
Ĺ�q"���Ծ!=L�D��hw�W�kn�XS�L���Ӣ�I�>bE�1�V7�ҡ�Xٻ�O��h{�uɰeZ��W�J ���^���}'FS�,ЭI1��c))��4�����%��W��ڑI�u��0B���<�YI���>��H���+�];wK��&F�Գjq�Q�?�k<�(@�r��S�<�+Oz���Q��r������~�%t��������d4�?|�Fg����3�Ҍb%EZ��7|�xf~|������Ӵ{�Z3<Lm����f��z���lL�~�x�;t��1qQO]dtk�5��F�Q#�2��u�VF�3��4?IW>A��Wi��m4��P������B���פ�MU�4yJ{W;�.u��K�tef�񂐮��j�BmOF~��i�t<~�<�ޟ�!��{?H�J��~�,}�;�Ѕ�en����߸��k�z�fY	f��$��-ū2+/\ʤa�a�d���\�{�`C�
�r�$DGG�п����`������9:�h��� �U�h�R	9��?'ʛ oϼv�*�'4�b%={�0�1��1�������!��AnZ�O�s�� ��+͘Q��H=F��oZxR{]}I�1B eL����8*\a�PȜ�����:��z�A��Q#�a� 1~Ơ����$"�B��e\@+�3�Z�g���Rt��M�%lDwݒG��,�<������d=<��U�zPg���b�v29%����m�'��Z��Eär��qJ2���aK�h�G��G���XM���#���R	�j��oh�,6�N�2�^Rp�9���*�2A j����:���eP���/<E_?�>7�1��p!%�p/�w0�C~lM$2(-1)���7ɇ��пq��۾��o�B��3�ұc����X�F:b4{�^��c��	v%(��L05�!j��|Q�����)��뫋3t�����Xt�� ��S����3t��I��w���D*�aá�(�þ�h ����c=�'J�~���:�[����ڎ�;A�tS@��_�qKP��`p#+�s�c������~ߪ&H�,J�B4Ӥ�z�����1�Wf'�~�τ����9�}���B�G�W�`*ȀA<M-�R"֔!�B��WjQm�GF�^kJ3�?>�M��GE���W�f|����45���k�9&���%�D���RK��H�|p���8����q:�*�g�i�D�$A�So��x��%%ţk��@�a�5��Q��t3[��&�!����YmX��b�hB�6=��U�����8�i��YL�saA���V�m�2
]����Y*��Ԯ
��"�F�Ёgb�nJ��*�`!o�������%{/@�:9"r����)��!U�~����_���д���DH��VRʹ��ف����J���mM��z�U �C�-�+��b.m�3T�Mq�ޗo���tJ(@�졨�y�쬎y�kL�>�(r�	�Ơ�k�u�xp��� 
A�LS�V�X3�۬�N���3��~���ёQ��S�"��� 4KYv	ˈ�y5-��(�F�l�t�|�:
� 2Pi��[j��(	����4��5@ВV9�JEC�ex�+��(�q\��q��d(IXوҌjY�����#*�)/�j:թ�:�����vIn1�Ԧ3�M�I1�&�0,��w�]�RXVY@���o@C%�<p�K��&��U���]�I��"u-�/Nq��W��$�?�5�Ǉ!F�Au%r&\�F�+)�1r"�&����HM�M�H�Q�F�Fg��뤲��$�⡧�p�L�F��T�"G���X��v��!W��n��V-d��3m
VR,��T�,���[���@X˕l���	�l8��TVcc��U����&��eT獖�� �r�-	%�0qؠitfqk*�߮�[�bk�+�H���=�N���y.��U�3�0��M�n"��%�"7��U�F�E��W��މJr��{��\�7��Մ[[K��(�>|��2Mג�k�U��wa���^\�'?G�a���g]X�"�;d͞y凴��ۨ}���ъ��EO(���؆����#�D�z=��qȀnR�W��d'��I�!3J�j�2�j'^O�:f��R���s�/-o�2���eg�=!���G�S&�(�b�ڈ�$ݓ����e�rz1A�^�h��'lb����0�&]��^�:�Ռ"�/ݎ�<_'���p&R��\�b�=�$�����-1��kʄce*�=Mp�XɎ��y�,8���K<�F"l��h-TdH6Yn߬)^�W����C��ņA�$E<E�شlK�}\µL�.{O.���c�����L'�z�xQ,�xK\�@J��<;YI��6�Q�Z�/2��v���n&ʂ�w��3�+���*�%'��c���(�_h��O(YE�6�+rB�B"T$Ɗ������$[�C�n�����Jކ�FZƋ�Yy���,��>2EB�Ģ�Zi	p�"%��>M���j)��P����_ƴ6����F�G/�\}���'U�Yf٧,�2Ri�1;2��u�`�P�ϗ"��ܜ�C��PF/�L�}�r"C�r)�$��%F|-�.X�B��4"�(���Q@���+%-�^�U�����;rY�PUHr��I�!6n׉@G���g�*�{��ʱ��GX����\.{Q�±w��6�udF��A+5d1��=Hԭ�g�>ԋl���;%�_�jPqk������"��и�S�
L"�)�&@8%�i�gB�z��Z�W ���
<�ÖE���=u��:����B� �\ߞH6��:/����˴��ȭ�*/<�d������0D�	bld
�)�T�.�t����܎Ǜf���!wG�*&ୟ8���_��~�%�b�"_]q�|+�V����b��_[�)rWq�X}
3��%���(F���o�=�)�)�`pq�H���jn-9,$w�_�z���B�&CY�&�߫�-@�������+��"��;���]��/��7*N�$d���"�+��Kn�0�G�P��� {bh����JZ��U�[m����%�W!I+ue#l�D>q�&M��ۂDˍg21)�c��<%���A�3�%-����()�T���i�x�=3�:�ڸ��߁Ied�˭�{����9o���'q�8�a���Y�Ō��k�_�H�}D��(����6bt���g+Hp
������t{~���Ԓ��B^���3��]�d�m�Q�ڌ/�x&_���{�b��b#��_�d�.~`���`��i| a�4�T]�J/�x���)S 
!��B$�ȍ��E$m��'�o�H�t2�YYD�uhmB���� I��u�:b�bU���ǧ�nO�-V�_��x-�rbBvS^qhF$Ҍ��'
SnmI ��tMn�e[�T�����j	��h1�*zRo=�&�D�p�Z�E������[�is�e���	1�{��e�dB΃q0�2}]��.ҥ�#�
=)qHO=�?��!�V9I�(�TFc��w�!ۜV�k
���8C��A�=8
��Je6u9�`i��_&��v�M%B
e��ˏ�!w =��;�n��o�2$��R�ח߉�F�	G����Y
�˻�z�d:�)}	��6�qL\O��HD�BqS�J]rX�����Q��6LF�V'�<�O1�h:�dɧx�S�?<��@o�3�%�z`qۖ�q�!Ҹ�=�&�")��g��x���H�!�mGI�P��r�g?Eq�B���-��e�|]���$��GKW%�j%۴2/�~��p$�n{���uqP��k4c+�l(��t�45��`��V@g&H��p9�-�wd�cI�.�%HC˩���kj2��&��B��bFz�,$e�З#��a���Ы hi�bd7X���1b�_(�cB�Ho�oO� �A�T� 	G��F6�B� jj��
��ݐ�M�(�C]S�ڼkQH���L���b�.qH�֦, i�{F��	S���	E٨��<���͗�),9�FG���W5��kU�UP_�d�T�uC<�p��^��B��l�C	rm*M �$ա�_\[��/�kW��{y�
�.V$��X��0
k��1�օ��gJu���V㺸jZ�匠VT�) 8��D�9��Ql��I,�b����@��	�>*-�ǳϷG0�*<#�)
\�ҲR��<k���4�� π>����۴i#=���T�3�����\>O��4::&
�$����A&�-�?Lv��s��L��,�د�]\׏T(g�&�bT�%4m�4�jJ��	���A��Ny�[^g�d$7)Z>)ŭ��E��:d��4���D�}d�d����\�UP���iG�0ݰm#��Hh�㰉�F�&9�<, ���Z<���r���0����n�����/I�I�Z�d5���gÒ�j�/Fn��ާ�P8��]5�d�'�Hгa������(R����)�� E����x�����:-�����k�Y����p��@��f�ˌ���º����F��b,��=��T
Y�@� ���P2�v"K<������gb0�TB&&�Nk�lR��f��o+�a�_ ͢�{inA�]��b]М��,����^q�{�ef(#�p��C��ZZ\�}�5�c���@�:����M�����kI���}==�+���S}~�6���7� a/L�=q��{���d�q?D�:�5BO���V�D�Ȩ2RW�����0d�2�h6�W�DB��We$N����t$%��r,��Yl1�D,g�N�@B��B�$�5�R.��9H�R���&%��\G�W�I���b�co�J��PG��
*� �0K�KI�_![���@�TA'�uZt����A��bg�� d=��`IϵL��=�l��-�S,�$I���+I���	Z��fP-ѐ5.b�dz�3�,b&!(��6������q["�p����="�N<W��</�d]�pH<"����F@�q?�߱�7)��,AZ	���8t�����\�RF�����qGU,���@�|5C�'�"s�o�g�\�C���JW*2��.�V	��!�R>���⑶��nH�xhG?O2̼�P�P�s����]�C���s)Q�x��M�cA�,��O�޴f�ɕ�D6�Y�7y�fc�����7�Y|+�'\d�M!^AS���_{O�`.��FP'v���� <��-�&<3��L<S�,�"��)N�(Y�fx�.(�LZ��z�1!��:��ǎ���$͌���۱v��/�2��}X��/PGG'���9s�>�����K���Іn�ob��DUdh�B�Ӯ�n�b?;WPOw�����p����h|�d�)E���Ꮾҡ˷�e�ʵb.2(�A)�Z� ��v���fJ�,dkvj��'&eڭ0^��B�R��U��{����
HR�U*Mͫ��=Bb��J���MF�@aW&hU� �D�2�.���+����g�11���)�*�j�<�"��p~A�@���,m_���o�L��2��_�%��WU6$L�([��1(�Q]���N��Eƣ�b�����*�8D�!&5�~�ȋ��ZJ*Y<�Gf�7"�&ɱ cLF{�Hml�����C+�!E[R�2�I1:(#x)u�X00Kb���X��wBƚ��	63I�Ú��&��"F���Pc��75�$V*p���	[1*m�sSwq���R���bl��?h�K�,�ƌ=�����!G(���3j��Ƥ�b�#�u�O��"I>5-&&��x�����Z����M>��A��g�c	��^7�,�I.����D.
�BRH�c/	m�a���:��#�ոjU(��g慭��� �s�Ѿ�]�5�O�Y��g�H�Ќ�dAM��<����&^ՍnJ�IP�(�Υr�֫�V�*>xH�&V��b����~:}�����u�z�re��ML�'>�I����K�T�+J�FK����Ư�fS�)�A��Vez�(�t����%\��J)+����̎MQ��
M◤�!5�`U��U$�j~+��ߗY�
yy���E�tt����X1/N�Re�$ר�%�T��ȃ��2O�y~�V� Gk�so9�x)i�l�`Js477G��%E�?�����"�c�b��B�^W4�����)��Cu����?@�|��\<���	R���V>/r=	��B��r����>�ķ�D�ƿY��"<������J6���ܦv�(K}F��1�7���X��1����B`�#��$����&}ҍ��C��EQ�c�7�\j������2�ڳج(�P��ሃ�r�j{C�هds�<EU9�K�;��
��@ ���e��C�C��qE��G�3�lA>�?/k>�&� ĩ@$�`��)^��jB����4�#��Ȱ>�;A��Wg���Ίp�}���%����D�5mD�œ��I1�k�+�⮸FY�T�9E�.���'C�-����{ ����$�q�{{����QĒ�L���?jnZk�.1��sqrغ5	�ށp\öF�-�l���[�������k:�әcV�X-m�����]�L��-��KwQ�_���ߡ��k�WD[6o��~���蟾�eQ
��V��r�$i9�.D�^�X��EY���E���ezff�*��Jv�lY���r�oS����<!�X��J�*!$�wvvN�]�tii)���a�ĕD����0�8VH�Jt�Wm�焑���h�4�ըT*I�H\<S�!%�T���[���^g�� �J�*a�Ύv�z�F/_���q\M��=R�⢑ɑc�����@��~��������3JFϳ�]/ުȉJ���&�4kf�\[sY���ڷ�������42;�����Б�2��=�P+����̕�tf�U��d��a�E�c7���-�`{>R��e�Bw;�4�E�~v;����jx�F��/��z�}(��� I4 E��N$!���d�?L�W��Y>��Μ�
_�7=��Mӂ4R6[Ak6*���e����ƛ��ωK�ib~FZ�$3*�֖B��<��w�^�m�d���q�-���%�~�ʫ��#���j*�2"��p{��z:�%>
4�8���0�g�Ev�1Y �[M�4wakZ���W�|/��a�9�
,l�(�MS'������"g��H��:=3M�JՊ�o��ņ6��l��x��D'm��|=�����w�]�|���|�M�&���*+���%�[�kb\9a�O�Z�Ξ�H�������@H�1�s��J��/�=���2ţ�U);���������HY��ZI���@bnjj����E��%~�1܆�i���b]�I�w�W%�2���E|S�HdF�5����FN.�[�}�R2�	4�㴃��dM+��t�"	L�%u���g��u���_�liH�s�<F��n�	�H���Z�H�bt��=��ۄ�9�"˾"����\�̷�~��.a����de�^�t�:�:�?7�u{���b��U��.;F��劬	�tVft��e*e�d��0� �H��a��\�O?�����#g�ҧ��9F�#�]Ń�I��@�]~������b�.���+�t֧��<=t�����CG^�G{�����=�aF0W苏|�Ν8B�6D{��!*�)1��)j�5e�������йK��{�1z�����a��P�U��$UL4�nPU{=���m���YȲ��o<��\�,n\��x8!tH� 	��
j���}�P��j�Y]��E���gh��dٵ�iaz�Z�iOh�2l|
mi�lU3T/{i�*��1���y�@B�!�)�V��Uih��1,��E:
�(!f�n���k�T:WRbp���,�$c���FM%�n��9O�Mܑ$���K�;;izq�EB����)���5���}�+ը6�0�5e����"�=Ny�x�V��ff�$�X�,��_��g���U��,��@���U��U:���F�./�C�A���X[V���LP��;P�J�\Vb�a2!�k�	%k��К/�,T���o K�l|	 hj�;I���6�"^+K��	\���#'6�� w�d{�gE2��7�S����I$��tk������Y~�2���!�$��:�h�������:N�����+aydz�M�����~���gP�d�4��j���&��r�����d#S���q��z�I�=�3W(@ɣ��mʜ�d��߲g�2b=76B�s��q�B����=[wЍ�����s�U��gw��F�;�Hj;�պg�>���}�����/��wʎ/3�i��jZѿ��m-NNS_����RT���?<E�
-U�Ȧ����Ѫ�����#@�\��mٸ�~�c���?�iz��aa�A����ϚH',�)��D�؞�������~��9���~�]�<x�9�z�*MMNҮ=;���z7=w�E��S��jP}�Њ����
-����ۤw�Zo
L���d�
�Lm��!�u�����`�+�[
���o�!��+Ֆ�I6���A����T4g�F��]�5�d�_.����Ң��2iZA<&��{5�*_�\����B,s5F@�Tú'h6m}��lJ���0q2�8�bZc��4Q���P��RBT�@I���vF:e�ReQ�QZ�ť��<�/�-�C�P��	�� @��:�MUH�3�HO��q*�\A�{p({�s�����@�������K2�)eP�/H�t{0H�Z�LLt�I��?�%�R.v�T.\Ʌ��QٰPIU������wwuu�g��o(��U�\�<��\'��O�/ƾ��Q�%F�9MC@P=T��� ֳZ-K�fݚ5R���y��!��]7w	�.b�?���kPp�#z_�)��[��M~�P��'�Uy7��WB-��{���8v��I� Ƒ3P�@�ϳ�
��@˨pp��u�\!
薍�����tvf�����HP�Ms�4]>��Ku�g�nZ�f��w-5�����E:>rF�N��
��v��E�z������AJ�b����,�yjϵ���G�5�^$#n�@�əI�D�,,#\�p����:f!��`:���&�Z�]<s�N��:�;:���(-�g���Z
kډ˷�i�4��׎���s2,�]�i���q/M�NK�pEo�$c�l�)(�+�=N�����C�b�g���fJ3�8r�K�75����A���I�H��(��������q�P����`E�=�b��S�L
���KM-z���4j��d��#>*��p�M)BXh�9/F�/��!J�ح[KzN���8�iO֋�$�(3�Ak%�Tm��.筕k� jAUX��J���P�l���u������]�Ps (���E���W�T>�=����$
W*k��%V�5�H1r��죫���kXI��>{��p4���h6n�Hݘ� %b�<��� �������3�����h��(a|M;�!E�6=��厭����S�x*W����]b� � C׮�g@��$���g2�Z�]�UeA9gBv���g����硣��Z�ҹ���ᗏ�kGߠ��yi��cxN��,K�����!�~zh���-� �t��HN���Y�{Yk�O�J6���3ZA`����~�'�����Ut#Eа4��P����w�TB(�4+,Lx�
b߳-U��AZݳR,��9V��_�����������H���?��ʌX�*+WLA}��O����Y*�����ҵ��TY��; ��y^����G��.�/��Ct����gT�AM�}��[A��}t��U�r�
��!y����h++.&������$_�A{n�Q�~�{���s�3�A�8dT�)�K�A�`5
�*�q`%���@�@m��B� �MS����׊�3�@���3�qW)qRQ��0��H=�L��CU,lP�$����K9�
F)�B˵�i>Z�Fs�*R[�XZdE1��ˈ���j-j��	U��`�Y�3��L�1�yi�,tRg['�g�*�E5>�9�X`ĺ�(dIP�*m$�2���lM+A���t�e��.��r�>`k���P�9	)tS��.XX�p�
$�KK%�g�����EA��|J���(���tG�,{��n�̗
��]��:��$ˆeÆu����;J˺X�֬^KWǮѣ�>�����i�3H���l)(a2H`�`��T$�r:0@�}ǃ�}�.*�A�de���|zv��響D�?�(I�Wm�i�(��M�տ�fˈ���s8��Kw�~mڼ��Bz1�����jz��'����VĘ�V���Gh��z��%�T�Z @b�/��J�U��;
�a�0��iO� ��, @?qL�9��C��q���"�tw�ʕ+���st��ـ���3��J"������,=z���
����"����`���S�W�䌯�]H�!6QF�$����}qךvD�|��'���1b,��i����j��iF���=\�*�Y�����������-�Ⱥ/�*��K閛n�m�����_��G�V*�{_�D�ͬ'٪J�7n튕���a�[����'>l�8ܽ��v����^)���E�IR$�l����[��M����\��k7��{���������䨄e���]��#�F[7naŗ�J�{︓nݳG�BŎn������/�+�����f>4?x�j0�;>Q���3��Y� �<��R�d⥯9,� ����|'��l�!b��W٣(t%���EQ̤�i�4'D��ٖ��~�и��ĹC���Vx��aQ�ˊ������-�R�=���z����5r�*/I#>/��T�#i!�5-) �a$xq�Ps8�p�P:�ʽ����:�ge��9F0H�Ayud���e�����99�Fh�F�-,I�Fdrq�=��N���<躹|�|�@�b6O+zih��Μ9E'��u�6�:V��lN�P��ף�
�(枻���ZR]B��l,S��F,Ӧ趱}���* �!,��o���MFfWzA��)��pmtY��$ה�)�z�?3�G�t�,]�2B��>ڵ{/ߋ�[�C�4��>3jR�p���>��(��Gmʹ-�3�E{������3��HL}x�zj+,���R�m�aD�L8��N�#۶m�[o��C�/�֍8o��mķ����	h#�_m�+�8a�%sv�&���+�%�GS_�r�2Ȧ�ti	��dLqZܸ������yC�k(�揘����j�2v����c4��Rb��7�8U���'��X�ɩ@C���]�@���/�Co}��s�.�*��@�s�~�zZ�q�%�R.�o=��w���t���t��yAyvIR�2Q \������v��DL�����Cb}�r��z�^�e���Ї�i*�"Aa�'Sa�/)_`e'
+%ɊJ�L���vVJM�W�xh���kSVz�u��{��B]n\��A̲!B��;ug�i����}�v�A=�bY���a)�G�qٮ�N9��ᬏ^�+Z���[Cjv�Z	��sB�~�6(Z��,+�T����M붳��*���k�� eQ0��+� �|�ϓ�{��g������օ��?&ٛ,4(X ـ10u��]=Td��I�U66��::�exn�u�cř��[hα��d������'0yee)ڔ6Oı�:��ћ�G�.�C{��Ì��ep$���y�#��HIg[�,�m��������5\�c4Ti��Ƣ��cŊ4Z+�+WӾ[����/���F��h�T�B�è��Z�E݅���3�Kp��4�P�[�n��6JXb۶͔����cc�)Έ�������xi�8E�(��K1)��+0F����B��	�:�h�?����N�9'���u�ʡڸe3�|�(F5"��n-��	=��G��d�����n�nȩ�	ѭp���ɚ�%��;GN�&��/$������~��ʭD�C����E&ʓ�й������T�3��G2FU|�u}4ؾ�s�t��}����!,p�x�v߰K6;ǖbz�.]�H�@g�d�:��}w�6v�^c����y��0ɇ,�ʠH���ܸG�U��η����zz{e���w1�M�s�^�V΍k�Q�X���Iz�����ht�Ʈ�JI�葬B�K0:z����������s����H�S5����r��-�vӽ��U����+W���E5z��hߦhM�0sE�!Fna�,�����Q!��M��|��5����+�`�$:�4��d��|�r��|��D�j��eiYp �B����C�L_��*���"Ji*BآY��V�����n�ca�1��W�Y��k�7�o$8�]��;��gŝ��ncd�{��40����(�^���iAM��<���1f�tSb���dI`�5Y�$�TW����ƶ�=��7�B�cT�MgΝ���I��J� �n��K�\0Z�Sz�A�ꍡ���E6�i����)0K�i�\ 	=����w�x���c�c��܋�D��h�P[�!�0��=�c�6�T��G��\�H4�A��5\�n#=�wЩ'ip�0�^G����C^���2*��c�A�W*����:4�k��v:[���{�n�e���_{��]����wӉ�ߠ��9�,�)p�2�'c���$c��:P/�����lg������?Hӓ�ȧ�l������ec
H��Q^\�E�$�ڡF;���^����ƹ*� ed�k����һ�K
T�j��5�8�����z���֙�B!���-F�L�$ϼB��Z1����-7���W����I�b��ʚ�az�;�F{7n�Lu���3�@m��ڴc�L�2C��M7��vH����Aн�.��w�U�ȵ+t�}�R/#/��t��4�ɂ�g��M�L��|���M"(�Y*슭^1(�pt�*}�K_����Z���J:m�ő�ͺ�dNC�>�u�H���Y���b�P�Ic�^&�S�����_����ZO���&V��]��=��ĉ��q� ���oY�f�FJ�h�Ua���@������;�@�|
��і&�������7NPOw/��u*JS@M�����Y]�x��o�@w�yy/��3KҜ�%ܧ�1�D�[��,{���C7�t;]�0&q?d�ڂ�G�C��@Ə[,q`$M�
�Tg�B�4����܄O��!i�^�r��}/˨���Y�hx�J���9MƦ��l�5.�������9v1Y�c��Q@�~��"�x&j��}G�	Q����K�#�QF��.]��a_\���qV�Z+��:�Zo��N&�z��0�H�%9��}�粒�y:w��`��u���V�g��\�jM}�pAs�P��+����G'O����+�y�� �����{��6&��^��R9Fd��֑��gH^ˡk�5������I%eZ��._�̊�j�Y�{ۭԱb� V$8����h��8<LT�ke�~��lB������&LC�ջ!��ODB�s�#U���tkً�+p�%�O�Z��%�ب��%�B��!e�"�a!])���ѣ��y&�NeVNSS����� ���|N�b:���=��'��%�D���2z�z:{Ey��8�Px�rh��ؿ�^;v�k^�yxh�XSl�4������G���w��.���s��.H����u��� ���?�퀘����-[���+ƔTMDWr�C�f�umf\�Y������V����vq�I\�����+"�87�q�qj �^����Ȳ�PH�~����>�aA#X-Ui��mt���h`� mۺ��\�L3�3�Mj����!�}��A���i��@���	���J��-͠8����}w2�������%jgc�Ni)��⒒�kR�.m[!Gs�����۰�d3�Ș�1gK+0�y��jʱ�ݰ~�^����e��JVBu�u�PJ��_����N�?>?C�|J2�PySId��qW��HdK�|Q�{��%��0��U���}��4�T�2t��3i%�A�G�Ѣ9�G���EO�W�,�K���}���Q�&B2>5K+�n������H|\4����Z.씇�X�G��gX�_��(�� ����[��9M�I�/Fy:�Ht����YvM�rN���Xy<P�����0�D\���+�G�Ǵ�k�ͤ����[���S�$$��^뺵���ٳ��$>�`|�Q�Ȁ^�4�z�ҡԥ�~��kE��T�3�����U��~�0�I%����T��~Zk�,��u�a������QĈ���'_��l�R�4�ZK���ibb��z�IFx��{�b�}��oѓ�>EC����q7�_���\�FϿ|�Ό���ӣtv�mZG���C{w�(�1�l����w�;��Ni9պψ��N-Z7�ڼi3�ټI�	mZ��Q��t�[�@�]Fn�B������q��)�]S�D�q���dU��6��$V07o���x�=�d�:u�5��F�z��I�ڋ.�I�q3�#e�' 锶dH�,�1nu�ٶy'�H:�:�K��j_�LM
�Y(ω�g{�b��v�1ft8�0/��☞Yl� iGI�ĳ�t��oc�� <�({Tbc#�T�h�l�����+�SJ�a߾�S��Ǥd���*��w��b��W���iFSq��F��\���P��G�-�����S�"�3��6BpS����J�q8J�	�*��m����]�x)��x�����פ.8F@�
�r����J#��ZI�6G�ixZ�������<F�7s����]���ZiG@�,�Jv��gi��I8�@��
�������''�^��#��G�x�e�-���M3���n�iF���qn���Mi���Ƒ���_�EF�#�Fs��]clH^?y��g #��ޗ�{@π?��{$>o��V+�(��N�eJӶ��hɕv%T��,��ŗx(�t��� �;3~�^��]�5�6� |]:��-��WʡR~��̚��*4�h����@�I��u�#I��z���G�����볇��޹}m߼����U�XN�%}��y���ct��qF>s�u#+��n�tYF�e��骺&YV^���m�[��������x�}t��	~}=n��=����OI��.v�ׯ[/��ݗ�җ����o����z�L#�77��?�Q.���mUlWA�|��
�G�5uH�/O��%~���r���1��������h��*g�r,�Y��6l��n����I�Z9D��t����2i�z��ieq���S��**��Ŷ)��LX"#wnɥŕ�ǃ}��&��������������
uw�y+#���������MC�F�����"�/��~.�@�{��&������2}m�:���/ʤU)�j���%Y?�R�&]LQ��o^��؋,{H�6M�&���Xc��!��t�	YF�$�C�gF'�P!�8w��F�׺��?'��@�3�p��6�[ʷ�_/�XյDL]����D�!�����R8��C��@z`�M7���)R�t���< ����kTp�_�#�(vժU�|%Z�n�(���I�<�%�y���g�1�3#�G�<�RGq����<$={���A�)t����r&�Ktu]c�T�T&�z��B��Z��uww�ɖ-���uh��n4-�d�@��}���8$@-��&�~�9^;+�x^�=.Q�7��	�� Z�CuYŝ��2$Yv�}r,H��.j��zعe�q�)�B�V���(F�Sݾa#����i��Z���i��(��wi�[�M�j�{�H����t��X)����d�+=u�$�6�Y/�����=���+� ��s����6��0b�%7���ei!$���ZY6$-:cu��6/ Ȏ�ڡ��~�z%��-=s�J֭[�®�K�Xp�!>�N��gea���e�JWT��⺶8]5Yb�XCt %�HF�K��V���/-B��PUif�-<�������yM����!�����Aj�i���u��	�)�f�i^�-�:���y���3P�-7�Ȯ�4��^��+r"��{έ֮��P��p��qC���$�P�����f����U+��\�F(�fV��T�9�ٓ�k��"���:*�+R�	�X���Q�3[�)����7��<����.�Š(^��D�_Gg�V�����pq�r@�� er��F1kj?q?0�7 �<��:�����`��#%��!.�7�kB�a�w3QK./X)Q�%��*�l�l���b��c�ע�ó�2U;%+�2�H;�7f��`m���h�e��`4���R�z����	�:&kh�$l��L�e���C�F)>'NY.Ӗ��r��<�K���}���_V�T�[/�/�%5��\?�V�^�T��dk�xd��#Dq0�:+�|�S;����������#i�S������s��-ed�s������� �D�������g�+S��&|�7[�� �̧�����+_����ӎ��Y��%v�+�լx׭Y'(���z����t}I'�*��v�D���+�x��>�P�1"3�Y W�YC���>��\cŔ�τb�b�Z��~���r�سtߝ�Rg��p"�n���k��w��|�߿?�aik�q�6u�z���l�+s�4�8#n�� �@:�Z��K��h�d�6�/�j��1�
��ꤳ�O�!Y�r4,d����GYW+�S��h`�z��g��[�GD��WK�B�	֌�R0%�;�������uvt�K�!"!����VR�~X�� 0:��A���*�Zdr
4���(��A.���݌SgG�	1�ڇ�~���"P��|T`/�-Sr7�ċY�--��:��;�)��vV�m�LaP�@��P���L�NQ�3M�֮c�pR�8D@�0`�gg�]+�,�,\Qڏ�o$	��_��x�C�y7��Ƙ�Pgg���ڠ�  �.�׃��5�O�to�J�w��If5ߌ�J�(h2����鬆�7�4�b��gQE�J?���R�A�Hs�k�c'�o��m� ��\A�qo!^g��ڵqA�)/#M*Pl~]kۨ��sr=!�A�5�&����B
��i)Mj�]�'%�ӳ3ˋ�+Y�'���bႋ�S(��)]:H�s]��ѩ�atӖ�3+Ѡ�E?}�h��m�T������_|��آwv�k���`O?}�g?B[7n�����÷�N���4�(Q�5h��镨������a��[��`S�y�)������w짅�����~s�t��̭��FjLafSZ*�ĝ�5f\4�T*Ǯ=8S��7�7�Ͽ�yz��giú���~V���}#��8=;�m��	e������jIbPh�DA������Ff&�?���B#S�dIvA�6l��U�I�i��^/�љ�g�T[���k�rr�Va@H�� �)�𚍬 �i��#�Q�G_�&fY��0��F;�|���䙓43;I�C(&�u;]�L�.]��=�h� �q��t{�C{��Ez�T�U�4�s��Al���]�����v��6X֐/��^H�hR����ԡբbJ5�6j1���h?�(Hŭ�u�P��%*���W��% ���1�E����e�,9�,���ϕ�U�| @�h���j�H���������k�V��&vC���x.g���`� �@��k����_f�s� ��X��W��|�5�{.Rw@Y��	�����ͤrٽ0�F�prQ�0gkB.`@�n'��P����u
������=�,�g�zap��'���6V+����R��}ȩd.���k��:��3
n$��4L0f��`:��6�Ă}�s����Ŕ��c�?C�c�����f��yp.5��v��4���GC}��m���sg�F��}���xvq�(���)ٲ���e/a�xa����{%���AiN�+�������&�>�B�8]��u�`�Q�� �?���#��(Q��>�i��?��jT����?ȝ�;־9�K������Zf읝u����/�k?��D��E==����~��4'�!�X�rO�������i�/�+W�o��r�i�^���r{���Z[�'�Y��'&e����F��o���t4*x��g�>�yn������*�~F>��g���~zaNN;.�x����K���?�y�vv��/�X�z�)9�����ǎ������{�-���������X�܄����˼�fcJ�3��o� 3�!� `��(�z����e]bOí]y��/䱓ʚ:5D��+qMJW�]V�pN?�%>�����ݸw[n��k�l�n����PK+�md�2��d'��śo�?��}����2�A{���i���LO͒]1��-I}l��16d��cW`���;j�FNJhԃԞ5�Ib}}[^}�u��(8$�-���s����Y�[r��-�4�pu��'����iG�=�]݈[{ۜ�}_:fhGM^+� �%��(Vy�(��U�קgʪN���8��^[��=�PÐ=�:�bt���Ť(ɥ�C4��Ύa���� ��Ľ��G>�x����n߲I/ޢ�9�Ǭk�����1 �m�|����<s@)��}�/�:����t�D�;>S�7f��\��D]�`NN��N����5R$Ō<#�� �7��f�3:\4��2�nNXg���ly�Iihf����#�yo�Es�0qkFt�5k ȭS�;0qO�K@�4�f#~�y(v%<H���Ɔ,*)_^0>��mUO�~^-�cP���|��iT�[����7��_~�k��w_�9}�O<��|�����(��9�4{��e���U���J<� �������q��/|Y���/P�K�|�I9��������eW���Ԍ���0Z<�Hx��kD��D#�6�핋��o��yt���G:DNjZ���>��ћ7nȷ���|_C^z�ġ���/e��Q9s�Lkڳp���t��{z��;w���?��ɟ��,/�p_�{�~ ~�q�X�(VQ,�y=w��A�x��]��)�0��,An�[�#ib�&���ɩ~�p`�"�E�"�;qR�:���dXY��u[�O^~I.jd���AcJҨ���exf.mc��f_��A9�xB���V�g	��A���1&��9#��l˝����ޖtG}��2��!�@��i U���_|E~���D�>Z����ut����9wJ���i�%�Ԫ��yjB0=����z�*���9������U+� q)|R}p1Gj�{����2,"Mf�����m��iۀ1�qDf���{�ZcD^Ү����M�9ůn�וØ���#����r51*���ܑ�*���uody���-|�!s%���g�߃F���f�n��bF90ˈ˖�,4>��	,���x����fA�o�b6���m���L!Ѝ�M�����\>��Ž-0:o���b�69	��j��+�����W!#�.�jČ���n޾�8��ޖ���w��������y������H�j�����=yᕟ��kD��wߔx���k-�z̖��+�����/���8tL uA�vlr�KH�}�#�G�?J������4��M�����2;13)�n]�����dS���ξ���(,�2����KG#�4��-'N�/�֗dcc�3�`���>�i�0xKs�����_��Ώ��w.\�?�������E��tt[#�_E��ޖ�����	��4;3-�����Lit���>%o\�1Дpɂ:�Vݦ�ư�{x�m5�w������3�� �a�51�����FG{�;������~7��//^�W/�.��[���;/L@s�~Q�dA�J,�C�����������������rg8�Y7��~� �ÈD��Zo��.W7o�Sڗ�~�Z
�G�� l���ʢF�C�w$����^�S��ж7��O~B�Ј�;G�� �����c
e^tom���>���h����m�X"��zN7��1"�E�%*�"
3N�=�����+8�[Y�U`t��\�U�KZՕ� ���L��E�:�0@��k6|���X��1 :)�?��<4X�kF:��XmUTFF�11NE���,�Q[V��o�?(o����Ƶ�G{��T�?q,�� A�� �>�i���ڃ�z�8�Mא��/o<�]E�%�o������p^�ܠ?)^Ʌ�����ޕ�W�it��B���%9�FX&FnC���Ʀ���{���'�]������L��x�3r�0��xP#�����+?}��?��<t�,�N,-��<��Ú
�jzPCڃ��_�җ�QN�ɱ���[�{^6ww� zWފ��#�ֹ}�tzMu�eiaQ����4�M������`d1	uqeY^��\��.��[�4�%j� e��򅟽$���w%�h�A;����'[���@3a
]o�m�L��)4���quL�����j## ��h�+�}��:TfzES�7oʇ�?)s����>�����<��	������r�����*���h�����\Y׃�јA`eoؖ[������|����h��Ʈu�hd�xt��X�]����X�ْ-��!���Qe�o�)�[p����=��kwoSUϽ��e�`��cl�)w�3�u�Miv~��uj�v@3B!$����;����!zB�9$&����nU��eB��!j�Yc�>������ ��)#�`d���
��Q0���(��7������+b�2�nm�
M�j5<���`<��Vª��pRo����&~��Il㰫U��5�����"��s¹���9����bi��<�e�q��LR�߽B,%u+��m	�v���?�}�l�hm�?��%�@��:���`��D�E
f_7���Y���&yᵟɛ�ޒ��C�S`G�9�F ����D�k���?��<��g�-M1��O��ܽ�/ȭ{7�|�srr��)�B�aQ�B[JT��~�׾񷲹��)b<`� ��歛��W^�/~�T�M4Wш���^mo�4ܑ��Y�h���An<�:�H�'/���>P���D;����Jf&��X.K-1��wo��?�>����Q:��Fd;VDql�E����i���kt�E$�����;rR#�SjȆr񝷸�65E�v��eM�w8�g�ז��8ڣV�K���z�I��RΖT`�}=��n[��|�|wKN����4�[����F]F6��<�@��Ձ�afQ8u�<C_�h�s�i�v�/�z��62���Nա/�-�-s��1K�"�;벩N�n����N	ƀ��g�#s(y�<��`d��`h��ĝQ�<���RH�?'�4��kl|��%B�Vx����Jڎ�n�P>�mں�v���]�b��I0@{���iԇ���(5v
ƺsj�v5��>�D����o1�{�k��ќ���0:d���,M5������?����c�:��Nj��|q�y��+#+�_��\���1
?�_�
�)Ӈ
�&�	ĥpϡf�0�7	C��a�R��P�r��saf�8*($��������7���+r��-n���=�`m5�L�"��pzn�]�QA ���@c̿�˿�_��U��vW�ݣ=0�������/_�f�����SS��H����bA����o�!��祗vY����`p|{�Q�GG��|�k��P䛝R֨��x�L/����;lnh�1ISC�N�/�\�D�������\�{���P���p/���l�[
Gs
����[a޹Ή����6�ۤ�!���]�f}*�G��i_�����r��M��k@����u�#�mȶF�=u�<5�Xp���CDc1y1�XI.m���4�;�i}��1����h��� J��3x���,%�4�֨/v�K�Ѓx�+��7�g� ��J���^e x�����;�(�/�	��ԫę�V��E�b�fG١��u��i������Ch��v��4�-5��S�@?�v�:;���a0.�(V�7k%����+,u%0��"��X%T߀�nll�����{������
F�zb�`�0�Y
Xx�p7;?����v�K#��nĴ��Y$?��s��^�K@��܍�A��P�y
�i��N,�.]��~&+"�P3���%�=�B��x��ь����e�It8����yZb�H���!	��_��o�U]Xo^�@�<�Tu��n\#�3�+��-y�Ƨ�C��h-np�>2�(�AD�=C179-��{���_"}o���Q�>�ۧ��`�G�I���S�~�]����^����XT�^���Q����Ct�bA8+[[m��˨��oٰ94gd9!��.�-5 {zN8�Cg�����2��F�~6���C]����8����F��S�O���۱	y���d��G�n�
^���H��Y���Gy�d��"5�]�ޒW~���w�2�<�b�$*�8x򦳐�x�Ʀ�g�"(d\e���������e~a�Ɯ@[A��� �-�d��ikQ�Ь���	�=W�tHU�ڍ9\�U����L/ȑ�#�`5�>~�FqscS����\B����HM(��#�H��)7��@�WNR�R�yv�2B8���Q-Dc?_�����f�k``�R�U��q�GgTu@R�z�znݺ#u:��&�ԬS:��&}q�ڵ�\��;G�
La��,8�áUE� �������dFg��2���}�)뀔C�W5z��z��
N����ZBfF�k��hϝ���ڈ��h�^��ӫP��1�͚��M>3���#�f|q�V >6��]c�45lЧ�����1LT2��h���q�B:N���Ԛ
�n��QĞ�:��RnTp%)(��A��A��Ц洊�.4gu5�F@����Q9�	�,=�t��c�7�`q�S舸)�gL@������� uW'_Z�Uss�O��}Cjw�����*�z��������d;lxzO?��<���!��?6'Z&��_V$�e4�
CI����MXڟ��/�@��{:�e=6
����XwO�����3�xn�|�ETSc�.6!0=�ZQ� ukӵT�(���=���¨Pr/���88�}�8���� Ml2-��&x�0bh��ϔΛi��~�/�z��P&��/8�z�?�ey�g/{/��}�ӻ����k�U�����&��aM������M�[7k�J����"qa�J�9Z��n8�Țdp���E��m�0��
�l0s	]d���Kr��r����� ~8$��l��{T����#�e��2[�fK!;0�����nL3/��خ<AN4��'�S��ȑ��r�}�A���Ꭲ�'�V_����?M��W�+�l�SCk8�zq!
Sl�P>�Brad[zfS�	���'Lk�3�i�R{���9:�k$2Do]b�Nyh���:�+�01qȽ�1O}�r��q R�BF�	gDM�	%K�I�� �4�f:���ޔU�$�+�3��b��~^��
��v����։A��7�?�L�����!Ҿ &'���D�Mr��f��`t�+3���n9?ߔy�ϛ�=4W�87��(��S�B�Ѕ�9Y�]��lL����yu�j��]Xa�Pj-���Y�
�P�I5��rlqQ��%y@��ނ����c���ܙ���"�kX#�[a�h��V�|�y��0&+KGx�����	���d� ߈�X��v��ի6�;�bWج�NIY�:��i �3Z�����Mg�3(np �G4&Rd�mm�tj9;���K�_�0�U�I��1L��b'D�A����<��2��A�?�g7�����Ufi�����֊��!à"�^2�� {Ma\'"ϕ��)p��~��s��F9� �����1h��%֔�I'z�y��']�R��qt�m�c��l����F/�Qbûm=�y��Eݞ�/8P)UƨM0V/aؖ6u����3=���t��J$�E�n0� (R����W�\�"������%+��KR�]F�R��CRcda*����y����J7�,��~�43P=�>x��anS۔�����^D��㨦>ar*S���3
�gi�e�q*h8���n-���r�9q�8.�y�g���w�D�*}���^�U��
"x�F>�� v�Ԭ�o:�ዑ��������K0>�}J�3�v�����q3�)��cæ��d��0���i�ϲ��5�jj���2�i7���7��c!�2<KF}x.����>�Q\�E�g�O��xr=F-�}�c�,*���{���B~nqA�=���om2s��4)W�2EE����XQޓbE%�ƑC�� �7Ի��c�NZ�X׸�q��=�bc&	
:���оXL�̟F�S�3�_keA &v9Γ���\���V�����o�k��)�V|�116�b�*���w��N5c$�}�1�$�#�=v\�Jd15+d�.щ���([��wS�/5RtONZ�E��,0WZ`�����=���f��O>!��?�F<W:��I:�'�.���s8�-1ּ,VER��_���.d R�Y�_)��rU��d�^�2�=p�V� �]�&�2�o��'��o�Lk�xV��б�Ad���91�χ��(Ja�	ɈR��a!`�����gs����7�+)9���DE,Ǫ�maa����B:���(/),��[�/�{Û��ϲ3�CO<I	�W_yE._���ˁzq,V.v�)u5�)b#�6ı�����$q�iXX�np QE7K١���2�h���Jr6��A���$|i:��P���A!%�M'�s�+2��s�,8T�9�����@ �W�I�6ǐ1XG"+�e
]�kdjz�)6�Al��^DK8&��iq|=8n����z�1�@���EQ*D��^�x(�ܾs[:�:M�Z�qHk���/���"���&�BB1(]G?y�dQ³���y�h�8���~g���8\7�k�9,�{��ﭮ�������Y��h�?h��W��0CKvl�a-�ߞ���3�w���g ����P`øw8����,�(�>Ϝk�ȡ)|�Oq��N������轳1=�Ԇ`L/1q�	~��h���\�zK�٥�b�@G��"[�g��_�l-.	��Ǵ�X��f����WT��P, �($ȥ�-0�P7���W)��5�I�2��͝�����t�I�u���E��P�YZ��zt��y ����1UJ���K���R�wd_d����^��.��<\&a�ԅW�yU�$�W:�@��V`�s�b���F����{�«\t�(�kpZ7L�����9>ex �I�Y0�5�%X��+K_��%s�b��+���G���=	F��{��"kKkBk��a���Q�&��8�=��Q���;����&D���-��9�iT�.Efӧs��[���F�����γR�9<@?AGT�`�K,*�dsy����+�����X�"!�`�?k��_��p(E���!�=T�= �(9<�]���,�q䟙��&@si��fdG�a�5����5F��F�z���<���2<û���<��-3����S���5u�8p��a�6�(j���� 5�@�b)����Pg@�B��]�
6�v�>� ��� ���wYL!�3�ya_U#�~X�[ח�>��-�> ���Q�}߀\*�����߱�h�ۨ��:�V�2S�
��h�M`���p臇���Q���Az�B6V��i�{N�u-�O�"��`cw����V� �P�P2�f��qj�ׄ�HX���P$;2,l��:��~�7����s�L[A���������
7bE�'ǌ/���E��q�Y��F�Z�r�xq�U"��:�@y��!��8{��>>�Rh%T��ޅ_�f��KpV��8���� ]���/~.i0�I�=�>�1�ynh=�#�.��l�` P�P��իϩ����6�]o�K��D��>�#���������](и��|�I�P�"�ic�����F9����Q �ila�bMΊ-�)������׭l8d��eri1u#r�K}�Rl��k���;�K����Ш�nL�(! ������]#]GA��S������u���/֯/�qp�(�q�/�Ϊ�&4�Af$}�"(��|��[a��n��۔YQ|��?/e4k]��,w�SV��fF4�F���?J�@C��HOV��Do�q�ho��U���~@��P����`�Gji���i���*xFXlY�Z�YP��h��c�\@>� ����b*<(��G@eA4w�y^;��BQ�vg�_`�v�c��P���Ƈn��%��Kadb74Z	����Z���a��*X#�n���XЎ�k��NUXd�a�݇�@)��7u@����fg}H�9Unh0ĉF�+ʃ�0�����0�l������g~�+�jl8�\
0{�`>ҩ�����"-�W
�!���>V���#8|#�/��8~��Wׯ��+�SdMA�$K8����H*8��?���]����;��̘�(W�����yU.�\������C���5�Q���DG!�y��,-(L��{=C�R���y�e����2&D�-���٤�����U)��e��!F�`� �����K�6���+�X�%Y�kF�A#T�:L�[���,"�Zg(�Ǘ�=�99}���u�+��{��|����ѹer�Ձ���E4|Ǧ����#�v�x��^Vyx�J,�Y�O����8��c��5�/f�����ǚ[]Y �" u�v��g��>������C�N?�oPɃ��a��&c���1s����qQ�w�})�G�a��_E�WŔ>�Ž���V#�<	Wj!��QT �v�JJOu�e�1e�B������wE�rAD��±�J�z�����zE�Пn�]y�,;<�ᐅ�|f��Ի`�;E�L�3�F�{�\�F/�����k��R0�"�+���{�_��Wx/���M�����~�^Hˣ�7
G"�*,R�)qQ��֗ ��s��eG���N��G�f��5Fiώ�Ʀ� ��u��Ʌ���7`>!���MTM���Ź��������}�:t��HV7�DV��~���3���MK���h�+�iM>������O���j�Fi1��{[����_�l�aY�kZ�G�$�ȧ��Ġ��Q���/c�C���)��NL_]l�J��U�ٗ���Aϊ;�Xq�Ām<g���(G=KumH3p��.,x�|��5ٸ ;�S�x�<}�Ԉ���ۓ���s�N�3-K�����
�m�(�`�����<�.�`i�O0�"�޿�������y��"b�����c�����I�Y
%����}1�y�u�+*�Ai�}N� #�.׹T��ǈ���#�/����?h��U ��4� c� ����9�p�p=v������>�u��7�x���?��+���Q�'Q^w8����_cg#R��j{l�~a����5��Z������`��"7��ퟔ�-=B�4�٠�8b�V㠞����Ϯ�H���C��'܎ʽ(x����Y`\�]ǌ�5�G.�l��e.��+�Dk�k��/^���Y�mY�<���30#Yc��=�^�����cm(�ٌ� *ai�X7+~?����>��c�_�}�mL���˭�-y�ŗ�n�61�?�!����2+���A�Q 6*Ԩ,#�E��KYH�PA�t���.�:�!���7�Zbk~G�^gό��<#��'5��.èXQ�uV}�Ԡ�8��R�
��|��&����n���K�tL��Fr~^(�DN=C���v�&4'ȡ�ң�pm��e�܉�{�ؔ�p?�uƫ���~���%v�ZTГ�a�C�3�x�ϫ�v��x�V<�F�__�Y�S;�z�wf����G��u%���͋�8;�"h1��ᕆ�za,*�zA�����*"��Ǖ��7�.C�f����\�ቑy�-�(>����XDn��(�z16��}���d���B�W�rýF�%Q茲�<��B��H��`l��fՔP�2��>)�E�1fc	�$5ÚJطISE~�a�� �uWش����e'N��^C�6W;X�ׅ?O�Dk��I۝m�|�=�C5:��ȁ��S0. �ד&���'Ɯ��[bQ9�D?���9ε��~���}��Ҍ�����j{mG��\��iY�]��=�Q��ռ=De��XP��ַd����~��t��?D�
6���Ɔ���+b�C�������oiT
(HE�#Da�G����4rSu�v���-&�ʆ����]e =s�T�kSb�>
�[>�D*QZ��[��(�mA�e���JfxVX�_.WRRҒ�q�oߢlaĝefг�������L�.>���;"��b�v+���rhRv]�uR��=Ø3ܫ�T��}ܣA_�Q�:� Q�g�N+؆��d��43/Gg�ّ�s�eV�gJ�(���ܠ�
%A���=#���!�`�b\���+D��2h�e�`ȷ����$�88����Oa37�Q�|x�Bfъʄ���%��GΣs���b����f�k��Cv����0Q+h�]B7#���G膀#�
c���	aB��Z�BC�fC�&�k�L�`'�F&��۟�P�q�$0'��b�v��ϊC0�Q��n+�,DO��bL3q�n�*��=AЦ0����|�mzH��3ͼG�Sy���{Ɇ�!E!�C�|�6/�c?���!�L�SKX��ɋ?����r����:��VWWess��$C��7ސ�'1�o�}�-��/���7����^KǕJZq��<����7%�"�Q�2��Hģ�������Y�d%�	�lH{�k�V��O�E��)3��I�0nF("O�a�����p�8|ߋ9�Y��|��x�x�)�H�f�e)$���oݾM�0��0׭�V`�����E�7�ua���\�1J,�a�&�"�6����klۅӡa�I�7	�_�!�
W�`�[�y1���4��݂u3&Q�h���>�-6��� ��!�ϩ��Թ�s/���.��ch�	�zT�E��y��ƚS�� �R��b3�pn�g,��C���(�N@�Qd��'-0���c����>�a4g{�`���˽�-�X���MY'ր㈍1xp�l�l��6���V*^����w6edĊ�#�I�����
q-����޲'в̕��t�]+	Ye�"�׽n�S\��f�W���t3� ��P���ۘ3����'���zë�y�	��Ȼ�r
�r����k�Z��,@+$T��Ŷ���������{T���F�@"�W�pL&�^�|�pպ��wl<D�0ܯ�����:M��0&t�=z��i4s�!��i݆�~��	���c�����3�2�FDBt�i��&�e�_�z���'�4̋<�|���"�3cj�f�&e�_O}���{�Ř�~�ǹe��˧N��̜\�r���K'����������ʓO����U��7Ǭ1F*?M����h��::}ꔬ��q������/_}�z^�gayY�t��ؐ:t����{�R|p�p�(8�>���ѣ�l�����f3���.��/ǧƍ��� l��vf~��f_���އ��D���(�-��ܪ�� ��Y`Mmjo�)�z=8� ��g!�y�U�d�nJfC���.�ދ1�p���e�����H����_�/pW������1�7�$Χ�BH�xo��]�?�qO�>-Sz�߸Ό2n�E��0�(;(]l�=��gն��q����G���6\{id�$�9�&^�C���z�������1"15���x��`�7r'��h��e5��0�l�SD޹ukJ�Z�'V��"v�"k�Eu:�>�ɧr�9లx)c��ӏ<.��?���>z�7���#�j���y�v�F�ZP��Ȏ�O��E���h��Ѣ�E�7pumU����˽�w���1�͂�t�:"�+�� Z%��с���E�	��[N�l5� ���A�!�8�L5'd02�cE�+V6D���n������%��e0��Ji��p�@T�(�}��Rl�/�V����ԛ��3�kM��Y�K�&��e���۷�G,���o���5F�h��\�T#��/��w�~�Ϣ��Ae*��s�-��x<������pc����;�dwkWV��x	�w�dws�	9�ܫ��� y䚫z=��^o�Rڀ�O�4L5��j ��ta1+Nn��pi�-���@�6u� Fg"�� ��c�|\ڕ�e�����}����C����y#�O�U7M��<���D��;�Z������ys�Vl���N����.�[��~
�f@h�ث���S��!�-��:.p_�������4�C��[4��k�5���K݆&FK�8"��?�h�X
ʧu�R�F\#;!��E[��έ���,+tw��YBC�Sf�>� 	��)9A�юOP
F�~�[��桺MA�����1գѨ1�^���dlrB&������v[>}���{B>�̳�y�x�P��%�H�b�4k�⫤��̋��"���M�f�K$��i�ڌ����bFPj)jU���60��~�/� 0	k�WJ�T���\D-
� th�jiŞ�o[-^vU^.��m/]����Òu.��!�U݀ [��Z�'q�~��Iy�̃��O^�FL'��܋T�s6c�i� G
�2�Xe�G�Ko���u��ZD#��ܙ��ǔ\8N��w��e[6$�~f�
k!��;��׶FM���b�țY�VW�k&L ㋬ѬFs+A�֨�)DC+��(��Z��-΁]xA`�שa�9I���%�^�ӈ����x.l��x`Q`�q촰��0`h��b�`X��a-��o�܋x0�Y(�lvK�i��.h�ah�a���ʵ�*|���(�bPU��Ygɠ<O;��u=u���4~X-����o8��y���N���9��PH��Eu�Q��"|���·���=�C�$���Q	���HL<a�0B�8W>��A{o�dL����P�f��l��~?�K�/�Ï<"��K���Y�Ih<Ѱp����w���\x�$AF/PB�(,��}�xE.����{���t{�_��7orq C�&�9��)p�A�@㢯P����e��ך�MS��8�1�b���e�1,y�5s����]�I��Pڋ�a�J%@?��O38v�!�?�z
��C���x����Ao��S]e�H�%��WF���Z{d���P��uDqnD���U�^inϡ歙��(z��þoD�T�%����:��m��[I�.��A�46�h������	[�5�d���Ho3j��2I?o�f1�#�q����4N�����TW�]U)�Š�Q�R<���giɇ.��,;���x���Wp�YFq|�e�l���70Y�r�ǜ{i�B�ru���X�YD0j�#M]H��J�9�[`�Q�Q-/拱����zd���P ,T�l��<���ז���D�����`0��1�a�Dds�v�jX�"6M���`x���f/-�lmL�f��ڽ#��o���/�cKg��1�H�a�����K���^�[�-���^oW��i�j�-BOx��7�f�H��()��fR��o��?~A�����ߩD�� ёD�nH�������Cou0)d�2h�s���FHӚ
ﰝ�"㩦:pa�k^��7���U1�a	���*+�G����L�>^�G�#�_o8�I
�1�����B�4:��l��a�}b$ys|�p)�"$R�a�FgA)AM'[����ҭf=+6�\_?�y���dA�����L���c���Ş~`{��]���� O��"56����o�?\ލ �)�[�F�16���s�-*�z�e����B�,
 U�T0f������)`��e�G�.7�j�C�bL���ҧ��&q\�ɡ5�М���+�H�*�]���[�p�⚤����5��q�(8�ܘ'��;MK��K�[A?Dڑ_w)�Y��AA(��I�%\vZ�����A�ದ�
�lh�	I��0��{�C�c�O0�����*{�g6�J<[����3�<V�V1�y�:㬦���\�qC>��G���	���&7��Ȼ����ͻ�O&rewU����L�'ec�+���QWDy�C�6�P  ܬܼ8+��1��y�=5�=�3����|)[amS�>l��6�*������p��H:�233ł�ED��DŐ�8iT�~���U��)*�%��"�4@qA��R�C�l���0����>Ҋ4��z})���V!���zmI�'��ѣ25>.W.]fJ̑71���ᆞYT7}dY>����K/�Lu�:�A�i��࠭�uV�[5��Pu�����	����3��v���~>����O����Sg��V���C9�ѱi��\��Lѳ��埙�t�	��m���m��4�4��F�Z��!���� 8��Bd���r�[�FQ��a5(��4�t�+K��H��*T�ȇu�����s&8<^`~8888A��ݓ���sA�+z�Ñ�B-+u�D@-6-e�Q��&��(@���$9��=v���빍y�o����7
qƝI@l��}ג���V�Ė�lݰ���8���P5�<����Y�~���ٰ��S r�~N9�)�٩i�.�����3�_�찠���{'X/�PJ �{K33>8<T��:���9^�*��ؐ(�l���(�c����ު�}��d2mH�?��U?��0Q�^�gt����e�7*��ڐ����Hƣ�<���dzb�}�wnޑK��� ��{��
*���B��ߣ���#��C�=�4�4#b@����-5.*+�a�AXƵ
��>��� 1gj(9��Ϣ�u_�zȖ�c�m��e3d2���2B�o�=�H�c���xSOa�3�ei�\0�H�4��;�C/��6�
U�`d��b�2�L�ei�.[8 �4dj #r��;�r���r�ز�9V�^g_9?F%�Y#� � ��,@d{�zcj�Zs3r|qV���l�b�j�Tr�S (�����{��)�U����*���������bv�u&h�{�뢱`GN,�ʉ��6��H`������$r.n.ͱX�.L���=5�=�ޱ�fa��Swވ����Y��`#�F\9~�F�Q�,���LOس���rL�-uZo��6��`hC����skg[?�_h�بg1ը��sgd~qA�76%廙M�@�l���>����_�/�L޻rK�Ő������EiL*��u�}D������G�= �� #�I  ��IDAT���%�"��B�FQ߇}D���țo�%k�9��(d�F����k���=�:�Wa\[�+Y��t�8&���ڢ'?�Q�}z��%�i[A	�mVL�{��Ls�·��؋�š>3����LW�����敦�#��w�nh��CF��U
Wř��JGj�>�`nfN~~�5y��u��h=�a کL�B�,�r@9NzR���/����D����_����^�4
���B~LDX����F�ߪw8)x�86y�~>�g�3 
6fM������%�XƈX?�toM&��_�d�e�}�������o�Qs�G��C�gt����6��~�{�_Ӹ�f��Ӫ���e��.�唨���)j��˱���ı����s
l�"�HM�
P}�����g���v���2;=���q��Yw�^�:Ad,���[��ͳ��(Cܰ$f] �F��%�f���L�ƚ�T��e�(��t ��P�&؝ǖ�j0<r|vZ��	o BE���C}�ǪiJ�ר#��'��FfvCwe��=Bg5_�v�^����(b�G�	�lh�./-ɑ#G( .�����iζu/ܾq����ӣ���*�����88�-�!��TmR��q9�JKs�{f��[C��ӝ�P�037-��:*o���+;`�����k�b�,�1u��r��t�WgY��U���Ϧ��Έ3�~�7gp��u=���ey�S��՛����m�*�rR�ܧy��[��f9ǖda�!�����J�5�(͘N=�5��M�u��?���&�^�,ۛ[h�!���GG9L�bp(;P����k�n�䡓GȄ����{���%�5�$�,��295BK��dZ����^�}u����}�Ɖ�P��.�3�+�_��239�tN�}�{`��}�>��@�%�X7��E��-��9z�(�T���!橱HH�>s�q.��0ؖ|���䡇���}iL@�y��\W=��+��Ν{��w9�**�B�m��Z�|Q�ƍ�w
w�#����_����Đx�E��x��]�.+|'�M��T�&V�!-e����Q(\���y!�h��w={Fn\�)]n��"?���+y��eSK�6�O�@�!�>��s;.�) ���bS��z��y�p�BQ�~��#��{�ޓ��o�Q@�Ɲ�����g\�8�3_�T�1���}�K5�1u�ȣ;���UBr��z����xuL���h#"�{ro}S�{�#ˣ~�Јp�0�̒	F�>��VS�ᬗ��4����%��4j�=/�%��ll��zS�?a��48 �N|��<d����F^�F��/X�D0��Y�:!����֥�i�����3�,��!m�3���O����EDWo�(��f���k��f4��3}�:�!(��9��u����j�c����7o�K/��]v֡������<�c�@�z'��&���kڕz��yE^P�����=�hS3�]��Q�Ew%{�A�
���u���M�f���PF==F���]uL��<����5�i��l�_���/a����0ͷT߭Y�"�<�a�ך2ۚ��Cӆ���9�Z�����R#N�d$�0�p�MYt���DLc�$��褣����=���}���ʹ����vL��N;&�oݥz<n�B~c�G١�3�%, t�\޸lM,��b y`ͅ*i(*�����&���Y�Ţ.Y�B@���VcLS�9N�������k���j�ސ&)5rg������Ѓ`���<��ic���t����!l�\��E\0���tO5�kB�y������a��*�/��'�x�B�H���F9��.������QF�i�����=�����[thx�1B�Yb͖On��+KOfZ��C��QO�6r����F��A�b
����(�~W���s`ٚ��5�����ƴ0/Is�S�}��m��J����e�p�&ge���uȂ�戵q]߈\�aQ���99�YD�],MsϜ;'ׯ]�{�cF��w��e�<�0�x�����Q�F�w��������P�Vtqit��/:�&&�����4�`]�A�D��U����y�3�di!���R(Gլ��C���u�.��0-�m0�5g��u�lFj���a���)bJ��˺m��qR��mM���/���t�X�:��M��9]�xrDڊ[7�ӆ *n4�-X�7�/���<u��6�OyK��M-	�0��௔:,
>?�=�P����tmA-�z �N���Ԑ��̀�p����K �� ���}%���b�����.< ��'�ڕ��Ʉ�����=9y������	�u1O:.�i� p��@��+��2�(��O#0 �A�Aɸ����
:W���jCD��:�;���FC�m��295C	 ��.aD���I�C
�4u�޺w�&�r��I��, �dw"FA�FSBd�Q# ��gN��c� ���ʣ�M��H�o���qF�x��֚7/D$��ax�൱�NgI�WbE	�p�0�0H5F�����T�E�	��x� ���Ў����c44|PD���%��5j��=�@�g��{@/P{&?4cԎ{�V��>F�oN��{�i �FĹw�@F�rB35�r'�'Yb����F�*��&������UF>�I�*w�v��F�B���RυED0`L�61 �|`ȅ��c���H9On��D`z�{�Yx!��u����'��"+�az� N#�0`U#硏�OÒbz�Q�w@���=���b���!��*���������[��+j��{����.S���7��{`�3�����k~�O���)�K�O �<5��s�mT��|D����U=�6	���=��W��O���Ď�E�7	���g`{Ph���+��HBĖ�6e:C�$�Ʀ dq�
���Xb�����F֚F4�yMo5�hAq �,�%:,L�02n�����K�v�'�υ�<l]�m��q�ZI1���O��,%�B!!p��σ�T�'E�U�e��"&<ԇ��N��)�!��Jq��Y� ���
l��п/L�0C��6a�5�s����C�ˆr��)9u����ϫ��+{��qj]�S�j}��f|��/�&.�A�`f��nVc����b���T�h4���
��̬*�.�J���;�i���n�	!M?hw̱��KR>&�F.�n���]9D1���������ݓ��;�ա�ӌg`�(
�4SZDW���م��@5Tt ĒM�(�K�*�N�M�
p����ל��ZᲯQ|���6{�z�y�y5ײ:�h,P�Rj�}Kű��j��HZ1o��iǢ���O���tk�h�������Ѵ{ ��7��Uc��'��]�������˂>IS�Z����KN�vdY�J���	�H���z��&��U������cǿS2"�0Q�ŀ!4b�k�:Xp��Q?�)\�F�Ŀl�g�E�Cvb��@wF��]�!�0�z�"�^��%}㔮�]]�-Ȗ���Z�l�&�(~��}@P�����N���F6xW�����Ұ}���р=Ù߸(�K!ҫI1�3qSl�FlST�#
@D�.b`V�iϮ,a��m�qa�����[.�ڏ�m��*���Z<n�\�� sUS�P�d�0��~ї�����V��I����,-,r#!����Ѩ��á�wc�kV8;;G<:�x�O&�`��殆�g[�[u��v�mع��?���u^���<�D.&�$��Z����,�*�=`o���]?�}Ӹ������SI�k�E>��~�Zz�M�����w߽d��ܪ�0����%�<�zdi^&Z����!��S�0���ۦG��Y؀�Rgw��=�b��ҍs����ݦ���e�ÇL�O�>Ǝ�4�B��=�Uy�4 ���ȼ)�2��3(�$���]��i�I�ac����52��zЀ�Հ,�ΘQ	���T�\ �(����g��\B���M�k��I�f�9���w5�3M=��X���
î����[po}f�zn�����e��E�g�{`@F�ZL�׈�Sdc���&T ��|�[�z�З���-���7"@5E�CQ���u㙁U��bg<g���|0������܉���hxn�e¦����	%°�yF=�JL3ӸNcu�wej�!��9�\��&Pb�o�>���A�I�n��7��!-��T#Y��XD� ����H��h*ךWk^�aoS_��\��*-:4�R�����\�ߋMueS]�ء�#'��Ŧ�Ɯ~���'#RsО�`?9@F,��󀛋E����U���&�@�<T��a󌫱�ӨF��D�x�8sK��bp�GA�=�{{���Ý��b��jb�|�ZZ�c�v�	��0��"�
:��m®�Tȋ[Q�tA!L<��qb"p|Ĩ�~��m��@��23'�~�#r��i}��4��"0�o���)V>15+����r�=��F��B ;)�N����="�����j���d'�MP��^&؃]JJ[fs�!`�0� /�����?�sޡ�8�m�r\	��cq~F>��O����c
p�Q�pM0D����b�2���G�% ���������Ʒ��/H\oz���y�Ѱw���9yꩧ��<#�������76�b蚬xa���!kkz�����LF��l�P��%e���⬜>sB��Ii`�4#T�L�h�
s�Rd�N�Wp���{ǵ3a�8�3�ƽ�o��O>N�� �G�5�3�=��H��
j$V�΁���&�3_{�u��_v�n��2�df	�}�3O��ţG��qR�:��h��w�H�+N
h�3�QP��_������lc�u�k���:�2(���'��m�~�Nܤs#�Rh�ٴ�^zYv�>�n��f!�t�ph2�)���VG�K���+�7rt�֛�Q7����>��;*
1�W]�QLᘻ;�p�8o�>�:�%�V�ȇ����ո͍{F��#O���{w��{�L%HO�{��>{pݰ�{�#�A..1���Az/�Ȯή��-&,�AJ9s�w�E��BI��R�xk��\��������r�|�v��; ��hh4��hnL�ʄF�c]rﰈ{�:�T���<w�� $��Fl�pAgC�I7RWF�[�D:e�kE�bX����g�N�ܡ4F	?}���ӟ�<K�����r!���4<��)�����$Æ�Z�X���[k776�w��҇z|F#��'��������A,vȴ��%�g��(V���ܾy[N;��7&��_�yg^�,H㑵l���N�u.6Sy�ѳ���
�,�Ùe0���s��� �BU޾u[޻tE�������c�6�0l&`�1x����krd,�c�3)@b�>�&��6��%���B7�i(`m_�yGb���!���p��<=)��ȞX��3�>"c���:��e�&oȉo��~]c��ؤ�D�>K��x'����J�a��ԔL��}��Y8yZFQ"a���qo��P2"��ӎv����zF�wF ��:5)<�"�X�I�3��\��������pW�ʻ�xh��gl�0��=͂߶���-F��!͑D���@�����ў<��'d��	�c6xե��o����m�����o]��WnrM˧��ה �YYt��^X(ha�@��_�����Ze�n��0�'2̌�=Mr����7�O��7�8�cJ�]�{Kv�aYʈ��[v9�d���" �!{_��gư}Z��S����l��w��� t��t�6V[��8lhM�bt·MH)�����ִn��uss/"=�4,m��{�/V3v�=�����o��ʙD\c���ښ��2F�A�'�����#lR�b0f�	t$nL�p�6��D�9�>� ��禩����ӌ�б�h��5�P�YH��4U�{g�ꬦŐ�˝��,b��J���8~C��H��t&'�NP�b(&1塍���c��a�n|����ʽ�W&(Z��5a�Ȋi���Q`���f4�H������(�2�lm��;S���������Z��������+�uy1����?vd�n>f�(a� � ��=�r�f N}E#Edk�;�@�L�Z�^��"%�>�A��@�ڨ5׿�/+��u����(ݦp=�0���i0}�A:*v=��uP%�dftT}Vӻ��"
M�r

%���
�1����>u�yر�Z�r]�w@z��
1����6��Nh�u��*�<N��?��>���Ƚ5���m"�&v�M-�9A�%EG�S���߱�ג���ˊs��[�g0����7ؽ�=)�l�'��5q�R��]Q/��O}J�g��k�\�������Q�u+��5Wԏym�X����牔�OUh,(�T����'�0�V�A��*愦�����D�y��Iz�7/�eE���*�/*U�1�C��bҔ]ě;�\p�N�`w5u���jr����´�fEԧ���d�5%��]�1]����f$�4��#MF���:���eh;<`�"�cU*j�J�X495MQ��uF�alH8�BxƝ��!����ѕ:�����o�3~Z�?���F7�3s�l�q���oȥ�WdZ����IC�cջ��� !*Bt�������UvjnFϷ�Q�OH�ea���Z6����`��k���4M���7���� Tc#�S1��Aa*���P�<�!����Ա2W�Q�mbr� ����"k[���youU64R	'���l-o������8�X/�DI���4����F#tbM�5X1`
��s��Ű��_탎ܻ�&Oԟ�Ze�M���]�FcRY$��E���:ʚFh0o����#)ܲ�w�
W���!��i���ٹY];e��\Cͨ}hj�0Z��M���6{?(�O�{@ѣ��B��7�ns9�8)���tF��(�yA,Q��l��kl'@,B�%��L�Lsey�N,��A�A�#o��kvcs˜2+@�<��`�TT���ؗ���FV��șs�{_��zac�v�ίd��e!}̒=<��v��dd��>բy`�>��:���Om�6��H�:K(FDl5�<�V�����Z���H�OK�&�\��
ć^���U_�!�ĭ7���=M�m"&.�������2���;ۨk�<��&��1�c�ֈ��Ҕ�9���n�."wЊRfl7��ؓ� Ռ�����+Kl�#���5=5����zB�n�#q��0��7��M�|�n�6�^�*�Μ���dv~�������hF���W^a�4���#�eB;3�(hh���9��r��-�����/p�A��j��S7��qW�;.���M��K/�ѥ��_C��3f?(�7>~��,,�xL��n��A�$�0E�U�N��:���MY^9B��͛���S`l�N����r�@�ͷ5�;z�9v���j�lC��S@R(�yք&���I&D�h���{l��=L=�R�m}��r9��j��1b��a����Ufl�q�Ե3�yKΞ{P��o����
�}$M�W��2ʙX�,9"�+�Fms4Xm����f}��\��5�N�z��}G������֦MN��B���0�L߳���,=��s�N��(fR���ޑ&�y�x��Ӡ���ҥ���^t625>f�X3��D����&���$�:`ò�,���bQ��ך��^�[�o�=��gߟU^@Q��e\N�ȳ(����襞l�b��F?��[Q%w��g�0�4-8�y�X� ���0�����8>�"��`�y�PX���k
iv�&��ٝ�����!zV�ů��j�e|Q�P9�:ⴈ~ǋ��M���`�ڹ6��>ǻ,�Q�a�� ?�9�rdR��B,3�9GfDqJ}�T��p�b���K�@l(���@�8�h�T�F1|�^vDs։�DBl��7u	:	z�衟�M353-�48rdY�n��A��$M���{�	V��Ð�H�7>+t̕m�v_�~�YZY�������Hx]F�$qn�G�R��?-5i���
\�����E�����5��22Ko9����-ȇ���� ��ds��؝�5m0k���7`���j���8a�p$��F�OQ�8���C�2M��"�5��j��3�)~�3�'ģ��`�V/D��4�?�����ɚ��QQ��ŉ�5��w恇��y��$7��Z\	�c�d��iu�G?�Fvz��L�<��=�$q^�
��-6������У祦N*s�e��|�dA���Č+���s��Y��_�'	�?�*�'����^X\������sQN��:������#*�w�9��?���/+R@#lx���<BT�k4;��,#؉�9���?%";�g���W���sR��{�.��{1'r����gW��̻��]k�H]w��B^ᕢJ�GȽ�F'��p�m���6��j눤����Cz�1>�ɲL��4*��8��i(�K9@0@a:#N����
!dYɐ(�>�=O�լ��H})�$b��ޟ��	��"�|=e�˂F�+SMiECN��ؔ��C�����̠A[�\���c� 0�Tk�@�!y�� ����Ss.�a���0?/���,f��6�����3�oF�z��:�z����gӔ���@��7�W�P7�@��p�+���5V<�1z���N+�3v[H"�N�	�Ig��I�⦌͌�SO?-�K�r��>���2 ���K1��T�j�;���(b)V�ѳ��6I��Zc�X��2۱;���k���c�>+��){Ќ%9~T�PjA���C�5�x�32������6TҢ�xLHL�� (:��h.k�H#��Sp)��0�����29=�9V��f��5j��5�2�+�=#��4
���}A�IꙐ-��_أ����cP�|�a�^X�~4cCVX���CƃbR��a�P��-i�0�����Z�
oX/2֏}�9�_�{��]�.^C3!m,rZ��I�8�9�m���q�JGn�챛�����N�/��Oc/h����"&e�UR'M�5 -%�Ҁ&��~</qQe���9̼A����ml��c	aLB/�*&��n��HÔZ�9�{�S{��I��f�2��4^;��� BL�f!����ɖ~MQ�`08MP�
^1T�����D"-�>�2�E�����?�����
5prk��5N#K����$�=��SO���E?@	hO��`��@�5"���Q�(�Ǣ£�&���&� HE�����2m[G�?��ٮ�:�ȣ�J/�ߟ�������gϙ 
��M�+�ML|�1&K�G��ŷN�ƹh�Т*VIe!�;y��Μ9�.`�`4��!����Э��Cm ,&���l��z@�>��G�Enװ��Qa�e�6�:{��7(6��>�q9u��;y�"O�>� �����t���(�g2BQ\�4�iq%j ��c���v�zˆ�E�G=>8U��|��T��V��u���{��f]���CA���&�~���B=�w'f�O��P)�@"/��H��dܠ(!Df��P�]�x�w%�������c(��(!� �e���Gl�۷uc�R�p ���:-���t��hlr��3�
�Yݬ-[U\-����Q.2�Ff�D)'���M�l�Sԣa�L�%�5�@��tqn�]���؝IDF����hݳ:\��+�Lh�/�,�݆�vml7pA�	W����t{o��y(X.[��6x���*���D
TnD{F!�2c6��݊��vx��5�,~,,)�4�LCgof��f䅌�bY0�����b���cHi�x��M�B����D
,�0��Xd�cb�H�'4�j!���R���a]�����.w�z2匀�F¶��G0PF��(q�����4Vg8CL�rXk��g�`��xD�3�����7�K���}��-
}�;&X`Da�]@�\o�w��0�jS�2e(L�#e��P#q���s{�Oo�#Պ/!Vm���������Zz��}�g�r�	�D[ި"Aʎ��d-����k��ʥk��tC��0�S������q��2��m�`�H�,�Y�7.\�'&��A�2��غ���=��}�w��ߡhK(�F�[%��1:d���Ǯ���)ؔ���c6Wk�]�M�� M<�V�-`�cjxO�>��i]vz]b�W.�P�CD����/R�r��o߹K�D�Ԍ�L�@��1H_jdW�C;AȨ<�?�N��#=�����k���$D|@��!�D��✆�֭U�9�8��Xw��6������C�	�s����?��lln��Ԅ��KJGVC�B�0\z��Alꠣ���9���r獪�,��:��h/�s������7��,;���޷�˽����^��Hds)Q�42F�-[��?�/Ðaa~�o?����m����20�P�,Q�EQ�&q�^Y]�]ݵ�/�v�����8���/��5���Y��򽻜'N,_|tei�]���o��l��l',�!n���s_�����;�>~�BJ<,eɢ�)�h�g
S���ӽɴEI��N�ef.���?#�{�srg�.#�A�oŻ��E���7 ��d1�<�Z�=$_h�����7U1s#Ѹ������Di-*�}����QIa8�n\Ӌ�ܐe(��=��
u �{۲��}Y]®8�aa=�@�Bf&Ԉ��dY$��8����O��u�$����
p���F>˖����4~뛃2�׮��n6&P���;�������$�h��-U�Qi-���EeK�Q����x���IL��Z���^�?����;��21ɚq�,�m֝�
�\�ɘl�]H��@N`x0fB�u�z�=�=W��<X�a����(_������|��y��*�:��Y��F��3�����(�+v��	㺠kinX3��y�����	V���*���iݚKu��BWi�����݅��s�����,�����7#��ѻ����
��o~췤��G�߱Z�!�6C<nH�%�Μ�0��������zO�t��ԫr%&*u��<X�?��w~����s	�{��!���aƇK7�0���]�D�w܍���u�mΡ�omn�����P����s�Aơ'�N�[h�r�*EG	��4�	��a�gY9��%wb� <x��ľ��u�����Y�\�$��e�<��޶zv�E��+��H�cz0�9���rM�߸Ao�f�� �P������n��>�;2�J��I��| ���t���.&]�׾�1aV�L�ʗ�l�������|�_��7G�_y���r@ڹ��i�B�I���}�1��U�r16�"v�`x���;�TKb�tetr�:�����Ԙ�/��ӗ��e�{��

��jW�}�\�ԕ��� ����F�d�B��9zη�鶔���Aܔ�	�I�PQ3f�2�#'T�p}�\f�G*�ݭnbyP0,��C	20,т��� �b��m[�vgjQ��"#�:���k�ep�L�����@XX,�b�4����{Ř��F�i���b��LIH �5�4�T1�Q�5qzpx Up�Qb�sX",�0X�ŋ6?���̲�V�GW�hվB�*�X�p�d�֎K�b�X�9W�yz�'��2�yj��yP�QQY�nK���;2"�s*��4R!��Z{@e15�,�a-(ģ�н�s���Yϫ��6JD��pר�Z���ץ�>��ؐ]�js��Ƒ��1�U�R����xQ��J6&����˲�n�Ge��ᅚKB�j�������Ђ�"������W.��m�5=ds�JK
�0���D9k�3YZ�3�ͪ�Pa�O�#�'��$\0��bi�d`����>������vH0�]���Q��1��������z�����D}`L	s��i�%�+A�ݾW�ᄮ��x���O�me�1q�H��J�w�o�f�,-����i��7��ʑ��E���_��rO�viQ������$K�{��M���{&1�N��1�7�-�u!!�V0a85:�,(����hqG��L)���a�@@�9Z�L�����1^�f8����qAX�Y��g'�Lqʕ�W5S��=�I�nP�(4 t�/	���O�Kj0·��m�ZYT%���Wς�W�W���Ȭf�J��uy�u�(���ݲ��A�nX_�!cΥ0���1���WN�J�J/c�Q��j\Oǹe� ���y`"S��L���Rʑ!�%6��+��^{���&UYd6�̃T���T�Xh
m��Ks�y�9vck����,��1_-��3c#�9�N��{=�3�JSͰ��p������0��	�`��K	�ۜ$�ӣ������:�N�� D֚�PX��Ʋ�i�/��D��%�6ވ�\u1j���2:���.�n%�� �J5GE�0#�,yHɣP�2��4ƕ�̑��{G\˵� ��=L:���|m�n. `�9�q;-�j��u���&�@�-!���әU�T�j�ͩ-�0U�#�K2��΄��ܓ��Ϝb�C��*�U����P�U�mN��~T���`�P�u�і���JY ��P-pb sZ��&��W�%��ș|0ё+�+�l����e�鶀��"��N��*�i�獒R��5�<�%���4�2��GQk.�ϼ(�,��[�RE�X���s��A-mE�=���%�bĦ6��L�U�����-��X��D	��'k�D)���<7��녭+�1Ĺ��"$�֦��m*5 ��(�h#\���p���E��r����o��wH�_'�`[�k�'��|k?0V���x>MXNb��K$W6���J1^%W��f1�n�cM�f�� `i���s�o�/�k\�(�#˞D1ST�
�S]��25�{�jh�t�\ Aق��x���+���o-�?���d��"�6��/��Wr{;�,y������C�}D~�w˫7n�_~S[�`�6�
�yyE�]�*:��vW�"�p�m�a�!���瞓��m��׿��B��5Z��<��
��G������_��_�}��C��Abd*���2��hfU9
�޵4�u�����ˇ���g^���D��Z�BGe�G+@X�����n�,��.tAJ���A!cb�� 錾j�ah��.v��9�m��[-.�d���
��I����[0�Z�R�4X��E����pLd�J��}e%�X[I%c|����6Z5n��%ҩ�5-�wT���i[c@|f��&�-S���I�.��v?�bw��/t!����E������ʺ�2In������s�ׅ�R��u#g��H�m�Y��qJ�:\�"
+���������4֭��.R+�,#�WM�	'~A�s�f��];��^�a&Y�I���u鯳e�S4��S�ض���*e2���D�%ɍJ�(sb�[�7V��*�,S/�LX}/�aa8�H�<�nD�Ly!��/�X��g�U�n2xV@)��Ceۈy$ā�yRV� �p$���$����ߔ��E�w�) s���y�#o���������`��������{ī���1\�fA�e���N�ÂJ��?���0���,-C�b�	J�?��.\� �x�;H�r�}��kjk���K��b)��db�)�r�4�yyQ������'������`�GkĐ	�B��IX�S�c���X��j�&�c�&�d���w�").��c��eB����C0�Z���&�������e8q��#M!
�pr̒�b)�~׉%�V�s���4[L��UqU�ݤ�:�	8�~Z���0K�J�v���O��Iba�R�����{�'�t�y{�h �g�(��7*$/KW(~����� GD���'V��j$���1�أH�Ba]2&(�5+Ϋ-}=E��.�}꾧��~�=p��j�1IV*z�����C+nᦡ��3 �ia���t��|$S�w���8A��hY#7�Z�i��s�V��	�*c�au�Q'��͛M7�T�*k�ÐX�*+a�\c�w[V��c����$CX@�Ϝ����^/����=�&L�G���ޚ,���ſ���3מ��K_�{�m9���yG�]�l,���]�At4��z
���o|��YX$��3�+�pkֻ]z���������?�q����R�&�u����7&�r�Bd���@[�r-/䉍Ey�徬/N�����,ϔ����T�y-�w�94�c��`����:�� �N�rZF�>�Uf���/�ͤץв��[Z��T��%� �
2�Q�9�
7���ѐHcWÎ��iK��]>���4c�S�6{��В(�x�bsM ��rjC�VcRCL�~��ͣ���2�G�P�T�ҺkxQ3װ���W/Z{莆b��Þ՟�l��fS��Mx6Z߫�ekk���Ҍ
�s���CF�R�k�������ʸf�7𫢲ml"S/rv̪x�y�I�ޔ�C	y�U�7���f>DH��\�=C��}�N�:��a=>�[��+�V}�PP�J�]�r��
q����ƅ�\�oa;��*�JCP3��Kt��d�3c�D�voph�ĒUr�,�����zV~�~V��{LTd,�mqn,�j������;����[��?�grX��G�;�t8%�zcAj9��F�M� ��na��}���5-��Q2,�T�di5��8	���4UdXo�=��}v�T�§��˙�\(���>�yk���ڔ3!}S:t-�����U���n4�����aƢ�S��B.���3^&%��I1iQN��v�E4�Cy#H×�d�]�������+��6�T�Z������HߖY�͕�Xkׯ�-�����9﹘�8c�B��v;f�]����Yh�<��lT�ub��=�a�!3��hiU�����5gC���[��Sll��̮`T������^�v�
/��T96���mEl�T��G7�P��V�S��(D��3�k;U/Þц;�yv�3M�/|~+37�;[̄9j���xb �#�G2�T�湷���窎��z���T�t���M�˂��b;���W��l��0>`�C������3���'H�t䑍K2���ڢZR�ԅ6�C[���e��c��)�L���@��Ĉ�*T2���:� �|�&WZ:�Ӊ��@u'j�3t�\\��h����AAg�=��
qdAa x(�����N�dR�,�e�y�5�J����rxۓ����3L�u;
�F����zŖ�TF?�%?7.�2ם_�%��I����C���J���ʭ���Ú�L����3����y�t@�<��3�\j��' �QE�$á��),�)�h�*���%���lZz1kԽ�F�ٖR�HHlլ���"L\ө+���kr�J���h��k=��n��w��m��&���~l����I�Lb����o ����0O�����+�ZI4�2�E�:NH8�����ys�Y?�*�ט��&�O�|^�.���|�Jk��&�f�Um�f�Z^R˽~�����p���H�h�OÑ�["�Z���0��<K��>c}m������O���/Q	رJB|��; y�{Dug��_M�Z������wX[(E�ʫC�$G�J �Bhi֜�f�KD�!T"�~��@���kqqaI�Ptp({���w��	*S>��&�Jpz"�!v�N��2��7M4�:P���֬a��m]������i,�aQWo��������\
vu!c;��=�r&�
#���:B�%WJD�d�6#ffe�"Z�bTDi�����j%�~o�N��I�6�\E��R��(f�%���� �5f����3�Ǆ��Of�궙iwH��$�J�޵�k���4,�y�/U��R�g���j����M�|q'��ΙZ0\8em�E�˕�.��⵼r��vK�@p�q���EKʭ̸�%���*��'��?���t�S)���u�Z��1*C�f曏��ˢur(g�4�s��U�RoP��J%^�<Gz�Nt-�������y�y>�sc�"�s�u��B1�o�\+��t՘���Qf�"�OK�W�R�+�J��L&��{1�%=��g�R�gz8Up��f-t�l�$��=����m9�i�<�}X��w�8 �a���	�zj��R�#c%�@�&�W�8���G��Ɲ[r��k��?�eǅI��2����t�ƥ�JS���`K�(
�	���7A���;�b,���kK��7x�h��q�16���4�IK?�C�2cU�U�ni6^�ڵT'�c��.�@y{r��ōe���� 3��	Q�G���z{Ke&�~�T̩�µ���b<,��i�����OZ\�߼����sb����(�-j��6O��bi����*y��d�>��RE2s톅x���K-W*�,��Ô�ð�Y�㯔�(X�m�Xժ?��G��|�yן�.��B]q5���R�sg�����ֻ�����zU8򼾞��4� �Ϫ��^�}$�2B�`���)�w�/���g���ٟ�� (]w�2�9V$�΍h��y��P$6�W��ū�ȕk��֖�t���,�vP+�V���������?�#��؏�2�G���e��;���1�@Zg2W�P �K�M<b7��N���L��\ΟY&)���ڞ[��(�)wΖ�e�]��~�6��+��0�Œf��G����a;���������w��w`Mq�2�F�cE�:���Φ�,�!�R+?W�GcaGQ%��q;���9�%��?��<�G�i<ầ����/�.G�jL��kVy/o�H�	��cy�qT��nl�9o*oG0�'�H����r�k��x�)�(ܲ�f��潻qR��-�Q��� ��B/©>E%�~�hҶ7�gP��lN��5b����B���p"jP*	.�fM��y��.�^���_�����G~Z^�sW��������*�1��V���-,˕�ҿ�ݗ��.;�3X6wY�����%���$XN/�s�
�C�R������d:��`M����bG�,�
��9�2U���O��%��5���,mA�%��p��jTO��[�����YV	��I�'��y],0I
?\�c�����(6���J	Fƅn��*���	�hTa��5�⦧]�3�ACA��5��qVQ�~���VɦV�I�8��l֪L�=Hv����`�C:V�UJ��l޳��|��t;.4p�gq�$����5�p�Q9�(sd@2�b�4�:�7�>R��Ǒ��H�Q��X;p��9,z�j{�x��`nO��/V���4�1ږa�7%{�w۠�-���f�UV�^i�/�	$[ʖ,w�kO�J�/�_���u�'�Rltt;�z������.-`u]����,����v�.U��MiֲH�����HM�L'.-�k�_�+�?�օ�sA��Z�`Ӻʘw����}���,�����!	Ƈ�<Z��
��/&����T�Z���*U�1���} M"�:��۲V�:\��a�z����D�ж��OOWZژV��Kl�[D:��s���]k�U4��mn'�kZ�^�iQ7�?ދYOe5��gB,o��<i|�c�qo�WS)��:7��xos]�^�q�<�=�s��h�^��4�q�����a��n2�y� Hְ��B�<T�YU`+i�%j���;_�X����	
�U�D�ApݡKY�g	����H���vQ.TPڵ�]Cَ� AU�M'2[����y�����_h��a�\:��vH`�b�J�Cou������QEw���ϛ�c�xΈ9窰ѝ`!(Õ�%;%oA�{d�s��")�RVa3%���$L%�*:#뙘u��!��V�aP��4E���R�K���)�{�c��@����	�h��S��aۓnG�UY���3cˊ#N�<���1=����8k��6ϚK�4�1�n=��<9ΝM���4�����fV�<��
�^�A��~?�gO��yG����t�fx9:N��t�������O=6E�Ԇ�VĢ���@�{|)�"i��4e�-mnG} �,��hJn�̺)�"[F=T8�v�+�]�I"ΈY�e.��4XHY��A��?043��Tr��;{F>��?ο������!n�����w�~0��2���a�Y7�8��9���GW/�:�ؓ�^.�]iw��3BY�(;;�%�#2���W��%U��Py��,V-uÀU�6Å���|5��Hp�*�9ʄ�䂞eD`P)��De*Zj{ ���v
�L�����tOg��F��XϽ�����f�l�h�xR�y�y�7�H�N38o7cǧ��8.��|���q�ޒ5��9���i�H�ooUɽU�z������M1f�O<2o|2�J>�>f7�*z�X�X��&�g��F�����W���K�r����ۯ���{D��縐E醯NP~�K�pDF���aM6.�;?���%��[��������ӊ|�?�џ�~�I�-/���oˋ��$/~�y�X9���J]�`m=��c�K��Kr���ݏ�^P�/�aP�k���󹷳I�]��˲����l<���#�,��Gw%�E�6��>zCaBK�g�HSt RSd���t�O�~B!6��*����h��#�pK�dXş���Z
���Ĉ�˕�>w��7��(C�CV�TG�/�9�o�I
k�$Vfcd�{�3ǽ>���]Of�3���L�ϴt/W9�(=�}8�2;�~�F�|6�8;t�AVSc��+"+T�K���=��߸/�*��q����ļ��ѣ�qy�$��� �GZ4�`%o�Oj/��CmURH���rm���{�
?����2�o*(�sK������kg���=���������,,���}�Ȉ�|��6����X���d�ޅ|�_��O~=(����{~L~��o��p��Y�	,r�-���I+����d��ַ�)����X�zKt���#ݰ�,�x������/�;,vsy���#�~Pɰ*�SkwwPCeNP-���!&"%^0ዎ"65����z_¦��O��P�6
.8Σ�񈜂d���^hUFT�����,�J�Ӌ�E]���.+rm���@��=�����J��m�b��T&C�6��>� ¹W��d�`�ܬ`NC㒼D���-� <,�j���)���M-���u�:�*<2/qq4_Y��|?�j�%W����ɣ��-+�f�[�5��ϫe��f�F~*�x�e�9 �>RW׹Sa[��7��f��ϫR�{q5�%5�]	RT�t7�.Gp�Q���S��2��WtyI(/Z��*�˽�/ٵ��V��QX�E��<Q]Ű�R/��V���A��M�G�#�i���H��i���!b�	��խ�ըp,u�eQ�g���HKu�znU�1,�ܸ��V�w��/VߙX��b;�i���Ow��~��>ؑ/}����j�Pp���v��+?�?�>��?|�Ѡ`W�@���w����,����>b�n��Zd�^����v�x���=ebo�c�G
h��������GnPO?���z�%Y�ud�2�6j,K�)��B2������fd7���5�<]Y��A	A���),ݮ�^!d�����,X�`2D�1��G[c�wH������}f�2K,"�R�Zy}F&�D�	<^���J�L�-��o(߭T�Qe�������Iy��P���i�����J���l��}�-�lƞ�E��ڽ2k�+�s+.=�/�h�e3dD|V��ޓ����T֕C�K�ĉp�Z�����q�1n'h͠�P��ԕ��'b=�m��f=h;��쳶=�-���5W�Oe���!#'0J�'oQe��4sr�ʴ��7�d��������}^h*�A}�ӿ��q�C3��ENi�U�P�:NX�����vR��*�ɪkJ
1��{��9�����ݻ'߼u�qC�Oɫ�n���-YZ\�
��H�p��=�����GzX[=Yj���z���3?Df�o}���헾/ۇ���������|��o�G>�a9��n�TkT�|�mO��?!7_�5���M����Κ�5�mn��Qɦ�eu��ޕ��`�DMY���.fĘ��c���l�uYY=�T���D!�.�_U���	����j��N^ZW�	J�Z��^{�,��[����|n	z�R�BP
؉������=l0;�N�>����:�=��t�Osޙ{��.W0��;�}F���JfH%�x�sUiJ�������&�\�0����j�Lٸ(���lD3���Y�U��2Zh���lϫ���e!��kwCf�)@+U��Įו�>�d�����Qh�D�V`���=���o,��M��:�
i��q�ied��8�HCg�����%ڹ@�����jw�:���r��ⰌPs����7��R|a*����K������ܾ�����˲��&�g���׃b��g��Y��t�-Yo-�c?F���p,����o��?�A5dC��pݫ�.Hk�M�8�]!�`ŞR�E���/��^�~�5����}OV���_��6�I/�eh1�t�z��M߫��Ņ��]�=�Sa��`��ʺ�Ν����?,��-�^��[ߓi؄�[h���i�3��TGt-����B���d�^�ƁUc>r��Ę\fᎲ��d3���0� �hY�,��`���銘׬\���y�BE�B �&�%Q�{}Fس�1���qN�k�y�ްi��=Z�U�A�xǲ���qoy�����]���KK��w��3�Jn��γ�n��lS�L��B�{+"?9��4�T�%�5�~�ҫ�o�Kԍ1���YX�`�e=�@�/����8�ʹ3g�eK�ܙyT
}���C/Ԛ=����*��DU%�����xeL�نe����0�ڵ�*�7���'�jxpl7'�x�I�ᛡƓ\�d�7l�sA���.�k�ز-�$8Yt�̧Y�I ���ݻ��4�)'�����IyxnqUV�K�{��$����d.-Y�ɣo{L�;)(���@�n��N�]`Yml���l�=��b@0v44e�
�c��ܺs'��-��v7X�o�	�V5U�*Y>sFv�ñ��;lP�
�<;9KI��*P�u�i�ve�E�л�M���YT�x������/?��R�v�3�-P�;�ϵt
t��m�%�H��R����A�W�p.��s���(��b��?�dZ�i39�u x	�[
"
��p_.�^-5�{��mfXSA�7�o�hZ.1A���H� r�~eqIά�� ��ġVWW����i1��t�!��Pz�S(>(+*��<���u|fm����6�%�׽p�|<����	��v�����I�к��4���[9���	���cj}}�y�G�ԟ]�(�	�*L��Bi�˙�|�H�E�����Pń���pƆ*0A��l���餈u歌���֬�,G'{�5��;���LH�Gj$5�ѕ��d�MX�|�K,�O)y��#�/�\�{a#�t�A��j�8���aw��y_�\�,+�y��G�?���]���.���{���~Tίm�h���6`�>`�JАl�?��r/(����۴r��ec#��V��A��ل��);��E��E������|���&h��ܗ����/i�ڰ��*��;�c��3��$q�Hd���>�JX��I�0*�o�Ko�'��`�`��K>����o,�h"�Y�k�ͤb����z�P�%4���j6O��3�Z����%�T�2P���D��J�7T��4�������R�3��kY͜Wr����'���ül�l�U��:�`�Q_�s?WU�z��h��J��V9�兿C�Mv��Sļ{���5BI@���l�T�l��Ս�I3`����� (�Q�|ѯ�ܹ���}�1���Ӹp�!�z�*(6��A�A��k:k�pM��[]]���M��%����m�a?�΁��`W����;��r(�%��ϰ�>������K�,B'G�R҂�T�|�z���#�<��������{�4���lp�g����p��PA�����!�s|$�*u<�����s}Ấ��f� �aϵ�)a,Cm:[+ٖ�"N��L4���>+�?��|��~ޑ'yT����R�)��8
J�ۯ�����Vʌ�e�A8(��ٯ|����{��{�%�� �@﫰c����vtħ�%�
��N�!7�wi%�
X�/˅�W��[7�`o�q��7d)(���_�q0���>0p���v����C%E�\+-Q����+a���a5X��
��+;����H����~�n�N�*N(ЉB�@c8��T��0#	tƤȴ�����*��\��	��m�_*xB�*���~{s�e��M�k��P�^HPS�u�B,.��<k!u�Ra��O[R�
��3�Ѥő�Hf���g��%�<q��;gjkYl�X�9^��_���$�hQo��
�k�L..�	��``��y	9��S���l�T!���g�X*�{p�hx�6���n���!7��T8�a9�k��daa��&�*&���s*���gΝ��`�noo2FL勿�F�r�����R�J)/g�&2�_��^Zҵ���o�v_�Xp���J����iI�d�=ǅ��;�<�{��^&��M�Ϥ6��lY�?C�ʁ��`��5�]���_+��b$��ܟʸ+���r]@�Ͱv�6)�P����n]��n�V���8��-������M�G������B�Z�L};L޲,�WH���`tpH� �/ �;�y���bF�y$[[j@�^~�t�@���i��d��헲�;���y ��
�#[;a�'��n=f�ٹ!��=�}��ҷ>��|t(��V��'���tZ���T�"�)d�Q	�0.+V�e�3��#'�Q���w73���g_
���(����g���i��q�\t��:ޙ�0��	�9��I�<�������דD��s�0�Ow��� +�����wXQ���m�t7aIQ�Ֆ��i)�"���]��z�zx���W�}�����i�qp8
��x�	�ġ-g�DE����"1��Z�t�SkHK�rV9n4-�C��z���\� ����`e�σ1'��Zj�0���"n�k����V��"	����!�-g����!/�e�S����f��0�pĂǃ����BG�(	�w�cqԐ��d�L-EH�Š�!�r�l�=�.�E2$��-<���0y��P��3$��=���'�.^[`�f?��+��+Z�y�#ctje.&��c�`(�V�֩� �p�X!v���-�s�MZ���=� ��c�p�*L$������*吂�D�p��|�wL�g�=~�䠴��`�I�e�1w|�,l֕�éܾ��N���V��أ2*�as����C'�)]�)���CHc0BuU�l*dZba�8[BUU�c�Kziz�⮕* ��dzI� ��x��Gؖ�����lD��.�0X{
0�x���;N@�=��y�b�ܒYȟ]�����ŏ+w���5�,��=U�h�[�D!Bx?��K��������@=e/��/kq��^p}�j�p�#�ͬ���w�2��g�!�ω+�����a����

+�Q4D���-�t��@GFŤV��X\bY5���`� l��®��R�*I�jwx�"����6"hF#��\��.���-`�Ļ�����A�˖�!YW[�=	| u^ Kd1A)46��1�0�7cDϩcLo�!>Á��	QdvO���&������~`	�q�d1qAe��o�e,�q>��lHk���#��׾,?�ӏ<!e�����@���?%ۣ);��_�([�Z]�e�1?�a��Vd��(5c���]���[�����D9L�SCon�UE�[2�J��߭.O,��z�il��,R�Ą亐*�}�����ڭ;���q����l�X�N'�m�Ga����qp�$��l>�T�����o��QZf�JVy�D "�9sgMh�T�t%[+�Y��0�2h�������z*nēz�h�?�b��!N�T"�J�����q����f�.)�G"o��n�Y�AW�(z���w����n�ڀu��Q�pEO��^X�ck�o�2��1��J�У������?0���r>��<���lW�,s��C�f�����pĞTd��B����TVn:t�N�|�3kW�����G�L�i=O��@ܙ�o�&�$`�"$E��W�ʍXӘ�`4l���zP�������*�_�#�B�,Z�f�s&k���*������l%�<�e��D��μ[���9���^�_�X��2cQQ�Hշ0<�&�!���#�ٰ���]Y���c�;Kc�AX��ߔ��w~K�aⰠo�ߖrA�,�����My�On��4ࡺ­�NFm�2)��Xǐ*[��fe�b�+��c��n����f�f[�t$<��X�Jj��s��8�����7g�1�7V�4�~b���6��ww�ܪ�bw*]�=�hv�pC!���p�Iɸ��
Qk��l.Z��J�|���I(QEov���vl\�c�y���C�@>t�����6��l���[j�Cz�t���Gw%�1�K�4ߛ���r4�#�I�)��iſ�XYnNh�,�"��H�@V�Q#f�>s�#��P�Ӥ� >��\�b8��Q�wp`�23�h�ZY�أ�F�f�n��sG��ܿ|�]9䦠�n�>־�ͮ=���5���4��
��P�]�F� :aM�Ah��"�m�U�P1i\��4��J*W�6݊B�xW$ƺՐ��A���]�S��s-'����.G�C�����))nZ��8	�6y��Uf�+zT%Jv�f�Е��M������R%�XM	�Zʴ~��&�C?�Ay����[�n˯��?e#E_�i�ۭ�y��m���w�K._�,/��23��hϟ?/7nܰ�E�����W3Í���O?��|��_���1όPR���^���0����T��M�lw,���9�PRT���Kf�+�J�F�ʨ`ǀm��E�[�`Y�U)����r� (�,��[��K�j��ƞ%�� :ă�=����ʲY~���2�uc���\�1k�x����H�+�ܿ�`��
�cȚ�h�"�]�XдN`9�^\��dDˎ���,V��Qj_5O��E�����*����X�VG�1q��/�6���HKigw?X�CC�0@�g�^u���9q����N[{ϳ�f6<�޿�w1l0:��:I7W�[W*~-|���Ӫ������q�r UB-Z)Z	
�V��VZ|W+���<I}�ei��JP��wp���@1�{`�+Q�i���}����Ɨ׹� ��4���M�s8s�\R���a6��B��Ƀ5�A�jT��$%[u��s��w�O�������²$_�ꗂ��"��\�����̢]��m#9�8,�_��_�_��_�;����Q���C ~�4)���s����5ށ�i�#ޯG�x���pooN��v��JƝ�ŘZEw`jn>,�Ѹ�P1��h�����_l��b,�8l�$J��|<�j=�$KH�!�k���� �`��\���q?=żd�<ři6x��G��Cs,�����ռ�t������Xxa8P�m0:����
߿�)��P�z�8h����e����!\nXwi�N�)391�@ˠ�Jp���F��*ٙ1���� _,�I!]�ͬ�I�����B_�a�����Q�إe��L�[:w��R|��x-�k��4|�f=nT��ou-����u����|<��tF��Kʞ|�B���F�x���ɓ-�V���v%�	�c#d,�M���W�F�b�W����c�L��֖G._��<�.�z�!y(|]8sI��%Zc�!��Lޠ`�牦t�b�X9Qy1��t�|���'䩧���^z��ôs�-k<�״�|�����.-�M3�~��1��bM�2��_+k"�Q�I7��}�;�bY���t�U|,,X�� fh�)�¤T�Xĝ�U20����*�J{�FK��ʯlsv������ ����d�k��~�]V�Lc���t��MoZ%��|�9�nM���:��Pj�\��Lk�ݷ���5룗[�<�B��hfx(g���� �T@��VnV���L�\ ��kW�K(K}r��wP�]��,��������?#���ѭw��������[ȇ�`�8��#���������2ќ[A�U^�v�w����)X�����㜗�ƙ'�\>�����I^T3w�/�õk�:q�>��ƹSK��̼'Cdd�B햖䇞}2i	Fr0�հ�.�_���.ʓW��ӏ=!��/�B��DU9e�2�W��bi��AZ�c&E�R*�"a5\��0�N,
R���E�'n������VCj��w,$����R7�cDZ�UP����9�B|}7l�3�eTO�Ω<���+���"���Ś//�9�8bp�U��]�5��3���&�E��xg�؀��}�Z
�CB4DF�%�xVn�<u9a~�$,�*��,��%s�Eќ�y�J��7�>�PFKK}y����q{�dmss_۸O+rv,���l���6�RoB��J�4P�bΞ�ށ+��e��y����.d��Z�|�,������-�KBE�:���k�KShT>c��oP�~2ͅ���O$�GB28э<@x���[�1�.^?��$��eU���8���%$dlh
���F�>_|�T֜�H���&	M�����U�����^��+�5��~lʘބίrJh�p�������D�d�6���X�q�q�v�`�^$�V�j���0*(�Bv嵻��;/}O>��/�0��������Y� s,S8�2��(��}�G�'�'��_�r�=!>%��~�|�va¤x<̭`��
Ïۚ�b�t�@���XBz��6�=*v����ƁB\zm�]q
�)u�++,`��UqAɢ�S kvjU]T��v�
�g��g�ĊM��V
3o��R���A��6J@�PͲ@<�J*W�21*8s���ɬSG3��5CD~��߻wO.^�@Br���^
��]���`$��I�7f�;�5�yGv�$K��tO`&���r%+AZ\Zd9)x|#���۲�!�XT��={6|��90�^Cd��uk_��I;Xc
�k��#�F��-�����j�c��mz�����<�X�b�5WZ홐Eꍸ��]���-{�S1��ȩ��|m�&��'Vq4�雇[��a#u�YqÎ�v'%-��0A�ܱ��J� f��Շ��3�<%o{��Zɢ4v)����G��+r�������k���{�p[vF���#/�z]^_7�ܒ�;�eX��&���o��q�w��w���Y�цm�Q�2�믽.�΂\�p����>�� hZ;��`�\ۉ_y�
� mµ�f(}Ě0w��`Y�a
v&aQ���2 �ms�SY�l�	��d6``.2eZ�
�7����,C��pY�K.I�Y�ʍI1��I��$T�y�(Ɣ��_7�9�3yn��BM�Pl0�)N�L�k��z�R�MH�%�~2�>�x)QṀU��8,�e+P�T��P���b�H����&.��=7�pv�,2Sn^YE�t)��oq3���ev����0���w��ߍ���.��A�Y�4�[g�gTj���Z�Ab���c܀��c��;��2�,�%���\-2,;��������UJ]�h�zuO \�'�b��H�ׇ\o*&'1�"�M�Ţ�"G
=���t�h�*���$Z��)��h���?H�4����u~��W�߉��hx�O{�7 �A��������]��l�Y
�r��JNٵ�U��y��Y����O��|�Ƌro�+��9�J��	o��j�嘨���<ovP(��V_V�EiMs%�	�R�O����?�gV��3�<t������T���kD�B�v$�]*�5h��p�	�[��\�]�t�}tS���a�H�2�_T�,�z��H��X�F��5�W+����v`j3��̀M3s�iy��Ű~i�+�D+�J�ݢ�>�^1�������M�����U��S�	���9:�T��uθ�5ʬ���΋���H���52/�T�"�]�v�j��3����DzE)wʘ�����gu*��.�w$��VZ_4��mt%?7�R̩tŠ�-V9�޴�xzC|8.����&�;�٪�Qn��8E)o����"�sP���
�w��t,v����\���E�(�@b��p.�<��-��U9����RU�iw���i��Y�|��ӡ�]��9O���[lP�G�wKNܹ�M,9za�	�����f@0�LT�ܺ��nc��^]�Z���f�f";M��"�!ZGTD�`-L�  qwx��X���>��s6:�:�m��@�W��7�[�_N_�ޥ+	x5�`�>� 啵dz��u)v���ױP��2�W��&f�d� �.��W��i9�C::�����������HE�+x����쁭]ZÅ��ekg�ma0 �@�qg�;Lϲ���4�ts�"gQ��3�q�|�0z�a����U0|��m��+�0c)e)
ֶj���R2����_��R ��-���J'�%Q���!����Ƹ�a�̳ͨ��DE禵TU�ѿ�c]��(����)��2���,��c盈�S�3K�!(U>�ވx�S��-��	����~�w����*��6�er��ʺ���&�[��pd�{o��Z�u�U@*xoU�_�e9n��Wɦ�6��iKK�)�>��v�z�NL6X|8���G�e�O�kK�"������h���*��(�P+K/}��0C�7��V�z���ܚ5E\X�='UeGCQq�Y���^C;�Օ5��_�B�]����ݔ��+��3������G>$o���W^�oܐ�v]nݹ%;��`�2���q�+7.���m)��'AQ�"
$YZy]���lY���o4��t+(��&ZY����ߎ����9��
���6H��<����KOIe�@΁�`����'�tJSB��@�~��0��\A{ʭ�݅Yq�(ٹ�����=7O�s�ǿ������X��ud����{�fު��DE�b�{��x�4��Hn�-����ӤL�ZVb/+Ov%�˚�'W��ƿ�E��=��Y��[-^����C��w	A"F�(��zC3M��fm�vaۢ���5��1�*��*4�F�!Zx�|�Z�@I�d�i��N�\G�BE�`�c�=�h��P�{C�Ly��ټ#����j(�2dyY��{3�.��]����3��ū��ÏɵKW�wF;�.-?"�]}��to�<������|��+���=)�G����/^p��=Zm������r�M�:�8�]���ɑ
�7\DŨdR�+�[P����4Bn| ��������	3G�B#�C`}c�����T��V7�#�W����W�d0�+�����Rr3n�&�M��{r1c��~&c����Rڧ9�s���#��SYD��轨Ǧ
�J4�[��9V�^	���Js��N=��j+1�3�g�]
�f���Z��_�?f�ݕM� E�����>�	=�C�hn���Q���Xi4K=[��F��CB�yU�Z۪���>���dv&�@��h�Yk���WWV䩷=)�n���C#02ZJ ��h��H�^nJ�\>'~���;�k ���ii9�J�Nn������ͦ�/+�M�Rɵ��
��>Ϲ����a������[/W.�mȳW�k��+�ɕ��i�.������G���O|��?�����eܪ���V.xY��Dh� UP*Y�����!*���*V2�2;�`���P	+:-��\}��p�ҔL!E8n�ﱹx��7�S8�Z��..���B�$!U� ��t7�,��9d&�!�("�'y�.u�R��$���3Ou��j��q����J�qn����;�q�I�o,*K+N[#3
��U��lç Eʭ�_����p�jy�t��BE`�ȁ[���J�e܋�$���qeL�
Y��V��U�0߅ ���q�Xj��r�2��~U�?��G�	�wz�ْw���nY�kc�d0yG���r���4,�t>�9�_�����u�An����&�RB~\	��H�I�P�߇�_���$YK�1�;�(|���X�j����c�]6�"���,ׯ_��^W|�߇��[jɫ���/ߔ'.=,�^{Z�x�Q�v�a�z�rP�$E��k��ޗC�;b��7_��AM*rpp(�%.�l7�$+�q��I-b��Y0��V�C���;,fp ������F����H��uT6��E��Ru���A���a]N�+�exg��ݺ6�O+���yF�B��b��vZ�4b����c^Ib�[�IG����|�'�;�P��s�����������ٹs�Y
�u$xP�iʙ3k��1��Cr����/+�a�^���5�%w����.D�������xO��u��G&�.m�(�۱�@ �o]#�F	��?���k8/>�E�1$ׁ���]Cd `i���r���T8V��W�i-�5������Y�U��#��ϗ��I;�Vb�`a)q��:B������ X6�٘��#�̻�i�f8�6 1Gz
Q�VG����Ē�)/��ޕ�_}�V�Pb �-0�N?�ax�w�^��߼!��O�����>��g�-O<�6R��%�)�FXsv�uak\LB��֕CGx�u������j��,���X���3���SI�(�2�;���4G&�J��cUk�����"�Tz�q-��3�lɞL�7Uca�r����ъ�{��R�y1>��6��p���	0DꝾ���8��[��I��
�y^\�sN�6�1!}���bO[[_a|�
���ȽɘP�%��	�mog����9�tᢼ����?���~h���~�F�d����衄��
�t����2�Ne���x#��+���`��m��:0��������g<g����?;	ϼ�w������.���Z�2�dJc���r�cB�E�6�X��he����&��/Yw��|b�$L0���ݲDW�F�.�:� �F]��_��R�:)��hzL�Vc6�C��DhE,���Oj[��*�;�]�
c��o}K>�?�$��$�Fd(��a8�1� ��v2��^���_�o���r�ӟ���=)?�C�=X��R���T����I���_��I���^9��N���-�p�G0�W@�hXW��T�������5��$V,���+j��ϛ��j�<���m}�� Z<�fD�>*:��J��k?����hbؚkָG��ٌՕ��3;v�,���?�O�3��'>!������{))�2����Jb��f8�qi�y��{os�=����ﵸ���XP:�ڂu71X�R���0\�
tkK�����|�*�M(� #��X����#�P�p~'u����C��q'��T��ՠ�Ϭ��haD�4Z��2��[��O�Mpzl(�}�t$�;���=����+c�C�� z�^X9 D㮞�T�7��2�)�ˋ�>f+�%K+c9w�7!��Uƛʍb3��r)�8%Ή� �.�w�ѸbXgj��t�3��YH���L��%O�t]kDe^iEqyt{��0��r�s�*Y�oY3�eV����������/'T�\Ho�x-���l2��|eA�n!���Ʒ� ��f@[b3}a�A- S��O��q�1]��fև�ws{K�� {U��Z&p� dkK+r|�lY1�C��%.;ᡷ�N�e�q.:$p ʘN��L���UN&�S�ՖH���*ʋItܖ*l�FYl	�.�A;S������L�EI��{=��b��Y�%��Y%S�NOh�v�n��S2����0�^�L��C����׋��/��م�@�Kb�����zH�m�s��S����b؄�R���!W1H��x��
�Q`Q♈���$X< ʣ>�jɝ�������X�y��a�R���r��ue����9E�I�m�� J��LI���d4V���|n��m^���@R�L�z2�9�ٽa��"/,
�%�n�Pzx��`}���\�ª�W\)\	����-@ƠY0bvwv)�Y+#w3�{euQ��w����z�l.s\G��z9eg��B�����9����E��Cb�o��2(�'��������I^�L�QU�ogBkR�`��~Z�V��Ɍp%[�e��
� ���5�%ğ�]����ݭ��ϔN/3Z�����i'͛�U�0p=�:��H��Wa��!�C/!�����C��.B�0Zݺ�J1N^�(����@�rUa!�.����+w7��L:�A-)����)�\aWLMk-�
�������,�E��nj�;���f�­��lކZ���VF��P�6��EYu{��Cf��s=yn��'?��O�'?��Xf����Ą*d'�]�bp�)�f��ߨ�c�~��Rh8)(#��Ye�x�C����b�-��Y ���XA�ńD�%�q;?�����ëT1A��&6vYT���l��;;h�	%�E�;[�Q�ăB�ƕ�Qf-�,**�P�^%\���W����a;�r���Ƅ-���j�n�m�+���b�9v!�dsk'���9	����2�2ܲ�-�z����4���%�aNz���ey��k�P+�ƪ5٧�GR�q�N���ܽY����Ol�9G��%���<9sk63����t�Q��Ls�4���]��b��	X�cV����?�S�C+fѵoM}\�L�`�O+�L"|�u.2�쩾w�l-k�1���J
v�n�a'T`�u�ۖƢB������
�n�	Cf�'��56�
w��˕:�+���JStDH4��1v���T����T� 0-
�L��Ը���b�f��ػ�ޯ�X��1�$;|���P���w�V��BXcSk�o��i�'��u�8:��'#��v�z`�s�-[l|�n���V��I�	�*V}y,�����܃qNX�޺�N�(:C{���kXӀҭ��͵O��b�J�0��kH0DXِi��5C�p	\�Ä/��[��b͂��V<ƴQ ���y��O�(�`����<Kb�h�уrx���W����"�k8
�-��=U�lk���Q��ߥ�¹�R�5�;z�u��z\�������|,��d��~��NR���7��b:j�U������$ǫ*~���Eך8��0P� $._�\�}���	Pl����~��\�3g7��g����f��ww��k�Y|�qF���`�jr����#c�I�C� ��n�& t�l�d#;ny�@X.J�Ůt{K,�TNKb"i�	�;���5���4�$2R�e��C1;���� |q�Il
�9��=���|����0�F�Y�%Ű`A�����mU�ȥe1e�/�P����;��+���@�+X'#v��\��06;�(��9�t�O��a���'�����l~����;ŏ�`H�I�>���A����0 Bk���/W*�N�įI����k���������r^5ƴ�Ѿe��B��a/��C����5��jWj ͳX�a���d�x-���f�Y봬a;Ӛ������)���/�X*Yf	��5��B�ep����n��Fw����'S
/����Nk��S��v	m��p�ֺ!��`îp��9w�ܺuS�|�*䀤����<;A��{ϿH�	4�sAI�G�i|�SxX;p'�hgS@Of&�3�l�n+k�a�[B�\5.����f��+�.[2	��h��
[�1>s��u:r$k:6�\�_���xC���sc����&;�i �M�<����L����Sq2�b�'���\8�LoA��iY�(��8�C�$�NX![[[,�jo/(�ñzv=Ƭ�*�/�yp
��@S/
�U��%�����Cna��'oqLj���`�$C�c������K�3r�*&|5$J�vi���F|cu��7�6)jf*��*#i<�1,=$��g�3�B�	�Z$��7�1����YE#ʁ��o�ǦR>v���?��4l�2�|'��h��e�'���Ә)��_L��P�ϸÚD�:��H�K}B�SKߪ�<�DY��c"���� �;�N�I6/�d]�x��?�7~F.]�,���� 3���-7���T��o�.��]Z�P�]yH���rFI�8Ϣ��v�K�� �]��L��p�v��"%�Qa� ^�;�z��tîbhE�L{��[Q�"�&�����*�sG�v�����ʂ��U6#�f
�u��L�խ�PS�aӒh
m�r8I�S��s���P3�����p�aс:Yv�{�,�V{��v�t�1'���hI����t3̭.��
���&9t����0����ܜ@�}h
�m�`�����I����(-F �X���L�NŻX�]��j�u ���X���y����qR��a��ՠ�,�\X'���}�;T�*�YIc�%V�S�ՆV�
�&y}1���glz�f\�j�'���dSK=#�拿;S]�?@~O���yE@jhX'��b}3\x,��fˏ��������ꐁ��ͯ�!�H�~'�ra�[�X��#A9b����^�}f&�����pv�^xO���vA0�ݘ"�		W@#�ɽ�F���るcV,?0�t<�3�3*&�l�v��0R�$-���j	�<��T��+/�����mkL���~o��Mc~G�+�-u����
�P�oP�))���,��..�>o,�H��H��B�x0�e�;�0&Iv� �W_���Gl���A6�z��*�
>�o�nDx2


<�Zh��"V�7 6Pm���#�]Ӿtpq.`l�,�|���NG���󲼲CS�dއ�Y�n^H���[�i�j�I7q��ސ�&P]�yG��LG(xq]·2&����"zj%;��l:��x��` ��,���M*;鸥��[�Ǧ��o����2���2�O�L��gq5�a>/&��^�tG��������3p7S�^QZ+tI��*���ԓ��La�����J���s��ϑq�_���=wF��u�>cq8P9(�Rp��tH,�h�y;�I�2UY��F�{��:�R���L?�q�N�GK�w	�(���[�ι8G,T:M��889~�&�*{�킓Z6j������ȩpE?=z4��y�i�q�g
os�m��a�k���t�RZ��v<���.������VPri_�iyz2�����51���ޓ���\�|�	)xؔ����e��ش��Т�6HǑ����T����\�^Z��\0:�d1^P�ix����id�%�)���Ƃs�a���4���F�� �B,u�b&C)u�UWό�������|/`c#���>|�i����c|R�����ϞZ�5�ϔ�=C~y����媤F�b9*vǩrAŝ�L�V���I��T?�t�Zh�L�\�Ow����n]d|fE�ұ5�T�;r�������lPΜ� �09��"�Lbm�C{mY\^�'��w��n�;N6pf7I~�_A܋�+xv��KMn8X=���\�����
% H�%�[:%�`I�KQnL�7�A���DVh(�6�!5� ���Ea)��}n�EU=��FX��⏅a[Y�����VVVo2�y ՜M�AI������s�,
5Jb�D<��|�C*7C��J��h3�eOb=[+��X�\c`�|O�,[blW��.7�,Y����7U:Ax�, ]H$�V����UB�XD1��*~w�2K�c�N�%o��	�UQX|_rB���������ږ�7v��\�Cq35����EX7Cz��`�9�-жA��?�;C���lNcd���<�v�y4����;C�[�������jl�)�e^��"�W�}�1�}U���k@�^)��*��Ojum�b�Y0������&1�L�J�����UA�������PȠ(��8�?_�
63��V���X��7�&{����U�>6��Ͻ_n���Lv6�.-��W��/L��{�?��o�?�x��@-�.h�J#�q72$�IP\U֦XC$����C��V�^X��g�!&7�X��k�GBg�����_������Cr�n`c�D����{���AkG�&�xp�LA�x��F,	����Bw؟ӞEטr�B��(G�K�l���RNT�ݎ�m=/�;�;Y�OxwOq`�a]�?����<R��P�hK�9���_H."L������@t��_���9Tf��РUU����Aq��������������6���.�.Y2$lAA��5Wt�W�͋{�ak���FЦ��܈�&� �^Pz���bx�=Vk���C��q2�����2�3�c\c��AXGg6dyi������><�%!��]#|���Ly�>D[w��h8�x�v�3�β�L�f�H�P^������YT���n~�.��*�ѓ�l^����i*�̔}�q�j1�-�c��ib�]/��Z\Z��n0�����b��7ӣ���6���a�u$%FA峼�"�a���	_»��(O?�v�ȇ�r��u��W�$[��2��bi�`ڣ��/+�g���ЃvFڑ�-�Sb�H�R�/�����Nh�r�.�i�&Zx��I2)d��{=v:(EXNUP �����Ek�>�+!�� N�msHx1��xO�-��{�,IG<�U��F"Hy�W��s��}�e�'(�y�œ~n��I~ܢ�4�Y�A��꼿��X�0>��T�K�b�x�V�ɥ��"��o�����;D@3��B\Y]��5�
qT��{ �	����/�s����dc��Y�a�Ѱ	�xl�i�ܹ�ſ�o��5�(���
ʏ]<�b�N'������V��{J�����^�n�'q�>-b2�]DI����5��鹠 ���>-��^�l�=6�yBynw��ɳ%�J,�a��]�BmʗǊ=<���(�9�jʝ�[J�t�1/��&���Vr�G�?�dzdr�u8��B�L��,�������j����e9wv)�A������<�����+/ˍ�/ʍ7�X�6�|��<�N��;��!�'��]���X:�1~僘9�CY��n,����dh��b
���ۊX�tD˧��k�������{��*�EuR(�+~���4j��A���O�i�GI7�����0�M+�NKf��q������	,$z"�y��KF�o�K��ʡR��7���ͭ�1ܲ�.�����@z�A�E�ʝ�w#'���4��rsk�a���'�P�3���E��$��L���o�p�O��Os�"q��Ylk(����}Y�تg�Q21��rj�D�L)ںn&���i6�V�=�7x��"N91�m��,vk�c�Ҝ$MTK:6�%�������H�-<S�7���vO�-ߚ��A0�0���GN��ͦJi���$P�H2�b�ߒ��>$�<yY޸w]>�����/v�ʥ��?��Is������l\�_�o���7_ ��E��V��B��
iƔ2�Ϻ���7��SY�r�=~��	p��-�[��_P/��ʹ6��Js��D-��&�4vV���5����a���𫳐�X�R�J��+ȦU�ϔ��V7�yJv�{HǈC�&�V�R���f�4A�Y\nN�G�mZ��"�G�޿�ʲ4�]z�'o$&��BGY/��\�(����S򶅚��9�T>�p|�a�xx������Js�x4Amՙ�ϫ�"�ȓ2]�����Բ��la��?�r%���։9���w�j!`��]�3'�ǜ��BO(��Z'����Γ��ԴX�m\������� �<�ɏ��L�!���1��N�"3䄩�2���<W�`�m��y�'�*Sn��΃EVi�M��"������]y���r������}��_|]V���g������͛7Í�g�b2&4:��zI�z��f���ҒGw��I�d��#�
�7�>���@|���B+���QqTBI�?R��L��q<tp���i�h��ͦ[����՜{��#7�V��,�0�/�4�
R���
ͅ�������ĽY�-�u&�v�s�;OUu�d���5���m�5tKh�6�!�6Z�6��`���n��n�Ԓ��'QT��*�V՝��3�^�v�8�d�{I���9�s"v��{�oM�Z$u��56r��9U�d���[�mZ�U6d�A[)$݂���w^����� ���)�{�����w�=�LUe��JS��d�����5��\����)}���z^p�{S��3�WF�����k���d_�u+��,[S1�ZR-�^*SekXf��2��?�&�Z�����e��7�J����m��H�s:�Z�[�:��nȹ�����IvA	N�KD�����h����B�̚���N�^~��t�u��Dѣ�!=:8��nP��#��w�g�����}��U�a�;lN] �R�,5o&Q�[-X&��������_`S�-@�f��4�Ř	%�A j�<3C
��F�b|�&\S�G��&u��^����Җ�S��i��D0��`Q�<}��7k���,����5�rwT�c�����z�ϕ��*��!/y���"2����ֽ�����!����}�^�9�T@�}���J���,
&�
�h�c��J�W.>�tm��W(�ʅz­�5���}��vo���'�\*��s�����6������d�yn���J��'|��c����_�ʁ� �ˠ�f�FH�*Z+�t��+�_ݦY���GÉv�E>ݓ�o!GF���h贺�e�UL�N��2��y�Q���Q��HI�ߴ�QQw>�ˠW��I�����3����5���.<C>s�<:��V�篧�'�)Ҝ��ާ���,��-=MZ�D�B�jg�y-;��D��hȅ���2>�j~S.wq��F�Q3��}�n������ocLqX��#�|��W�2�B��v�e��?���l��.S0˭�E!����a��%����)��G^�HȎ홁���'-k�ڮ�=PC��~=�QjY$΁$�[�hZPou�z+�4a�ü>9����I��R�O *ټ����)fv��ј~�*nmoH@���;��ͱ�i 	�:̙gAUu����J���#���)Y
���������E�����4![ĠW\$濭��!��e_8�{5KQ�d���?ov������"�ya<?������ZzjEu��E.D;���W�Ậ����8U��K�I}><�,s�j�I�Ug�z��&Ī�d��a񓋙�oJcZ�(�6��yI�"~�N�T���4+��^-��*��I�)���R��[r4�e��'{����y�uG�Y�	I��2��t_�͛;3%&r+^ʆ���4�����޼DYع̭T�6��H�*e�y#��UZ��)�H7��_ ��Ј��b�R~�^g�Z|�n���I˟�7a�&$��ᄆ�������ȁE�[�Z�/�U� 9C��_��t�|��7nН;whZE�	���.�ή��$ז��e�C)�t�ҵ�����M����֨WyMGȵ̵#���Uf��7�F���EP��)��rt̟��H[9 ҝ�����M�4 3����*q��x�+l!;�=��B�R�?�I�9����TwRV��q�s���bf���s�J$n�r�5W���k�w'=����/�_7�߷�C�����?�h�f�?�μu�#+�����ҊW#l��q��E�߲8" n.O�}֘��D�7��1�#E����''h���5���+���LxA�U��"[�\��BV���_���F��J�V5��gW����L	�p��,�LUT���`˸��?T��N�}���ZH�x����&����^���{�Z2���{wh�����1"n,�Y��<GU"�UK �7��W��ɑ���~�~�������>~D9ꫧ��
�h�,��Y<�c��SmH5�N㈫�^���8<�f�!��e!sˡ�-���J���P��!AD��ҥ��2ꦬ��T6һ����7�R�UGL���fYҴL~͂=GͶH�4'�o8
���ԿY��\�C@XK���Yf�VՅX��-R��<��(V	z�,��#�Nj�C�}�	��r��(��g��B�Ru���r*��G��e�O#��[�9�C�y�K*���o������@������:>�hv>���):P�+�JxU��Erb��0���:��l+�
�fP�c k�|���SoI��E���#o���;�n�{�ta.|-���=�H�<�SCz���_H��`��<9H/��P�G�A�\�I�CWmݼ��)��a�K�7���t��V�*cάo�g������g�������8<!��GjZ�b�#��b=e�5�f�}�MqVzNp�S?�yyo���t���}Y�x�fr��?/�|�7�~Ջ+҂���n�L��PJ�/YES��Sv$^��\�2�<��B�"�:���|uq�R_(�+���>Q�5��Ul}%O#����˾�>��3�Ȥ�I���Qt[a�b3��A�l��������畀��XN���I~n+�Ԅ��67V�3��Yz����_}��܈��>��M[�r�vc�O��E�Qr���x�My��_�"=|�@L�t�dG��,���H�dDO����)��]1�f*��Hh�N,���R�~���/)cd���w豼^��ӟ�)�)���	�nz�{���5�o�\�$��c2w�>R��(��(6o�%�A}�-#�mHQĜۅ[/5��y����7[�6���B�����4K�Έ��?�4A��z���L��B(�]�}���es�*�ӌ���j�m�D��{��I����x̍�r����V��JtzOiJWw�A䘽1PY#Ҥ�*��=~a\wumM*�m E/q�䳢���;N\��h�T�k�C��>��� teʒ�2Ч�����M�nG��bZg��A�S{�ɥ#8'��VV������EYg��ރ`�X.u�A�
�d"�Uq�DɞN���42Mq��c�za�A��.���2G覄|V��?�;����\�-+c�<LA�A�.l�G���t�h�*_���7U���������l���
,�s�U����Ԓ��B-=6���Jl�[YզvT������Z���2���Rhw� ����t���h���J)D���,yn~H�q��0��-�����aQ`l��_LF����e�5t����40A�����yRT`M�;/�AUy^�#������[S�7��ʬ[J�m���`XZ����5��ݭe��^���I�:n̬�Ƌ
�n�pŮ��/I�|O�=�je��y�u��h����F<�j��~��{��[o�����{��$@���aH6�2�``�9,��Pj��/})��b_�D`��q�@q��*�r%m���cb&3�|[hjU���f��%�2�A�/9��R�\�s�e$�^j���9��R+���ᦦͥv���D����\PH��=}f�>��v�B���`�0ۤEo�cK�����s7NH�+��쮫�摑�qa�M�a������ʬ�~=��4�̔ ��4�I_�g]��e��@m!��N�Ő�BVck�<�0��T��K�ɣ�DgI��H�;��L�k�V	T:bU�'qQ����IĿJvn�)���L��Vh|K�7�]��X!���<���:Y���:�ŴВO���)~����>�Sc�O#�NXc���5i(=���\;��-h4���`��m�T3A{|��"?~�&p�p�h�W9zY2,3_sc�Re�d���p+K�8q�܏���:��~�#�^���G�b"�g�v)([v�i���H)���Re/㔲W��̑";Z �_;��ôp#-Un�:�l����o��D:.~���E�I���˅t�$�-޴Y���/4"A��P��������w=��{��	�����Q���r+��jYE�?SO��E(�*B��K)�4HY���*׈��6�QȻ IP�Հk��}��V⊜y��\H;:��6<�&Bv!�OZ� `�L��&�.�AI�h6�w]��ř
B`�"Y�gr�0�r!� �	b��:���Բ�"�.u�$��w�j�F�t(6N��O��/s�OHn��<�C��t����Z?�N[W/���ЭU�D�m���`P͂v"��k�zR���LKi��� "�/X�^=M�@d���;���e��y��\D�C5>�<Mк+j���T��9�AG _������}�0�C�	Q��L=�@Z�[-���̇9����j�rE�7e:*�:�&�\I ��]J�,�/A��kDSiJ�<m�.h��s����ο�'呼aP]Nk�At�����)D�E��s�7���G�թgn�ʟMkiuFS�cW�{�`�*< �"�2��<�6_��)	f��:)a�k�v�BZV�*H1�A �v�mm_o�?�h�%�|�� �cf�>YpSH�!¼�w���>By����լ��z@�L��+�ye�*1�+I,����]Ⱥ���	����-�v�,k�'p�����۴k� ��t�@�O\�x눭�C��J���������>m���SMx��I��:�$&�����
���^�K�v��,Wd5����ڦFd\j�k��R}!�Ю�d�L�s�]�Q�̸s�|�a�(5*�H4����(���-��9��`xs�>q��@H3=�	9M�~S�mw��,��8ܛQ1R�/�w����{T��1��A"�3%F�X�J���NA�u���E2��pp�v;}�J��+mxx����)H�Vd�ϑU?(���$��̐	{KPc��L�Y9��dJ~j����D��S�N��rвJ$-'�醠�|2��G�Tn�Z�y#߻��A�[�ﰬc!"�J��f"��q����hvf��2�gs����z�|��(��	b�����ڣ��(!&&5�s�<W��j&�D@������ ,}4%�ã��������ѢrƖ��D��h�$�=�����@>aǪY	Zݴ�7��J!�������̈́@@[�h��n�%��V�����y�Ii�Z[�d��y��-�s���Ĺ	vw �wA�*H�����������v��:X��h{A��M[�H�Ԯ�&K��B8�]��Y��/F[aO�f����~<�@/Ka6��֐�,X/^��G^}�>��K,d{���/�;����/~�o�%D��ژX�|-����~��������X8w!lLkIw ��\6�^~7���p�/<��_�������g�l�E�b�,0[�6�;U�s^�i�9�u>��~�~��>)���W��
&��g��y�t�ʕ���o~[��p4օ��������k�&d�����ݤ�;,,�B�s��-id"`5�`�d���н��A'���wx�%��?>LNm'�h��l��h}�<]�~�>z��y"��q� O��!2!�&{�&<:����&",&���u��İA:���M��������O��u��ɔ�)���5�_cu�╖���=��_bs�X�l�0���l���� ݵ�Y�̞��)�V"㝉�Q���
����.'~^��NƔ1�т�1�,Z�x�L;�h�~.��c�U���E���P�JZ�&�c�.����Q�m���8h�h�9��y�6i�z�J,�8'�P�3X����R��Kq�蜗ń�O���@*�kk!���A�y������k�֚�h��<�#���3���F��ٞ�g:�Ӣ���i)�:�� y�`3u{���^���7���4�����'?~��рNX0ܺ��~t�=9�;�]
�vh�� y^ӽ�v�����I7��(��M�g��3'���d��.��Ȅ776�h��F���,�6c�	����EX���&�d��h��/ɂ����]z��o*Bc����A7�� �������1�o��o�������:�k��"geD+>���Z���J5��l��/]�D��뿡���_�roFJE(D7�!�A���� ?�Ҧ����K����O�o~���PZ��^�%�xΝ��/�ǃ�d����d@����}�o��5׀-PzP�jZ���h��_�}�g~��<�`+������R������	��*��
�v�Ok+�����O�����E�	��F���~��3��s?�s���}N:4r��VH�Li̤�E�h������'�����ʡ�n|��T�l�aHJ˭���
�w���Ѕk�������p�Hr�.?��Y%���p@?|��������D����A�,�5�ϋ���?�Z[�	X]E�����?[�bi��V{��|g�������+O(#Tn,w�2��Q�����������_�,�x�G�؆U,ܸƑ�u����xD?|��E�$�)g��T��L�t"Bd"dɐ\X?�Q�9u�� �����M[~tz=ZC0���'��t4�6:�=O���>���;��[����}2���t�'��F7_���"h��L����D!����bǄOQ��_<'��g^�I�L�'��XI���G�sh�t)�A(��j�������!]�|�ַ7e��R���0JW��M'��$�t
mA�������B���`Zj�L���.lӕ�)c�&��w�̑H �H�%/rCÅq2��ҟUh�B��甅���F�^{�%j]��(ঠ�:�����'��F�v+��=���?�՗�+�u�\����G��4Ĕ�/���]ߦ���M�����l�&�����n�%��MUSAy��c�<}���"����L��1�>�	���/����Ư�c�,Y���ĳ y�����sTM&������M_�җ������k=��<��_@���ӟ�(����j��I��`�l�iT^!G�PY�������������ߕ'nY���aW"��Ȣ������?��u������oUzJ�W";��o�B_������ޓ�����&q�H��R,����/]����/h���5F��pD7�4S�ш����У���ѓl���p�������ǵ��CĞ���0O����Kk�{m�k��2ʷ�ָ`�9���G����mM$���`O܁8�����jm�t����]�񢠎�� ,��)]8��qӱ�)Oo
u��?H��u�0��ms� O�-L�0~k��7�6簙Qb�T��\��ʡ�)#G�t���Ç�.����>]�z�ֶ��'���N��(`B������6����"ؔ�:>�7(5�x����ӓ��^꯭Q1'Y�!�h3���t��+����߼�.���rnAhQ�Yu&�0�y�n}�>��i�Y�};��<-R�Q�V4eU�":�B�Ί �}F��^�Q�
[xiY���_k���#VP���/�kluuV�1�Q���ҹ�lKǌ�4>�8�	��'����֭��A��˺E�����<�=�ş����Gh�f�	+�J��h3��enQV�'s䤯�U2��2��Nf�U���@ pt|H������E:8:�����ȫ.�X�P�8�V[����`��fS�bp�3f�H�: ��2>�'�n3��P�'����tN�b6��O��"��|��wS9+�T+7w��4�(ϋh[�W����<���}�xn�Хxb��đŠ�b4{(1�u�O���
�O�q� ���R$ks�Ε�s��%eC)sTLA��aӀ5n�EQ��X	2M����N��e�_=�J�Y�v�6y�y�vxһ+krS�ߣ{��Z�%�$��i�R4���ޖ���G}-� |<1��nSӞ�@1��H�Sm|iNh��>�,�:�q(���7��w݊#EҾY�� �JD�O�� �?��G�_�A?�����f���6�i	�=J��?���z���
#�c�7 ˌ"*�rgV1����n��O�����|�g�j��X��f��ق=T�)�F�� 4!|��w�����A�kt
6�2(�+F����;����_�%�t�0�ͤ��D���!-��\�h����D���_�=�͉(��T�阀���*5# ]Y鱀�g��6���q'��pKȽdh�O$A+E<�H��yrȟj�%f��9Z��bHڶH���(��t�����+���v���Y���B׷.&APr<�6��}����DR(F�Ri���С����w���i��~����ٻ�:��jP�����'��f����/�J ���w��mo�"�y��HA�n�>_�Y��gFĮ�8S�,=i{c���?'
�p0�.��AЭ��X�s}����ʸ�T����%���,���&�-�xn��ʾ����!��\0�{��t��Rd2pY|��sey�pM�|�o-<k��A��o���18�:��2���g>E���Ͽ�����mu酗�Є��Ν�Z��u�q���k��Q��!7/�m%I��xP'`�u���Lx�KJ�j����1��-X�q��ε,oR�Z0�K��J�������U����,��sm{c�n߹E���DY=z�X^��Q0�N������FO��͗^���Tq���<��,h��e�'��uE���;{���1�$��lndT����Z�P���)����W?Jo��]:�s�ϑŒE����(�U�z����2�n#d�ɍh8��|���|\���f?�0<�O}�t��ޘ��3��%�ֹ�ri����;��ߢ�������ӘZ�ϱt.m����X2lڭU�����ؒ��[b��>���Y)�qFv���w幠Yc.-�3u�ZA�9�fE&~�i0.X�}���k���7���yW*-��a(^�v�/�Pܾ�sYJz������bd|��Mlt��76��u��S4z��Ѕ ���_�{|H�>���M���w����_Y�ѐ�1*� ry�5�!m���o����w�|���?|Y�����^���sA�w0����ۥ�	�hF�G'"�s�c}*�ѕK����ߠ���7�����%��;�м�5��9e3Mi��Ǥ�	��um�je�T03�Bz�æ�^<�����f���%ɡ��/|����o�΋a��p��Y�uh{k�'g(�RJUkJ�8��+�ڙ�:"��Y&����bm��<UΚ�~���"�U�W�l�h,^��2�נ2���b�V� s٢�I����ի�3?�	���ܷH_��vӌZ�����H� $���X�ۄ�O����dwW��.o���2eB�j
��wJ�)G������+�Օ6�~�(T�r=��n��Y2?��р��Xk#b�XX17�����C�J[zȢ)o,d^ �P�,�Ӗ[s�|ª�*a�l:���_Y�����FҰ0�{�I��D�4	C��i�㚈���Yy����t��ҭn��V�Ǡm"�����"%��-�6)؂0ș1�� SH]b! =L��\;�{��{@VDY�H�[�J�HWK׶�Y��W�C2���Jm��ۮ�bUb�a��|<�c��;!����-[C	Zͪ,���ed8�J'@,_��X�4�B���X�ZQ���]�����o�s��
~\�OAP�QJN(�y����O�,=~�K_�����+����m��1�&�M�k�Z�8���A������׀{@8y�N���������1з�z�'e�p|���
��zr��Pv����b��k�[���I�;"���$v�j���oŢ����7�7P-�7=�EK�P$�]$��U��x����.�������5XR�({`BBM�U"��J#�S��2X��F� ��@�9ҋ��K%�y$���K/Q��%7��Ps�A��tʦZ�]�Uz�wHm�*<�Z���F��E�6T��"���cj�Whuc[ƙ��B�)�*��}fY@�NX����֝{ԻpY{9寖��+��i�G!�M��=g,�;����#���Őe�[
V[�q���-Bw���+�2�2D���s,5�V}� B&c��3$�-3N�@����ڡ���H��� ��-�D�4 J���{1ӎ��u#}x����Ǌ3��Heૌ�Q]H�u�B�:+lq�G�؀�A3s�W�5�>�JJȦ4�>��_ni���H��۽
힌wL�e#Za@&�e�dR�FZl!"P!c ����;�'�˻8�&�|/�<h�����k����*�
��S�"ISʰ~�*��w��?�^g�Y恼�8�b�F
���&K��3(ۏ&�'� r�T�"Q��S�2��O�6�b�UZ�#-�+�5b����?��M��jO�j�U�����Q��$AA�R�iے{��E�˦�+'6("����Xe�2Y4Sk���
�`j���*,d���ltE��ܐ�UcqŸa��Y6e3Zl���/�D��e*xm�i��Ql�F������D����8�;�����x���O�_K��E��;�"��|�X���)O�$A����eSuumCHɇ�P�FT�e=zr4��{[0�O.�oZ�DR���4U�S��,��$����z� �Ye<�p�r��v�p]�8OEw��~�6u���:��嗨�D�%!�,C�s6jT}$�uV���E�� .P&ʽ',�Ɉ�A�u���I뗯��`Fw��	����$Y8	�����$H�6�*���ZBŚ�	����<p��.UN��n�	?�ۏ��:'2l�Y6��P�U"�Kك�����rk��� t#��Ǌ.��n�ʩ����u6����!e������Q��B\#(J��uk�(�E�[_g̲T`�V���t���kvek�>x��wL���ڶ�p�����q����*+g%Xd:�4L����6V������+/й�����G����,W3���+i4K��z0k��ɘW0��b�Qۿ(t������6ꥫ��j�	ڐ�kV�d�81���J���:mk�,)+�TTa���8��+_���G�t�5�O���V,����Ā �޾����בW���j�bŜ+4�GnIα������$�-����y{6'd=��-���#�&Gӵ���T{�E@Mƞ��_��Fm�*���X�i����=,|������}muE������Ts ��h������pNl,�M47^x���У�c�mY���>�OvĪ���z豙�Qv
a���N��	Bx����J�%�2H�K/� ��%b�
�~�?x�=A��!��f��08@?Y5�M���`��h,����,�7��ᱴ�G�j��}p��e���4(�8�<>���[U�X�e���z��+A�=��-�	F�2����c����y��HL,�_(s�Z��0CKI|�d�f<�CF��i�7a�`A��$�����9�������'�Ǟ�3 jK�j�.\��{�X�D�����pw���y��r�~K�a�ć+>gMND�J��퓇<����K���T�S�H�Y�Ӄ�C�9Č�"��tK�����8�,AO�2Ӽ]χ�ۧ��σʟ�ʥ
��m1rfpƿ���V`-t{�l����)Dqa��mx�	&;�|VZ�3+����P�m�Lk�cmX��_v�"]�L،@=�uʎKA�S�hn§4v��M��׿Q0�~�#��W4���!���k��<x ���7��ӓ�]Ax����E��G�N�FN=)Z�c��S�l��ߤ��<����a��I�����V��*���
"S�ZlG��Yi�)���d��9ߕ���(<�?��?�|T�$�!"܊B�#@q1K*���-�v㺤;� ��r���#��"y�_��Wt�3E?]�yy��_�_�N$��`<��I� t�;g��TY������ث�I~/�ğ4���W>J��ݧ�?��oO2$x˰e�����^�{��w����3���drlU��e���Wip�ϊ�#�|~}m�}h�+j�y�p��ؐW�p� $����`��,�l�R��E�.�q���K�DIa���E޾}GKrlda��1�VZ��kC^p%�G3q��\z�9a�by���trG�n����[<�~����	�_���{Dּ��y^�`��{؁�CbU�Y�����ߏ����&M�}��jք�E�/`��0 �X�C�G0�e��������:�(�FP��ҕ��B�"RmAx��>ޡ'_���+`qa-b���mYd�d8��ۓl'�_��������H�lt���R!��n����%�b[]3}���<7UL�R�HE@�t�"V8 ���� �k�.ȷ�v(�8�:�wx�[����8eUP(KSG��L�[vMXYMZ\=M����i�w�
����w-P$0qd���R�-e�.�ԲX5�������ohb�RL��lT�?�&9A@q:�� J�[Zu�Wz�R��4�<O��{��V�����WDp��y�����Ţ����3�����x�#���e���`Y�F��#xV��_`��	+�cT�LGR	�����?��?/(���H�Y���-�_e�_��LZ�W���Wv/��P������m:���o7�ȼ��C��Ch��H4��M�ω�H�	^�:5�B$D�_n AlSz�c�{��޿u[KC�9c;����R�S����5{�HK��4	�,��|V&@έ��:4"�vN�X ݹ�H���?ٓ=�|V(ʕnO����2��i�����k��)mT��:*Z��Vum��_�L���mQڒ���)�O����~�L���M�8�㩸W���m,[����6Eɠ��Ռ�=u�����}V^*P��B^v:-��UW����PY��/���Y�������U�����	�S�S�q�cM=�m� lK>�F^�\1q0w��Ӳ�G�WO��٣<A/�fajj���Ap�T�����-7d<Uͅ*yr J�ŋ�,�Y�$_��gW�Sm�L��ɹT�UT��tA��)�.���P!FSe(�3���	��k` �iS�;Ll��}F�[�k��h큲l_:�J;Еѱ��%����yԪ��(Ţ�7V)(���HQ����Vn;����ʠE�}�k�p��>��,r[a�WXHwx�O'#e]���^wYxN�������]gA�����My��`4�1(GishQn
!.f: �"  �*
bfc�fV� �"A
�WP�%$(B��VB	s�נ���_V�6��\������ofUr�g��N5~�y��oHm<<��6�	A9��DQ�7\<�����)�k����\}Y.A�kj�51�i�@�Nr��rN(�iA��B<Ȟ��yLb��Ab,KL���tG%��x� R	�C�	3�?���H�;@�_�q�\��tW\� ��ϋg)q#�S�D�3^W����������L]�Y���y�^�-G�Y����!�Dn�~)�z���p�fe��΅U�b�� ��D�����~��x@��c�8��4�S���Tt�J`m���j��k����J�Cq�g��3�Ct�.=�_(����9��!ޘy��T[DT�����sZ8���KP���3��WyN�кBt�s�+��P"���:�'�C!��l�I��H~�g��O]["���aL(��s�v[�¨m��Rk��V��L� g$��RFP�jv��@ݥ�G�51<s�6�	�%��6�ws�O�����tn��x�K�Nix�
 �@���\$� �㣁����l�����%/.)7�����3���M�Z�����P��j�&�#��0��a���p,e�EeI�梯2�]et	T� �:�.ȟ�3b��l��X܃�4�>�}�vF�U����$��O0��ZSi�2B�4�|�)P!hs�4�^�[��o����6�g��k~;i�^�j6�tM�T��n'
��x y�UҠO�Z��⚳�zQ\#��N�
 �󣓳�C�u=K���v���j�zE�89ָQ�ov��q/P*u�,�qPJwd.��b��)��%r��
&�2J�\I0"�SQ(��o�!��B��h
��d�4>>�"�6���t���*�zh�{�LS����-©�	^b����И��o�����9� ��l,����/}��]���F����I���J�6Y�@�n0�[g�h�R�*�|emC\�̝p�E��ߗT�A��πo����w�zH����V�a���u����� 2�
\�V��FzH<�ED�?-�������:d"�=��js��]Y3@��+����+}��7"�LU�\�_+��PS�z���;dA7F(���9�;��la)R��y�=����Mˍ?��{ěAr�"��KĞ7-h�H���?>�<V:��,�#$mL,6��q�P�d����˫�'�^&$�"ؑ�@"�R���R�N��L+��<��ĵ��+�B���h0�٘A
��r<U�5wG�H�t��F�Z3)�!��ϙ�۵I�%g�f�=z�(��$�6fT~(�* �	�T�|���"i����(�$厪zh+tX8�q1��ᱵ�M��x�-l	��G(�A>�x�]�!�C%s�J��B0P49MZ��"����-�P�>'�/A��	J7v����r���ښ �><A^�I�A.�	i̮�vu�6���C����2H8�E��{�PU�(:����bJy~�hv���8�tyS6�����φ�ە�.���%)Ǭ�S�,O��ݾT�=�q��V�\5�l�~�DQ�@���_���TB	����	\Y�9�Y�77����-t��v�⁏�w�?D���h2�M� ��ޮ�R����Bg
G�`���w�+s
�+H��r��Zg��������05�%�u�� NX������m��@���wh��(�}PN�,��+���@4������u�4�	����<~H����� ��u�?0R�2�n�A4����q?���z|�#~\���
�o��%�T��}�|���%�=O �̊��[e�G��uY����GOb B���t����w��=���\.��m	�[A�۵x���AP��J��Ahu�����vP|�\�oݲ��X�Y�X�<|�B.��
��s�[b���SH.�ڤ7��Rڴn+�k4�5���#Q�P@��9�f7����	�/�A���n��WQ�$�"�W�ց�3��\��3���Db7Z�����i&�r���C(@a}a
	A[K�u6����YK�|&������@p�t�����D�p[����J���HZb�T�X��h�jZ{h-���ҙ�K����gCy�fpW
Vm��]>���6Y�\�|UM<x��U��YG,Pwy�`����7������t�����o���G`� ��#ͽ�0��L���L\�v��Z|Y�����"�Q����|�E&���������j�l���\���.Tn�_"��o���ݧ�	䕚шvO���� �%��s��~+��Čg������tt2�T.�-����M�n�fo���@j�+���%�6�i��2	Tj9��ގf��(��
c�@��y�HkC
�L/�@@�l1������@�},k8�Es4I�f�mk�$����fZI(����`p,� 9�=�#��� �����1+	)Bԯh�7���ɋ��>�Ϭ�AMiGx @�C������Ni
V�6]�pA�4�,��	�[�Zrn���QP�u���\��=-WRv�ca��& Y�e%[$z��e!G�w���oD�w�э��94EE����t��Q���;�ԝ������$Z�JxOϤ"S������^���=)?����N|��%��<�5YC��{(���:9�K��<PU��@��!C���]���/���m��� (��L�}\�`�
z8f�����p�.2���\���m�`�Hp�EhI%��f��T�#��(����f�8�5��h����1w�TAP���l��������4W�na�'km}Et>7��#Nm���H�'�/4�^����@O���k�'q9����f��%"�H ����WJ�#��S@��B�Q9%]5ە�����N�R����K��r
	 u����U�\�H��y��j��ح�9�N�qws��T�K�e��N����	hBLC���)��A�5�π�!��2FQ�D|�� ![iR|$��*�.ˌO��x����*KUau�x7ȗ���	���iG�R%"�}r|b�!QL8dm�u�֖��m��:��|�ے���ն���	�H�e��'�dwOy�-h����hY�AK��g�$<�P� �F���h_,>"M�t����)���W����r�p� %>^��w]Da_?���?��[��
��p^��\�ueOIg�c��߽wO�-q�+�Ha\�i*��O�g��$�_�|��2�F&K�L���Vd�� �'���9��6܃�1`p'��o���&�BZ��wp(�������5���r1$�Gi�$y��ۼ�T|��-���3����,���"=���(�C�H��Dh��dM?.�R�"~�L��  ٽ0�Ͱ��*�
FLz��+�.�qB���y����<�U^�[ۛR�{ tf��d���U3	��,4*P�!��<�Vw{���o3w$��YQR��l�k=�ў=���/]�IHǝCa߇i�wr�P�Yb,�^}VB*܃0Amlm�� ����
!
���!$��]�6�"��*������ں���?A�@	�
���+�� xSTb� �aj:l�����d���8'��&��@Vt�k��� d�P��\e�o�����@�ީ���u��0˃5������ �7�y��O���3���vߡI�%�8���B�T;�\��#����)Eg��H��s�$[�-����YaETщ \k1�� CU�p�"�~<�ʳ�>��M�XQ�Ӯ��[� _JЙ����^��at�4��X� :���l���({g+��ɚ��*��՗n�}F��+�2�Y'�5�D1����%�f�rGw����*�J�\Xc��A�[ݤ�˗�� ���L��bр��;W�v����r�:�f��9㥬 Y��������<��խT�3M3A0����Ƴa��M�gV��n�X�c�;�<���h�J��Hqб6�s���{��X�f�{��ز
	hf�l���X���,`���s���!x�&r�Ȼlb��2ϗ	�扅�6��Hh�X[A��.C�y��{�Cr���"�B5��g���K/��w2A�Ǔ���\-p�#�C�MF��}^�G'#33K�E��x��E���O����/ރ�hRo������^[<_�#:B�+���k��֍�К��$�[Z~��M�r�J���B�K+�LSP���fg^���D���y�������V?H�&u���:y@eLm���g H���hW��T�v4�E2 �5$*������t�P�9#m��C�[��}����>C+�AY����Q�kd �S ^(�/?Q't�p�?�;B�< x5U��kE�[Y�<m��y�Z�{{�㗼UV�ₙ��k�5��퇇'���EA��d���s�hR�(����֖<���>��YN�q��
�% TҘ�����Z)j-���e!8SZ����ec}C��^��ñ �؅tA�3p$������� ^]���x���Ub[��0�p��TU��M.GRo��{�p��@V�l����
`>4�͛d_2� �+9��B�ϒ�rbS��Ȼ��A`�+�M��@��ZYQ�6<���!�8��6�����Я~�W��oҟ��_З��5��Y�h$cv��lY���L�j�4��^p/�/8�iY���˝]�5N�?�EP����겄]�:���N��'RH�g#�43�IZM��Z�ylUy�s�ʜi Sxc-�mm�����R�z$K�3�}��a18��4��H�%k�(�sn[�A9т���Ee����Y�n���6��+��q7�����	@iԃ��_�q��Fek����(���4�cb��d&��F��j�Fay�x���;q�@�H�5rf�ė�'Bb�si}�F������<�L�$,��Ԭ!�ja���#�N���1�I�h�i����KI���C��+T��y�.���A�e	���,�
k�M��Ժ(�R�p��K�+���������u��Cf����w��)�t��=�$Xu�P?-�<�T�I�q����ѱ���G�R���y������7�l�������xs��T��&>X���(���{ ��k�|1ݜ�;b�!�������i
A��A��1��>!u��F�9rAW�hߊh���=أ������%���2]EW��U�Aۖ:'�`��4]!�C��?�
��ų\��gDw�G�f�T�B��M]
�@�O�%h�Ģ�8γ�?������nF�h$c�멛�孰I<��i"�V��|�y�e���3e�ޗ~ފ\2� >R|Ϋ���͛�F��n��l�%� H��qZh?&��%}�'�$bF�jB�����~:o�f�������G��Iu"�?��]k�2�����F���G��ik�������RZB�f������1vb�o��f֮%�zϹ�p*I�+��<yQi�T9_,�K�/k��U$�	R���,�"?ҵ��D���{*�u�%�ٹ@6e�V���@�,_UU�بg�^�"x^� J��UL��=����ңU�!-kW�v�5���#�`|�2I�.`�*��d���J��J�V��3�5�>�X�A$8�_ަ./�"���QHvF.+�/���ڊ"< t�$�)��A��vA-4}��vXU��1a����Y(����/R�Ёu=�}�ΟۖM	����6��x�j�L�2�%���s�E`���zd�陎��B�k�����@!	���	x�vh�եK/��o��.�O�Jrcd0u���43�"'*Ž������T�؎����S,���M�ڧCY���(*�`�ݦ2�7�T�̷[h��J��!�hDI�:���TFy����f��+��[��<$xdi:i���/���dV�#h_l�8
	E(�0H������~G�(\������0!��8���1�〢p_��Jė��s_+��AU-d:���ߕ�I����^��
X�)!�����%�?Υ_ó����
��^\x�2�M���P��"�-9#�uMp\b�0$��>_���{)/��5R.��uJ�>�s�M����6��O���!���
Y����*u!����O�l��5a��w�Mb&�8�0��l�3I7���=�g��G�V��M�&@�	(=�p��E!���ʲ���=�VN�!������OZ���<|H����V�~㆖��d���^���I,�'��n>�R�`Z`�'hT1g~���<Z��߱p�ic�?�(�n��@����Q�m,�q���3i�c)���{/�k@�VQٌ�� Ӳc\m�K\,�X�)���Y���%7/�]r��Bm�(du�x ~xi�|�:�͑���m�����!;�$�c���R�Bz��suu
D�JW��Jc
�����%�ꙴB�U>�2ZC0A��2p. ���V�5[����ƧF#����g7�|V��r?�r�nkd��#�-5�����e�%�?���5~��h���H`��w7���cT���a�G�tT�J�w���!k-��J�n��d�K��d�C���� ����� � �`
	�"�y��B���R�����A]�>di<@���&>�6�jg s���Z���\��,�	< �,e�
Zu#��y*���OW���*QmR3*O�\r�A��Q0������Fz�����/�s��}Yj��M�R�Պ�(����Ӊ�3��!�Y�t��u���ģ-J���I�{P���b>�0Sd��!�r�db+�N�n"Ϫ�a2�}fNѲx�\��L�h��U��`ͦ/�-6w>f5߯Ͻ�552��&�62����aѯ�B����\�Y0S�JD����Z_K��畮��A�Z��&�$ч�\�M2G$H#B�$܃�ㅶ��S����U4b�O�>����E��LD��{����Ayv��Lf~���3�+���H2z�&�(�DR~���F�;.%��F+$2���ʫh��7V�,���m�z9i�f�f�}AR���E�W�J��=�&��/�Kh��l�����}��؈�������#��W�O��2^�P�W\F!����������!D؅V���mM�n��4���s��}����	�M\W���5������ye�EP#�@�B:c+��.�[��-���Æ���-�'�`*����^*dI��cU.$,�A����_���j�1'LCI�3?h�%� KN����~����K��������G���岢��h#Ѳ�F&�V/^�� ~��#9�`鰦h���k�a�|�C+�~:�L�:Z�������:I�h I�'y�.z���m��*	tU�̵Ր~�;��%s����K�g��r�l\ �<�&N���X#��,���Yk&�h��c��v���飰��i{�^&$"cK�I���t_m����c�3�a�շ;53XS�օ9�8�>&����W[R�{����8G^���t<�Z5��d�uv�������'X D}��1o,�Ļ kr3�O�`U!8��2n���J�wQ�
3�D1�_Nѩ�ʚ Ư�tN�D��xsq��g! ���~j9��^��D��?r�!��|�Y��/�Vʱ-_+ ԟ���P2�,��8/q����LX���ҵ+��B�'�,t��T߈ϓʗ2�Wx��g��T-��!s���|;ᒌ�����[��y��9�����ѿ�ҟ�����P��k	��
ü׺~gA�iZm3 䖡%�k�������jU5��>56}��I*kk��IH?Fh��a�C �\J��F�I�-jM�u(g"Tѿ��o���ڦ|FZQ'�X���{Ukçi�j��%׉��Zȇ����U��`�p��VY�
��V���i:[Z'N���Rg73
)��b{ͅK0BʕȀ2��l��v4-&CZ���Uz�ïҫ/�J�|���uA����D���݃t&�甙o2z �*��J�[e)]v�	�������4*d3�P�؎F���V|���<��3�����;�zYDX��˅t��*)�D�eA|�(.��N��O����!���Ƚ���6��
p	�:�7$�y��x7�ck%d��z�C%��i��{�LG����Q|����u�m�]�7��"�>�K�	YT��cV�[�N��q���kn)Q���7i녛͖��:�Eɗ��͓��ӎ�(9��ه�N.�h��g���f24lf�xG��!��7R6vLz�(\|�#�C�0Ļ��mj�u��Z��H�x2!��xT[�ۛ��y۲
�yd��#��}�5WϴBXtf��v��ң�p�:��m��85�S{�4/�|��*�DһK�T��y�cC����M��t�7��>�Q��_�u���Wy���i��%���3�,`V����yJ7���L��r˄jw��<o�x &
���0���	�k���PGV�@Tc��d���3���7�%e���
E�������μ�E$�n���Y���|�n�8��_��Y*��"����{K��/��>H��
J^�Z^!o.�T��2í����+U��5"��0g��"���T�z�JO�|����B6F3G$�K��K���Jl�9�I�ђ�iP�6~���FA0�S�Jޫ&��Z&)F�m���,3M�ӡ��.��$U1��A1�r�(ٮ����M��S�.Ni^H�O�M�x�כ���٥��7h<��|&I:gː���r��>s����T��!�T��`BV��Em�ySd�T�CL���֛�����Zi���W���W�������c�}Jڃz�UTw�%]S�\�j�eVE�F���t*�XY܈e�U,�q?���t��I��1w�~	~�!�3��m����@�"�Z�*�՟���2�D�_(��X@�3�T�"��?e��Os{wR�`k��r`���N�uc��-Xf>4�m�Z�����+�ek7L�>3t�k����N�ѝUͻ��Za�{ǟ�e'����@��YY��:�c-[[��,XHfu�n�]`�^oBMpo����\)|sKK
�K](�OJzn��Gm���cf�|Ǭ1���8z�FV���0���˸25=�\��F��Y�����(�.��!ű����F���wG�τL����Sl��-�p�{�T�3��L,/4_�ϫWƔ���s.Cj픞�e7�K2Qn�*Gp�x�1�k�b������F�Qi�ɏ~�>��O���EP��s�u}��ZP�;�h>U]�9�-y�s+)��T��sU�,^��;�ʗ����ρNYF��-�^zds�欨�꣒�I�LR�Ƙe�zf��-� )�"˟1�/�t��^>&�}M�9����3��M�B8�U����b�z��~��%��yZ��G�#� CB�R/���AU��2��H�N����V�4�y�$��5�
��Fy&����!�k���T2�)���e��E�c�$
j��e��ZM���µZ�'W$Dt�.�e�6A�Q�}4r"@��Zոӟ����+ ��8����Xb��f��v�h�2��ƣ��������W?N[��T"d�����T@R����#�}`~��s�e�'�n���;c�!Ĺ�}~]4�3��%�s���_]���%��Y��X�q,�#y�Yרh���ҷ,w㥐��
�؟��B�!s�Q��T�3E���m̂:�S'x��!x�t�\B��An2k�v�ۃ��I�e��B�m(�<�bCX�@h��l�m�N���\�@��,%~<���h6^���@s���t��P#57a��<������в#�TU�A��>�)w�J�$Jwh����/��y	�b&�BH�ڷ7�Sb�#.��U
C�<����(i�k�q��Z��9|@�����g���x���.�iC{��s�߹���8aE�5�8�l^��o2Y�t�a� ���z˜�Ҍl��3A,�c�_m����͓�S�7��-�[Zz����{�\�ڿI)
L��j�!B#�(��_����/�A���ܚ�'U,��vYYB9:0���o|��&�|�
�AU���Q�BӅ�����h(g oF?��� �I��sM5���b%��eGj����{en�Z৲�h��'-A��g�
��_��kst�ƮS�̟d��֞��cVH���/˜�g�	�o"w��x+�<s�ln�S��X�|���8��|4��y_wh��~e�5�/]��!hr�Ui>��-;��Dw��+��Jx��"&�^&Y:�xo�W������I��Y��-;����iR�i]��\���T�@�N�Yqm-�JS87���V� �?}P�C�Z��������!M������t��N|�Z�a{�`Z��Ա�d�~�$��®e}{����/aq�i^j�Q )٦���8�j5!��ZPp"���.(����ڕ�W͖t�vE��t�(8Ψv��'z�2��#ờ�#�UK45��'�i��������g�j"��t^��Ĩ �-_eű̕e@I�1A�+�H�2��Ƀ'ː�G}|�v�jA3T�&^��o�t]���Y��x�H�hF�.��p��%>I
T-�P.?S�ȅ�L�9-�Dq�E��*��\����c����<��:?�4�����u���J����ȟY�FY�|��}�z]{�,Uz�~_e�i;�WO�l=�����&�}��!,;O}��z�{�Ϫ~K��~U���yi�����Au��ʳ����ekӭ(�o����TF�U��D���	ǖx��.�����@��i]�a1�4�˻a���Z�M]^�F�.y��Q�A1��r,�1p~��Hҝ�LٙH�qe7_�h�囼��B��y��o��t8�^/�q6�<6B�F��Ah}�^��UDE[]���{�#�n/I�6�#�~[3�V)h����#�*�H��lA]��\�X�th�����Ή����MY�QSr�[��]O=���O|4��)(���(d�}�"�3�I�@E�թ����jͺ*��Gd��ֈd��.|+G�K��~N�yj����BT�t3�D��%8��Xv���֩a����+�Sh)H��l^�>�
��͟c���t?��E!kB2�-��?�K~O B�?ҩ�x��6��e���		AL?�&���]�7���b
���e郚��]�#ʿ���B�'�m;@Y�R�w3SR_
�e!��h<毡�S�Y��d�|1kP�,�%�9��9>�&����4��~>�~P��š�������j�&�C�h�աrwѦo&���II{{#Q 9o��V�>�ᗤ�����?<��1P�
~�y��LE։Օ�B�Q[Y�$TAe�yϹ�葸��Fسϻ�~�χ�h���dVÔ����zP����H��w(������D��3
<ر�)k
�R}��ް���T�>�X����������ߧ����y�g	�=o@nq������K�z�V��?�l��g��Q/c#O�9
���nNj�}PQ�/
Zy�J�Kg��y�X����uF�[����&u�ܭ��.��a���v�k��txtLw<$����C�*W�vi�cf>��b�8wk�.���U��_����f;��Y@2 �Ƒ��Ñu�Jk�ʃ��1���EE�E���|���{������R��c���H����>uz-��<�Cp�ʯ�6ᩭ�����q���`���Y��0�{��ĢI���(��٧d��M�,21������!�0��-.�0G�7�f���c~Ju1����	��ݠM�f:F>y=�9��44���1��F�]!�`S��&��Ɖ�#p�k�%���< R7RSa�|�D�q��+d���1��z�1��i�3�'�I��ߋg|�,���e5�d!�f^*W��p3�jSʷF}>���q�#���.O�:�4+�����>��y��6��K7鵏|�n�x��66���|��ƁF���s��mE6:��x��V*��P?�I����@/���2F�m�ͨ����@�hO]�2�Ӊ��F�(��ҽZ"�Ŕ���h�?�ѓ#�ʃ�j��]g�7���x�M&3��V����O�� !��m��N��	�Ғ�5����J����h�:��E?b���}����~B����xҠ�ұjd^xU]vJ͍I��MW۩��y�g��u�K�d�ЩAȫg�@���ދ X�R΃>'t�*�t|���c[��Z�����[v���zz�U��秝s�[���� �~ޔ`��GD~������}.
���w�4Wl,"�l��V�F{v�}G�ud���Y��o���&m���ل�]ߺH�����g>�Kt��M�h����׾F;�����S��K7JxF�vA��ʍ�t��6]8��i@�!��;�����tx�\@��NY1zԃɾ���D]B����{ڭ6c���wY�-�ڐ���\���{��g�{Za��� ����`�]�s�}z�_( ���ҹ�usA��P�Fn>�N�����ږ��~���̧G�j���Ċ����g�"J�1�z����!<v�@���7��zZ�y��5Z��g��%�*T���M����(!��:WTč�L[��صߔ�v��T�y��-��_xos^��>��V�g��S�s�}�Z\T�����g�<�l?�ߧs���������dU��WU�;��͔j�,��}=Kx�P�� ��]����@c��D��"���.ѯ��L�~�U��-I�:�?�����з��-[�"�\MhX�&w�.����c�h����?�!���7�����	#�k�.���6ݹu����49.�c.Rń��� JK�hY�n���ˬۦ�jO;{�х�$�k1��Ϣ\^���)�}�����Mz�`�F�����du�C�j�_⍝�#�Qˎ>[��K�0���X��yͩjMs��ϔ���8u��V}9�=�� ��տ�}�0���H]Ⱥ���iZUypx+h����.��u�G�ηOZv��L��~�i�w��
i��Oo�I���Q#d��=�bZΜ�#���/Y��͏�7]N�	�Z�K�-6���>*Hۗ����+�}����ߦ�|�����@�{��94��҄���lD�M���M�&:G�ӹ�F 'tww�������W.҈��#�5*;=�t�U:޽O�d ���/]����[c�[���}�n��>����{,d�BD���X�cT?S�o���R���a!�y)͆�h�Ґ�i�Bb|��s�x�N�Gڰ�߻��--o@&A����Q����ʩ�זJ���!�������~����4~O���"��hq��"^8�]��z�8B���+q�<Ǳ�:Ü=[�2��$bn��,YM?����B����]'E�� n>���}=���<�=�rDƱ�|���i燀ul�pV����>�e�2E���=�4R��d�#Ɍ��L�"�Bu�O��k;J����m8�( "����DϦԝ����  ��IDAT��~��n]�sk�҅k���/~��׿E;�����U�v"��tZE���N�Ƈ��o��|��ƕktt|H��/у�wY���7��;y�l�l��ݼ|�>�3?G?�ۯ���;4ㇴ��M��C���>��O�?��������%��?���?���]��z{��]�AO�?�l|$��ED�Ƿ��t{}��~Wۓ)	�eF���L�hz=F�<WW�t��I��&�f����t,�z6b4�JgVj%���9ZA���]a����K6;<JfUb��yB�{����TyǓS2   ��\�����E&���b0Wљh�2�`Y��Ox �"&�j�z��4��<��J�f�.߸ʅ�B0�ae�@�)�M�%5�u� 0��i�u��ܫ�ǋVܜ���W�]o<��y)�t��"`��3���|�O�V��<�в��?�7|�}�}=��
�5������c�͞$����߹7���ڻ��;� H��d��,Zg�h�',9bb�~����?��0O�˄c<�41�%Y�dɖDY�(n�
"@�h4z���5�rϼ���}�{Ͻ��4 ����,tee�]���~��c0�d���e�8��ݬ���(���4�i!N��\N�VK�ણ����N=�����-����?�w_{��_�VGX�	�QH-�X�E[LwD�unagO�ŏ�ȏ�13��V_y�El��؍ڨ�q��y��3��"-��R��xУ?�j�7�^&���7>j���[8s�!���o��kaYŖv��Q�n��Ɛy�0Q.<\,G������bqa�҂�@V��P0�=�d�j�H
�:�DB+D�=�G�v���M�CXB�C,�P��S3U����@W�Y�q�4���^����A;-���M?�f����}j��sXc�A��!�)��nY��KO���`�[8:$H�k�/o�3��Y��8�y
4��\T�)
o���=���p�ܽ�7����[��w�����z??�{}��Nl{���{���=�˞���1�ÕK���}�K)Ú ���ǥ�;�"S~����8�j�\zt�ݿ�K�ԉ5����{=����zU�~4�%�����[!.�����z�X��js�"�O�y��&��p��9l�Y%6��v��!w(h�����V�cuٵ��8�X��;7P%p�	��1~��0*�G�M�8�ēB��@M�OFbJ@��'>����g��lݻ�*h�ƣP�`yiVz���������#M������dL�]i� �ΠE��;�K%Y��KD�C-��y��S}�Ϟc�Nk��aتV�~��8����"�hf�5Hm�:� �
\g���f�w�x/��^YzL5{�s�Qy��q���@�E�<��:[ NM	%f֔��Bn�z ��m�j+��i�\��HcU+���	�k�$�KP�P
�����v���yT�[¥*�}�|����޽5��l��[$p"z��4j������l��<� �T�����]8����AoЗ���m���-����plڦ�pa�P/����K��S.9a��>��!�`��_��_C+h����͸��`s���/,��Ňp��qܻu]����p,A�^itty��]�,@rdiy��o��vW���KI�j�bR���'���5q�L3T��H�l��A��L#y�2�Eg���j�IWdJ�w�턁-pĶ?�`��(�{湼�E����'�ֽ����pz]d����uҴ�y�D��~�́	��_l���;��y��A�����vW��]�&��v���UV�p-�E������}����f�]i�pܬ�\���l�"����Ε���:G*��krw�S'��'ǭ��I�J=X6�3i@�g���<~B�p\�F���	I&��;��HLw����F����
;�t{Cb���YIa�յ�8s�<�|�@��*�"m:b��d��͋�cn�����nK}�~<�.�#'"|��_��W���A�]Ā�i�3Do�-c#��-�L�dk吲2� �S�������>Bb⻃	������T�(Lr�	?HU���T�N�qeůo;��1q?{-��j�}nɚ�b&��Ї��`��˷1���׼�ebУ�M�CM�bf�L0^����� q�d���� GW®=���i,u/�}/��vν��u(qZ@�{�gr����\��:v����0�6����4�6�jkS��I�ok�e�ю�HFR`�	��0��!�Z��TKbP�7f%h�{��:=R�g$��w��d�q�_�{��=8���D�͍�z���L`j�r&�א(�f���K�5��\��K���v[My��=��W��f�Nk:��f�҈��@yw:Uģ]{,�⹆��/|�@���ł��n�R������˘#�\o,a�����[{�:�3�
1p%U��!��؀.�|�ӟf�66�i�f�nBYѽ�QIo��&��B���M�{@�;de�L���'�C�`���0B��1pu������o~����G
$�a��9�\j�_ &���86}��ݠL\{r�\�G�&A�u�u?a���[��0O�Q���5��u�`�ԍ�I�0Q>8��ҿ�;���z�Iͽv��^����2��d#b����o�"϶$"���h��+V�c�&�,��K���|gN���Vnv���~׮]O��*��Z-�����~�����x���Zմ�e#0�E�K`��＀O>�0�}S���X�9*~�)�$O�mm#��"ླ�������5Є��mw��?����JGN���_¨���	�Ll"G�Q�W��2���Fo��K�_IHmd���ir���#+��޺u��=���67F(f��%������;P`f��s8��=������;E�km��?�;|p:���6�Z�2$�K����Z6&���gƂ?�k�y��N��ߴ����c^p*���a��y�;��%Ȝ�`�g����0Ӝm���N����H@vd%����8�lC�����vY&l�K�1�:����k�n�#O�e�B)��C�ڤV������t:�N�Ql�ip���+hw�x�����KQ�c;q��Z��,�.Hv';���cL����Ġ�8J9ꍍG0M��8��X��-b��'pk�Tz�  �T���m	�
U�^]śo��"I�������w�:J�K��&$f��Q�8���`yn��mb�E��8�}�I��
��ئ��s�$��C��~���/eb�=ODS�"�8-wjоW����9��I���9ό�_Q<�A��u�1©�ymq�"�Mep¯�eKW��<�p-�����$�sO���>��暽�d��<�9�4֛���4�{�3NX��6�|��^כL�=Ȝ��	Ȏ��1�K�y*�j���Jn����jS?���)���ҭ����7%�T�8~���N���bl33%i����|���Jj)3ԅ�EI]�>���۫�r�V�����T�Ҵ���\+$6�����&��_|g��.��J��J�,E�Ŏ:hcs��[w�DL�;0B�Zp�7K�n�@���c���ξk�v�:N�XB���r� ,}k���u/6�@
�̠�zX��lo��iJ�l��4��`f���՗��;��*ǹ|����"nO����b�����2uRE ����;P�N���"�����"��r=��8��J֋�<�/�f'��Tzf�l��-�LR��1Q|Y��p�`!���޻�S����5k9JMb�����Q�ulkz��R�5��]IK��k2����-�8��ԡ�0�$H��}S9sg�v����S/����F�;�e��ܘ�������0�����?�3'N�k��LZ�Zڤ��\�	 yF~>�iH��صL2�F�5��b3��D��I)A)S�{��.9[M��2V��se�����l`�9�V:��dc�]k=ۘ2S��ۼv�t�a�oݸ���:��:.�:/�¶Y��Y`�$��Yߐ8V.XSo�a�@����kW�&5^�7����g�38s� l��S��Q��gp��[�m���1G�e�Gz4�;��YV|��v+gN^l���6m�M33U�{},-,�y�}�ln��~!k��%�3��R_V�6����1P���t�Cx���[�}'.�G�Gk��G]"f�uDÑ�T�9�!d3����B��Z ��m�.m�wӅ1øΨ��h
����4��lbS��V��$�������*D����hJ.��n�r�7&��T�i��,��ٙcC�x��J)H)G<b�7$�L���}�s��ͽj˶����K���X���r�@ϲJ�އ�Ĝ��ON��7�:��鹂|MǪ��w�(5M���l���؋��;S��t�U`�+�jV^����}7{�d����p7Ӓ���Љ=�'���:Y�..�H˞���D"M�?�\6Ag<����zA��[�g��>��3x��ǰK r��5ܹuK[�q,���f[o��kwn���]�#v� ��[o�����{���cO����P+��`�	|k�w���H���~�.��hh:_j��8�!"�g��+��·����
�{luZ�qw�V;��:>�c��?�����e|�����fՙ
�g�w��{��	��g�i+��jz�G6��c�v�h�h��I��r���d��J� �X�? {�i�d���X��[�4�w|��.E��c�Ԩ�{=H����4��Wo��B>"L=�|����r8���֩캆�l�~&2$G��+�oώE��Tׂ:1���������.�,3��D`��l:���{��W3�Z�7�
#������y�j�q�|�2N�3���c��YSHR��^ǕH&r����Á����t�IF�+�h��jiz��2�_�'L����Z���K�귿�o|�kX9r��_�\��2�U+�Wp���Џ�x����5����% �J��Bب�n]�/�VØK����R.������Ս[��R�I%�TX�@�@��屈	X�aFCkT��?���g�ܝ�v�2._�nm�E�]�#g���Ï��~�G��#�c%�}��O}��gp��z&%���m�Xt�RA� y@����`����d����@���C~�?2����m/o�^��{œ�u�:RU�0G�|y��^rS 7��Ű�W���ʱ1m��M	�h2�A�� Y��/}`"s�m�����J��$j�kD������6}�̽��Q�	I���0U�>`�3I� {�9]:g�NHۊ�6}����yG8�ާ�p{W�8��<V�����J5��)S����s����O����abnq�p&�A�������r�?"|�0_�b������z�*��^#�+J$��e��֫������y�kmB�KI�����W^�:>������V�V.U�̓�Ux�KA�i�*�����Cס<�s}{�Z���ʤ(�,��*�O\>���]V�K�7,�ĉ>��ɍ����Uh�:bӍ��^���#8q�,F�!ڻ�v����띝�mn�~k�ACҍ�&Y�k���-��=���H� \���?��@�U=w��Rsd��eC�{/���O�R�|{:_����35|��y��$� H7��	�h>�Ý����K#\|�g�qء��T�t#���O�a��81K��q�����x�]n����=��̵��S���˛rP���>h�A�UR@L/��e�3'!�2�f�h���V�<�-𳧐�ַ�6��e|��3B�M�o��fb$�.a��JÔ��"%C��>1��6�,���wu���|�RT0C�{��%�oL��%`���x�qw�����f������'�4P-W�������CDL��F�!�N�kršS�/]a��o;��.����H���^'�]�;"捷߽���'���2f�c�ry�*v-6mp�ma���d}i�%�|��������u���@��v����V���}��?g�Iў I�ܦ�?���df�t$D���IL}�!	������N��M��h���M���tf�Bk�v�ScX���݃fϟ���@�gZ�z�';p��.샰2��ԉ��&(� 0��xM/:_3�L��D��:A�.\e�Z���j'n^/xEOXc��p��~&U�����͚svn�ܱ[�3[-3��Z>�Zg��7d��ߝ��uΘ��33�h�RC� :��n^1e���)b� �>ivS;��>x�G��X�i*����i��{���w� :VP���`2R��0��R��tD��;��\�j$̲�� n�۸�y�n��^%#�cV�q��Ƹ�Fj�s�%�"a�zfQ�mvИ;��l�Ւ�Z�I�4A�\��u�ƌ|fH?,4X��J1���:M�9=؀R���ô:\���qQ[&u�>e�ǟۃ���s������%�Oa�ʂ	;P��g��n���v�f6�CC��G� ���<�c(�Uzd��g�H���i��9a��)�����3Q�2���;w;�Y[h��+������`2��c�1[����#�JX�4��e�"�?y�H���.�{A�*�S��&���\��$<�4���~TM"�T��]�u�~[);��O�B�������G���\��4��k+��{�}�>̒u6��	�=�{\���lgr����Ц�T���lE}��K��v�G�`��40�h�_A��2���Ka_�.*>O�l��}b��=�6sBZ#���@�F]Wv�rmW�Ru� ��ۜ�f$U��j���B�T,c�A�CI�0���#&�T�M�G�>����;��Ip�'Kpj/ziJɥ�Y ��]��Ȧ���������c��~%#�Y5Xݡ��Q��c�a��,����t���ӏ�M6a\^��3��y]N�J�]%07Sj(��r��v'3������ň`Z��*w!��V��N��k����k�|��6N�w�#cT��p0J��L��ސ��3J�z������Oi�M�L��8�Ĺ�tJ�i � �.b�:���R%���Λ�}	C�f��|Ʊ��.��1�:��FCTS��A�65���gB�7P�N�	'ўH��07gϩ�D��e.��@O)[�T�;�x"~2�v9H?��[����c��,K$u;�����P��؛0$-��z�L,�����kC�X$�ؘBi!c�m�X�l4�J�Z(*�)�-�E�Y�ci#3�����EI��J� �,���������hB�v��7���ޓ�lɛ�̂�)Rn���{�*2��8�n��
�h.�'9M�5;58c����T5��0Ec�%�d��\Y�'i����yml�FH�}�5:���{_M�EylV;��pXa��¡�b�� ���~x�s�7W-?�,��̺'$�%��_���y�X,H��V@��j~f���=7�v,�'��9y��i�s�1XhJIS�G����>�9�v	;Nv�]؁M>HiS�G"�X���[*Q�$����&�(�:�u�-�Y�p{����G����l`kȳ���I���'FvR��)�2"�� �]���QP���T�d�i-A����e�H9��􉭽���u
����1$ߟC���V��T��
� g<�6k��k��N�7\��������f�T�?�C~��I����#�g*6!#����:�6 Q�L̥��61��8H��)ㅳ݄����Y�ɆuZ��*�_z`�,��e	��jB��v�z�.�yʺl�����e"o�i�2v�D�S&u6p�ܲ�D6�o| ��l:#<�� �H�8Ʊ��2,;G"T�KR(�GH��]YR�iՠ^-����K����e��M=���"|���@�����mP��  �}=���Σ��a��2Y͘H<U>�O�^bQ3�
S�i� ;�zփX�#�A��YŌIA*�[ 	2���ā�����& �3L9�f��#�M��z��E����33dy$�?Y��JPV�o:�&��n$=���ɘ0��6k�ܱ��+������{J ��pCk�P{�8�K��̚��
2�/��g��T0���]܁�$���N>������AbY��%�%m욑��)Vm��U��-� ;̆�L�.�K�Q�3�����P��
.�=�_tz,��tb��P����eU&;|��;9�E��	!�1�$�G�͡����(�ls3uW�s�4
l�<�sx'�^z��?26����N'����0��d�mz�ӶR�@�ӡ�}+��>#��#m�U�ρ(7;���ə�7(qrK�$袘m�%qk{N�bo��OjL��̡ĸ84hh�-J���-� J�;p#��6IҵD��8�X'-' 1���{RKa�6'�)d���wH�g[k�V�sv�Tg�k($!j�'*�5���\�[�ό��fI�����r��:4b�l� )��ו���f���''�9���T! g�-͚��2�X���6}UM�1���w2x�L��X�C'��I�Yٱ��ٜ�,1.��l��Y��D�����b��<$Fק��)��,��P�}�6���%aY���`4���n�1�(�42�B�yg�!1ff�c���ش�_Sn�`T#�,c�p����T�l�]�)�6>�A�7;׶e`��v^�|?�S����S��F��7�3{�9��#����ޥs�]Y۬�t���x��t�%�J�``�5��Yc"�ӊp/p�������no�{��N" ��~Ѣ2G��z�m���8��za4���k�U�lz�D)�����5ܨ�R��D�{��������t�(nI?�!�W.��qΚv?��	{Lٛ�$b��U��	v2���>;��Kt�H�:�.~���Vh�H�=��	L�xw7cBc1�r��	Q�e�9I��8Œ�H@�nl� B�TEXu�[��ᆕd~ܢ� �]�|�*ѿU��u[�_<������zX\�����J�>;�A�27mU\e��CP�H�o����bd�A���I��b��('��D;@������DU	]�3�k�1��l�B��r�J\��EX4��ɲ���͝&��
Ft���ܜ�I���%F��ܡ�����+��0���~�B���J�ϳX7���n^�<�ōc8�l2���ʂ��W'�$`1�	H9����Il�\k�1[E}�a�ǂ�,� H"q�ܢQ�g�u�hߕ.t��C�V�#�>���"]�!`J��h~qQ�|f`N8 /$�L��(8I`SH�I<�ӫ�f��u���69K@~��TI�.�*(Wj�r?5�"l�]���$n	~�l�Gb�:}�^�	�K�2=��L�67Kc^��ءl�`fMY�isq���&�|l��� �r����h�ے��1Z�&�Hcɟa�� n�:0���}&K7͛>�#�>�Ū���.nyˤ� ʃ)Sf02��$s��Nd;������eb�=RCXrpAl�b�96��b)�drhWU�jw���eS֎[�p�+n�2�"\�PՄ3��NG�8��6�����	 ��Ł0aV�yk� 7,ܴ%�C3��Sm�h�߰e�28���앙��U$R�f��cɔC���̚Z8�vnqA¼����K�䰷R�"�cҭV�K=��PƑ�?~�}~�9��h�\ښ��s��@����n|A/g���Q��c��͚��&P�#�E8EY�@�z�ֆ�c�jX�;�����ڛ���Gщ+R�Hb��ev޼^Lk�������O���\�T����w�}�N[���?��'N�,Ӻ/��n��*vL勣�Уq�/�~�^�Mc�f����?�[�o���ui���C�T��1�$�I����P�E��N�����`9V&�ҰF-����y����L+Uc'�-��VGI
�d��D�����D�DY(��(_����{�{�78�gq��Qq�qߵ���������O�v�(��dcx�5������=o�qo��`������ҨpL,�������G�,0f�:6%�8�Iۨ�-�"ag��!ui�~g���,�~�)�9v��`Y&a�1�c++t�L����w�E��p����z��w8
hJ,*���}�84��Swآ�0GbF�Κ��~4B�E�J*_1��}*7��.����:��1�W�X9��8��Ʀl�/�KtO,y�[��f*hw{R(g�PFcaI�g7�ML�x �5�j�{���W%l��l��*�����ɌM�D�XU�ƈ�S�֔l|e�\�\�����rl�����vWu�Gڥ�������_}���&���Q��k��	h�(QE��f|�J؍��[ 6��I l�0!�߹��v�/%Ay�3��j{!�i�+�I:H��S�bi�Xsb��l�!f�v�f�������<�/�ta��SV��g�[ ,��o���=}��w��;@�<u��1[�;�|{3�3���ԓ
&0Z�P0�_�W�}���G�Z*��ɤ���I��=�����O���¶1N�f��#Lx�k�G��ADlH�N�,wX�+�`�zI��`̠S�H��0n<��Ȇ!{�iqq�,m���G�����,������-z.�����^��/~M��l��S�O�FR���%�5��Ib޽;;;�U���G	���� B��K�"�M7xveG�fIr���X©
X^9�}�c(U�h0��`c��븷~?��&޼��8���ñ2�Xa�b�,�A�AQԿQl�[�G�R��T�`e���|����EZ�s(�����Ǹ~��\9��#�eai����E�k^кrv� ���~'�P���'�-���υ�p���ȕ21�-���;ľv����Z��f�̊k��E^v�Q߳E���I��`"L��2������Zf-ji�(}�1�ol�6T5a\�� 0�b��4$@i�����X͈�=�V�������2�z�!54x2d��6��E���7�	�k(�����j�(�/ym��KG�1!BE�a���N<���:���e6���ve/s_S�(MiI��죉,��9s���_�D���������o���5�iGj.�`�'�:���L��T�y��.��8���k4Xunj�7Cj<�BTh����������Qq�V��V��!1��2mc��4�$m�\�"���q�;�������������6��]�c�6�mH�|H ���,5
4�rm2[��+	��mTf��}1�l�ԗ�ԣ*�R+qa�-�lP���hg7�|gz��c��tn-1��8���%�>~'��;W����mE��l>9��D���4_n����b&��̘~>��sX&��	s�t���A��^ 8�[St��w]*�_c�w5��	���%.�䇞�r����N�o��I��G�]��u`�<�i&Uvh 1�W��K�uGjl4U�(�+E�
U�p�� TF�&�u�>��X�*g7�MW�	�Vs�>�,������v�s���We��	���&�7m}��,�6�8�3��Mo��=9��e	�z��;��sRs�5� 4X:���ېz^��֊dEn@k��s�R�tä́�+�np)gM�چ���7Y�niJ#e����D �#���I�o5[�`j
��Զ.c$�X�^T"H̿)������dck�4�E�>�Ui���JG�h�l*m�څ9�I��J�QD�B��W�~@U���	<���j�����[I*j� Re�F���&u{���W%`����ܙ�E���W����  ,�2vh1�$p���'6\�j,�jh߉�=8?P���`�>K�^E@�mR��U��;$��;�Q�;M���0�?%l�*�ă{k��G�է��2�$,*�ޅs�퐊?��_�ah5񱏟<M���?6͝�a�4�=z�#t�MR׶i�q+�=����w��#�ry�B�
�P$�!�
��"tN���c���ͣr�q�Dh�;	���Ga�a�z\��F�xø�aVI�S�y��\<v
}�Y�e�YE�ָl����]�M������ZmL�gB��l@ϰ��.��R-�ُ>G��t;����8{��.�>ͣ�D���nF�ڌ���Y{�_�E��xe���Gܐz��'~XNgj��ԥR�w%Ӊ����v�%3�6V�;?����?�㲗%�"'�pQ|�z�b� �^#��d�5D��<Ǥ��]i�4����'?)$��[w�r�|�٘U0�<&$3N��4�P��I0�L�:�Yz�/�;[8}�Ν;#$����b���w�t�0��1� Ό�m+<R#F�⍐-zq�� �䄜b*����@a�Mp�Hx{R�-D��b�������L�9���^�X�#��g?�xu��?�����*a��������ig+�]�{8{����g���	0����)�V�F�b������H��]�>:)Z��|���9�rl�0{C���Le���"f��V'�,�h!
cy^v�4���+W��ׯߤ�h���ai����&��Oט�%���m]^A�����q��(X�Ug�&{d��E�����X���w���2ۨ$J#-��/r7Ǣ"�����%�c?Tޚv���ǡ�{��t��r-E\k�83`0T���UeO7	�B��۟��ۍ���1�^j�I%�S�����8�1�I9�72d�̤}���ݕ^lO>����j��KWX�u����{�\H�{�@%�`eclS���x���3c�i����j7�ٵ�N�ج����Lov�D,y��b�tZ{5���:<H�o~p��%�l<?�J+��-=��X�>p�q�6�*�=2'r5����Id(f�X�q���1u�3~6��/� ��O�rX�{�ocS�M�>k�W6=�H�h%l�售�pm�M'N㙕�-R{%��k����1�����f��W��&v�M�A�x�����F�M���d!1	5ꓴ �s�;�8I v���A�s�����T�厷[(ժ�7j���Ю"����>t�T�Բ 5h<�khn��2#��aI��V�q���z��M�\{�-�-����s�m�;���Q�޺���e�޸&�q
��y��{o�6�j�� 334�Us|$�I�tF�.s�'��'��_���}Er��Hm��%�m��/�O%�f?{ӾgH���fS�ς�J�e��)��)�,��4��Μ��?.Q��aـ��0�p�#�t����e>χK���i$�y�$�=(M~X��ӳ����:!�^狄��0�:1#���E[�����߃o��u����>��v�B9�Ps�2�yTI�0�����RQ0B�����We��L2�3P�&�E3�uV��H�M&�8EH�GZR�\�]�'�@��9����|��q��iZ�!Ο?�nk�n����h�nI�lU�Y`�"��1׵w^��9��
�rB�B�����@,��FwH���m<|�y������`Q8�z�(vb�hP)�Kdg���%=�ҿ��IZ=4��޸G�]��g�c|�&�� ��n�
��7o�m�k�x;-DW��K��RS�x����۷XϜ9Cx�@�$�A��Ǐ��v����E)��6��Q�9���| ǔJ��nS'Ǔ���QƶѢ�11�0Eqһ��ʅ~4>�zC��l�c�3Q�����9�}z��e9��
� �1�ڹ��](S���*�3��ݵ���'���U�N�܁��j�^t�7W�1a�S��c��X+�Ik��s9k
�p��B>��h��}�Z"�}_j1�
<�U���s _Oj.�6�E!a�H�]ʌ���yn�����ݥ���AXL�Bc�إG���G���ǉ�JI,?vo|_a��=lm����A� �H�u<�0�����c�{�ⱋ�qfq^l�Eb��b(�2(�.l�>u��9��ں|�R.�E�Y4�w��8r�T�R���=�b�x\����nWjzr������W��s�Tè ���^�G1.?�
��ܐ���c�u�WoJk��V��m�����ĉ����0�jK؅��=w^q�"\�x	'N��
}�k�\_[�N4��Բ@< t�K��p�N���7'$B�ٹh�߫d$߻���5㩰��@��,I{Jl�ܞ�����F��Ν:�����	��A��Lg~2ϢҸ��cc�t�Y���)�N�LG�>��3h��N���|�{��W%��g�q��"X�"��{9� ������݌c}�s�M^sHkh�����8mb�	�H���"�t�} �l�Jn�;��[Ӭ�&�Y��c�ֳϊE�B:���q��iR��87����J�!��}�	ܼ`q�fgP"���}�}���>��"u{Ub���NK�pp�żk����c�HG�zOYD����Hp3��6��[w��HLV-��J� ���@�Y����I=�J��R���$�R�5����	-["�Hb��ۥE��KĔ�J�J�G��^��߮r3Z��޿���?�.� z������u��r��1Q{���^��p��	�-��u� l�M�����L�0x�����W��Brk����A���N�d2{�*q~������+o��ի��%��?��H/b��v�5���S�󄚚e�����Y��+�7�}�a#��:l����{f�ib�c�]Oe����s{�Nf�dy��r�C���g�
͉�����Ҥ�܉`w�;��9�����	�>��� �d�	�J�:{&od/�����ӤTh�y�9�]�B� i��%��W��O�ħ>�W_�:�t����u�-��
=R��77�j�b��+R�#�0�;���-�{X�,����N_�����m|�ɏ@�Ć�]�:W���6����,�>����=Ie�x�F��>*��o����{���eVp���//����P�@�WA��<J��~���RIh@l���6f�W�|��OH�Dww;�[��E1X��8~\�/\��ޠ-a%l�̵��_µ{w�v�V�Ob�Mʔ�p(��F66p�sd<��[�߳������I�������l[zn��C��Z<£���)�<�l2jq��Ml`���gt��mb\S�^6�y�|M�i��_w��5�v���Ю����,�����)'�S���C�Y�l���N��C��'ә�!�$+`��9��ľ��P�����.B�?k��+�a�n��CJ�fw���%T��I	<!���������W��w_y	_8��*��>"n�Bl�Û$�&(������@˳��������[�����&v�F8�r� ��X�E��+��k����x�{/�3/=Q����(��3���������mT
�LG��W�_����/<B�ZD�0���6�� �t��]n�S�P�1�eu����;x�w�g�yrN��I^>��}�)���ˤ�����[�s�x}�A@aey��X��4��07=2����^����i ��i�O=	��'
}��́�a���T�7�jW��"�%�n8�%%Ҕ�4-T���1������$��e��ڟPa]��{9���>��Dk�� ����K�d���,����H_��5&�Rd'�K����SS�$L�����ƹ4����{-����x_��g/qj�3!�1���e�f��PX�n�?lS�Cl�G?�)�T��ZR���C�+�~�o�b���7_Ǘ���$1H��X�$R�;�}�N���bv�@��ޘ��Sg_}�RH�q|aNj%���9s׮��w߹��v�@p�G+B�����:��{��oa�^o��6fkc��r�Kȥ�x��4����N<"��!����{Xo���cO�g?J�t������{bt�&��j�=���#�Rk�94	Ŀ��oK$�믽J!�����*���׿v�]ܻw�q,1�hk'���Jxgc2�ȷ����gʿ�6�^��,\��v����J�U��}ʄe�[�T[ݍ��tz=�96�M1�>��Fe�Ůؼv#aÞl��9�L'7��kN%�?��SEM���	{>�4*�ӓ�'����{O���)	Ϗ=W���H�q��W�>�����cz#ni��Ï0p�G��ZsBVΠ�څ�%��1��Q��d ��{��{�����ҷ!-�o�]���Vc�U�!���rr]�~����B�e}*�ِ�6k*�f@���'�@��8+�>ũ�=b���۷�V�CIW�x�bXg'����3���k�������5R�hE�-n>�s�ԣO�P�'�"��<�;����?�+7oKH֘���9��
�V��{���?�u:�6�-�HJ��6��{�m�tv[��7����VV�ӿ�y��R���i��Ѽ��Ja^ɘ���W���}A��K��Ϯ���Sx���������	4���2��#��P	0��y�~�[ߖ�s��f0Ŝ��7�n,I�@:�����rg�Q*�B��Dn����ð�i�̑k�k��7/�9X*[�%��Jϡ{�<)k)�Ӽ����!'�	`9����Ye�|63p}� Q�CP�z�� ����)�Z�ʭyq�I‒��ia.F��J�yW�"��T���f�U�kH��O��Z
�k�0����R�?N�͛��<��a�='�Ó�1ړ��0�3�0c�^#3'�Mn��5��6�i\�r��׀r$��,L�qe[�H�t�� �\sGsf����m�2�V�g֦L�z׀q� r^g{�N&�T2J�f��;�雭�pk�&6Z�X�+��:�U�^��k��y�R�J��M�#����dqsEE�g���r�\r�6[@�y��A� o�>}c�
�m����Lc��M�n���1ʤ��CU"�8C�/�����5n��(TQ$V�v�:��<�M��=5p��슘S�<�7.�C?oc@ל-W%��B�?����_�:	�Y|��i��·����Z}�kb�-��O��[��ݖ��El����W�B���F=�>'��e����t.,[	��	�_YV�O�:�F�rL���Y+F��S�6LT�N�c3R|*�J1`Ig��e�S�cW�[�B��|Ω�	[�6�DԆ�YX�y���fT�e,�j�|>Ύ6���G����)Kȶjv����圳�f�qCΑ�t��H1����k�����|v`����=�S�	��R��n��f���Yͅ�&�H�u��R�L�	Q2h��6�Ö��[�){vd����8I�ލ�"�]�Cʹz<�OgH�/���m����!~�g~���I���۷����۷8�_2��@
�/M�0��v	dzR��o��f�p��Eܹ{C�]?�5�>}�Q�KL0��v�����Lbǝf��*-�<��=A+�1��1�Ao�asb�b�'Ϟ��b���>SS䅟�K�������&�\��"�a��X-�-��m7w�g�C������!���O��{��ڍ[���&�L�G��?�}�*�F���q-= �%�omW���[�ӭ��$����T���9he�|�Y��]Ԏ}d��Ԋ���AV�ݴ4}$}��e҇ �8�jd����u7�Y��+�Y������4 ��Si������}��I�P.�i�yf�8m������s�R���Ep��-1�$�0y�n&�9��y�Ml���?�g��;�'��<Ⱥ.[�཰s��a�K�ɦ7k�l֗�'�YQl�,� �vf��\n7���AZ[7��r��/���;��o�]<|���C����3xs�M�h���	��Ի(�E�ap��6^}�XZ\£?�h߸N V1loH-X�Ŗn�6��"�CKO�!��!��Y���Ԫ��v$ݖ����[�z32*�tդkV���P��V�@:� f�`l��8q�~�~�ZCڙ����"��N�^��������X�/}����`u1p#9���=߀X�@�{��� �[=4�~��"6�u3�E爹�ddM�b���� ^�
�.o��t�Q�r���Q��K�X9{��1���<�}3(IW& ��T�� ����6<[I{u���u=�l��^%P��au�ס|6���:�Ek�7)n�Ls��M�T?)"�A�e�Y��� 1`�`�M8�2�����p&C�u�թ)Oq ���N��w�	���Am�ۼ�m� �d������4�`��!y3�r��w��d͉M���&�+8i�(�#$��8cS�A���B�1���iM��!�z�$z����M���+��?��=�1�޼K�M���Q�+��2��)�O��M'��m�茇h�z������揝F��-�J�T(�_;���=�ޠ�A�*g�~��\нuIſ�C�w�sa..��V�Xw	Cb�u.,�7"\�b�4��²�|��}�0tO=�è/��Z�\�G�?�
�1����[�&6].��o��o���+'q��1ܿ{�X�ڭ�؈�=�61��w�cqq���*V[�?���'&.�14��\'B0�jQF�4�fF"�����Z4-���ld/�0� ]����Yl��p��̤~�� K� �a¨���qZ[�w:I9?����zG��0!�)evsf6�?�y����
�l���ЕЛ&˜pL^�wE�:V-mZr'b���@�|zʵُ�Ȫ	U>�Il���[b�tjw��:�*��aM{>k��'�#7w�&N�,1�6%�U�?�-����*6��x�,L����j@���.Ȁ��\N�������c�n �	uTzW��K)5��j� ����~���R�͛x�� *���3���Fua�B�-�07��qk;��"����sP���k/�����q��Ib��;�֢ �$I�������=oCls:��<J�"1�Y�=jiۛ����3�⭷/���gp�����v��樋�f ��"5>,k"��~��n,�c�+��Ɛ"%��B�6��ϟ�
Z�U=����_G��£�L��6=#[a�t��o��f��B�HªG���{�6�l��;�zJ�U`�M3�����_m�5����w� �$vQ��4���H�Z�ĴƎ�%�w���`��fə���.�N*��G��
���Y���%�٨���5vQ4I��ʫ���8��X����M=G`s�M�jN@�P4��{�ZȼHl�F~���ʚ1|Pu&�"��E�xZ��s�ZI��H�6hq�~�R��#N�
;���D��e8���Hj�
�H]	m���-��#�Z�7�l��;ȘfR�y�	Df�dѮ��?6�@ңˁ|l6�	ja��z$�q�Tgڨs\���,����k��WM_�u��`�O��hH@q��ϐ�o�����F�4#e�z`T,6ݑ*ag��}��mz��bET������o^C�gz}��ub��(CRݻ(-T1Pcb֐��onl�
�����"�ҫK/�Ko�:V���WN��]@L�|~~s�x��[���נ�3آ{fv�l��[�q��=���쵀�sL��+��7���1V�oag�COG��3�p4}�ja,�
R�X���q>K�g#M��4lz�Y6&K�1�=�	�ulǲ���l�3��c��|�ɗ��Z��M��u��)�ykoU�:�����Y��Fx����u�Q��'��l����Rg���4�.���%�o^���̔�~~KۊX�M���T_�|����S��9 .P[�⏶�
��-tȇ�1��˝{����z����sk#?�Y&�W������ڔ��G:z�%���k��B�8��%��A�����^*P&�S٨��À��V�+ǎ�8-i؂���4؞W��S�����[+F�prnn�=$����FX����n�Å`��Ԙ�'F��ӿ}��.}�
	c*�����ZT,)˼�k@�.��oݾ���JN�áO;ƀ�3^`f��ڼ�4�j^�"�-�gH
��J��w��Zci���x0��lnKQNl��:�N��y�9�m���GO�j��˪>I� M�E�>`�L`j�r?"�'φ܆�!c��L�V�b-�m��:�Tn�E���(4\�g1�X;����{�4o��NA^+��y�1�(���b��; �$��֪0��rn�����1�E�1?X@u��`�����h� �'O�CدeUbW�?���e��lf��<�����
�1���۴�#�&�T�Ϊ�F��>W�����LL\�^�o"����ɹwG�LhʛC�e�H҄e,�}�׍!�~VP��N�g��t���p&����\������l��~l:cJy�6�IRn\�YR]
����;aRH���M)��R�E���
8fR]��yf�y)��7kq H���-:���m�o �5�!�����%k�+�Q�B���q�:��OcĶ�2o�P>v����À�ۂ��=b�7w����E��&�Ml$3����#b���	��
�F�
�F:r!�>W+��T[�k������.�2�4�Q�<����/��U�Ơ(堥:Y��\�@s�7M`=�����JdӪ9/߻tSQE�����v&��֎e��]n5�cq�8����!��m�Sp�?���K��|ʴLa�0����0�
mM�u({�)8tDd�XJ9���*k4_�\�>g T��F\�g��6�+�$#��i����l�-^�;R�z$��M'��[��q"���mk�iD�4܅�N�2,$������3we�)�1���eV������#{
������{��@j��-�I�8]7#m��ˇ?�~�-w�ʚ]�q:ϼF����=%M]-I��i���MUď�p)���y�0�i�~c!�(y�dץѴ;�ڟg�v�Eq��veu⅕�+��U�d��&�ܣɰK�c��Q'���A.�����y��{q��a
��x��{�3���H½��(s���lf���y`�k���vlU�H&2L slUZ�=֑��T͈`�5�e�p�-6b��4�(0ōy\w�ma��Z�8��u��O(o4r ��
�m|��[��;�MM��rM��������ݔؔ�v��|;�RV�N?s�p�Z�g�"=,�H�X�_�L9�!j��2�baua�<���=�2���bY/E%��fɻ��i��hf� �:��g�H�$�j�1���v�)ﻣ�LFyG�>x����G����S���o�����]�7'��=��Ӛ�:~����� p�Q���������ro���a�q���,K�c	1kT� ��26�/mp`Y��X�B�e]�����/l(G.}�ڙ�JڒD�1��#�*�蒑L�Dc8@�
�p�6�$��
)�_m�Xۓs	��ڐ���j���F����՗�_�l03k�V���Z�窅�d+������}"��樋�^ZIܺOsϢ�i�9�G㆔*0��L/-/�Kk�Z����ڱvf-�@sH�G�T�s. ]��Z�m�)���e[�^ �������hI��N�À䄗����wL3[����:������(ɚ��0H{�œ�²6U��0���#n9���h�J��I�0��\�`l�MVN�I�?�l��7PZ�k�?�|��_Ž�u��9&��&�!e���h�i�������EO��.%8�iE�̓�!���;m�]��\14��#o&���2{�Me�
{������I����8L1�h�!w���dU�gH�&�~�i$-H3Y-kr��Db(�]��E���X�����3x���t��/Am�&�Cu�
����������W6Wi�z �|�)����b`��_�5�(��f��[�����qt��S. �j�*��ٛ������W�g�ʔ�D�d�݆���e�hB�SP�����g�c����˃��l�A����A��׳��F�A�v>B���6f:��ĉK�d��30�-��	)�/�}��׷��L�s2e���]�����1�
)�q���~��:��Tq�;�\o�h wa5����
m�$t�hR�a��\��+vB+4,���
�&��́O���J\���c��\y_�zdlh�T�7��Le�U�z��\�^��C��$7z��/�E�G��A�ρ��5�q2M��4����i�qΫ���>�q��O�4Μ<��ƒ؝�1�_c'd,��вkâ+�Y�q6�F���Qe;}"x��@x��r�
Y0�p���(�;��� �s�����:�#67M���{O�1c8�����Ց�R��^�͏�^f��*-�a��z�JZ?:�5��s�9,S�7?���~ǃ���|ޑ+�蕵l�`�q�~ZRŤ`���6	��c`#k�[*Ϙ��h��0��7��D�l���}�܋T^ V{�l@���q��jA�RE"D\g��z���s�\�c�7�?K��Xk��7n��;�Ą c>P�Ȱe,���� ���ٲ��6s�f�����k��x`��M��*��X��1�l�QvFL�����Қ�|����\����b�"NA�XJ;�9X1���wUR\�7q���Cf���r��_�;?��}�3X\:B���S0�J\Dxp�3��Ġ�f�5,�.��,�8�<Q�RR`�s�8-�$�ɢ�ܟwn#�]�_�F0F���;X��:N�� �'܉"�H`mw���r��q�C�vz��v��z$B�R2uxͺn���5��$���T�#K��]@��s��z����V����^�m_͌�[k������@����&�C�4VV��Ê�Ry}J�\�.��-�0����&��Ms�w���5��e6-���*Z��<舗/�
I"�p;,r݁�n� �+V?��afŪ3Zb1�R�-ئi$�z�ia866��+2� ��|�3.���=�\S��2c!�M�T)�����4�es�q��u����V�����W�a$6�Hj�i�	�1z������q,�e���A�G�[��t;V_�O������1��`����	�f�IcPD�~�&X�
����:�M���L\fʎ�S�`���������̜@QV������_@�ۑ(�U^�x~��3L~6�A�櫗��o���`kؑ�^��N"�7tll�.n��Gfj8�x?�ٟ���J�_���m4�����}�O���R(j�<�E���	k��Ԉ�?������DfU��L��z��rbߦ�]J�2�kϬ+�7_�I؍&T�:"�:�z���q��.B�� }fw#��q
n��t����K�;����0����&ʕ�Z\���$�)bX�ɳ��˥�Y=�ޚ@@��>E�H@7��ؤ�}����6E���LD@�q���[����3p�?��r3�2m�2ר�M]6	0�fO=�TָMy���`��p ��b��.X����ȟ���:yY�1&!�̓Ϡ�X @7�g����-<����W�"���/�>��3b�Q{���h��Fm�1dbl%�m�c��D �D�yu���KL��ݩ�☴Re�*i��f������o^�g"����^]��D������G��
F�V�A���O��2fI&�<��-�H��OU�bne^ƕ��'�α����D:�l�W��f�]"s���LcǓ�;LhO�MG��ޝ�?�>���U��(xZ��,���ͷ�5��
����o�I�O{L�XsD�vZ���C�,���FS��<�<�E�)�Ur��_��֙㾢�)��KS@�8z�z�1�zQ l,�ɑ}�
�7��*8�Z8q�T(91��0/�\,�҄d]�k��#�H+��'ǹ�!�mq��qw�kW���}�1�X�
����v��"mD1*WضH�c�)��mj&��8��8�����{9MR���@���3�qŅ�N-.���S�3�ĄeLq�����|]�1x�fJ&n8�����'vO�]4�w�b@�zX�>g�$�&h#�������5�@�DU�����tz�K�/�3�����"قڵ{k����_�+o�DSB���㹷�'��0=�Q�y��4c�R�����F(+�� �`����ui����{0�=�3ˈӗ�b��yug_��wQ��#� ���8�S϶`4	^��	�aM��T�ӑ���\oC�N�;�!���o�zk��t �th�^0�"�F]YA�G(DJ
�IkQŲ�U\čk��B�b��b�'oL�\`��#�4If���UY�,�klc�Cn���lAV�%�)*ٻ����K�o�8+���M��h�W	^�m��"k��v5�!��c�J��Lg@J���	�;^#���z�v�I�Nd��컑,���G���D�"���2�'�hFr�����C��p��tr	M�nwOlf�dL�]�fm&��I��P0cN2�w|MJ)߻:yL���.0ذ1	�1{��[��2����E:7m���$�SJAI(��KGR�96p�Рr��@�0���я~��W�� �߽���^�
6ך(.4P�d�u�#Rs�v{u�X4�=�L��z���iиV37R�9l��n�����E�s�L��Q-�^&�4��ł���Ʋ��t���'W.����J_�t�ۿ�;���{�_��ڗ��Ee�:ys3�rs̀��=8�B��6ۥZ] a��AD̖��N���$�Ieg&	��ϓ�AUI��p��.�g(�W����������K�Fq�*��b��a�I������ji*Y�m.��m>U�����{�&�<]���d1&Ϧ���3C�������k/���'����
N�:�j�Fs�C���R-��*�"m�
��Y҄�=��6vZ��;�Ĝ��,$�����׾��;��3ܥ���IR7����Aي[f/+	j�M�Ƶk��/~?�C������ϰ`�)�D�DRr����gq��Yb��aʾ���^Own��=���$��MP��-���l�:"\�8�����{��4�P�<�2��o,�7
b��VI�*�3qX�b�Mr�>j�Zr�+�}��48[���ב�L��pF籅E�K3p�>����$��k�Ü�-���������k�:ϩ�<f��Dڸ�jsw�� ��^|�Ul�v1"uw�lQQjwWN[�3��|�ݷ��o�<~�>r�	%�����&�S"�h/򵀤��#Ʊ/�ǔ���ky=�^��m���Yǀ�d�`2��>U��dp-Wb\��+�a��bUbmXN�X-���{��� 4��k,�;��i���<w�$��-�y�
v�o���X���W��4��@f櫒峽�%9<Kc�����T)"U�H����������+�i���Yi�$��|��3���%,@���������ĩc������">����?�s��e-솔[T+5�����t�5)\��>-`	��7�
m����B�)q�;��:��t!���y���"m��}A4.�wg�*�
ة7�d�p��X��3P��-�I:�*2ʕ������'YB��5M+vi�X���W��Н����1���x�-�������,~�3�C��
�(��V��/���o��D����n��@%#*�HF�������e�86���-�?��_��_�*�i�rg�:�D�p�����sv �=���_��$MH�$%,�m��ę�z�	��] ����I4���|�;��?����2�eg��I�>W��(3�f��6��b��$�I'UR6��s�v�6�9G������^Qv�י�w�͹r@
U�D$�D�	�")�
�,�V�^���=�3~�սf��t��Y-ǖ(��H�")fA� �S!���Vݪ��9����s�(O�X�ֹ������=�"��,Az6�.'��M��G�Z�ց�{�ֆ6����`u���a�[]���*�!��/�c g� GId
#Yq'�fW��9�g��W�{�
�] ���H���sd�^���cCx�ދ]����Ɓd]�dh_��)��NF�Go��x�bu14:�+S7qw���_�u����8
�(�,j��I;���x�8��"DHb&�J�7
d�����h�@��,A��tP�9�R���j�o%s�p��ݹD��NX?	+�g�L��L����>��y�_���B��HX7�����[�6�Yi���C�͋k��|2JcRּ���%���b����%�_��o&t%��n����3*�ҡb_h�K�L������h A�������&Ӥ ��� 
g���
A��wN|E�՞�B֨
66{3���kF��#��^�����(���Z�|j&N���$lR��~&�f�����������{�E�>ǻ�^��ɚ���yi���:vQy�}��J�9g�Z`Y�gvœ�=|��	�<=��U��.M������P�ӎ�M2��zՙ�ub:��"m�&�\K���̀���,�gxI�3�Q2?���	���`i��^�d��_/���m��^IJ���	#�()fFs���[C.??��*ϡ?>���ԁ�T�Ke� ˤ(d�A�J`>�42��� 6�G'�e�զ����*U�A�y���{��&+�%�\U�ɦw�4ӵ�;8u��x�Y:�,�/^�(h��o����.;�.o�����H��{?SL)˥�#	�ɟ�d�-.m7E�4ٕD��D�^�Y�ʒ�#v˽ǡ�	�����x�=�w�3ᛐ�٬X�ξr@�GU��2M ���G7Yޥ`M
l�C��u�텃��O��j�a�aU�������M�0G@�2,HX�!lP��0���Y�]� .5'�G�����逵h��t6�m�ؓ#�x��WI���,��s����e��Adu�I+��4�ʑ����I"K�6�7�����dqɣ��!B��9��l�i!i���FB!aBt�ʆ�3���zd�p:����[���oѸ�������-��B���;_frBʹf:<n&���nq��!ev�B�~��{Q'�Z:Ȕ�q��)��$��H��H�����Ю�X�6elU�f���5$����鐄hN|0����!�*��,��^�X��%x��I�,H}���EߍX��:�gΙ�<W��XYrV	����GN�c6�/� ��$<���d$d�|���.�֎Ep��{1�&d',�����;�8��Km��e�"�0N��>e	�����u�SS?���+��Dr
�������"T�Q���K

��I&��|��"��Z8%��&��>F��]���3sI�kJ߬��{��^�254u��)���eV[�{t�P|^�Fr�6���s���ط}�#~+�}zzo��&��ϊ�Bފy����\����)Qzy���8�.B�\�I�(���H^�.eQ�:��i���{VY�,k墓qM$����=YH	�ʍ�����ywF�x�*�D�G����E���.0�*���L���f�r�>��5�\5��?�z_[�@yhp!NR'��&�9@B�W���>KH.�>��)�%g�����N"j�IK&]ɐVf�m6��,w���H��t�"�C���I�D�B�_�X���Q/!����5S%�Ca�$8Hȸ=���!A�T~dg�U�;�� ���[&��Ԅ��n4}��E*Hp||�����ic�Hy#C� Z��+n��5�eT�\Y����
�|_��t.�����>�x!E�G���C.�����
G��
��j��"��+{�d&0x�HP�&gy�ظ�˼����4d+BX���B�wl����b:��35�޼������r��_��w^R�s�ÂIA�����yI���_ޭ2?d,�����J��ne�5_)[©A��N�9�/���E-��lg�ZY��/�[��,6�
�	)t٦@^]O�O�}	���]6�-����,M`�R��.����'*�_� \�U��26��\��H�K�հ*qe��RŧTP��F�bל)�[.i/���ÎH���>���wF19=��hS%��)A�/_.)�Ê��}#����ҔՒ�WE������g�epdXP��F�s�v䬖mt���4����<Zc)���94��rު������HA�7��Q��I�GY|��L|g�t��͒d{8�BMe�c��ʛ�K�q�V$g3�cH�+"D�r���.@���I�TutT&&G���	�">����B�C�/����-��t�!i���\W�����qҺ�+�Ll�I�W7�X��/JW:*4��M����~>��T�ИmFP�b�]�����зd�ͭ8��;�2�Xb�!jw|�"����bs=�ҿ0�����c	Rs)$�xh��t�>�>�[rV���J��"���ڪ��Υ���rن��ޛ��-"	ZbA���G���+1��Pf��A{}3)���v5H�m�6AyU���R�iCm�����u5�:�nڳ��b||�9=�������5��*G
6�L�jc����t�i�fsid�� �}R��R]�p�(2���>3uь�J7*}�t��bݲt�^�zM��t��_QR>Ƶ�7��=���ݢ�% E��F�M\��Œ��Xѽ�P��ĒL���,2^��vY�5Y;���3�����˵5wu�욟U��F��K����t6���!������b_�<P���r�w�,�޾(��~*B��o�9��ꭰ���t�+�J�	�|2cxf��[[#%�vg9χ�;�腭PUMr(g��汶��|k^#E��n��\�0	;�0���e罉%=ش~�	IrbpI"~�[�B:=C�^F&�Fw�r�/Z,���O����K$DKd�g����#	LR�-��)<~ЄHHG%�m.>*��p����bA��H�l�uv!�@�h!�˼ݒ�葲L�Ǚ�������(�R���[�԰	VV�)�͉��K�� ��9,�l�ǫ?��(|�Y<���\�y�G'QJy�5���\W`zf�hM��4��h�o%���بX��m�Qm��J�8S@����3u�֮�0��9i:�Ǧv�L����>\�~;6l��7�Ҏ.��w��^�	��	={�-*v��8�5��1�W.vY��ψ���:8��B���.y-+�� ]>��u1D|��Q�4lz��B�Y8�Ǌ�<��cX�҆R�	z�� �fgp��	��P���γeA;��ghm�N[KN�����t�Uf����^1m%ũ���gR�;�n'aD֒핒^�|��sx��Wq��ϰ���o~��]@Y2��"K�L����B�))�����Ebt7�A��ҾKU~'
��Ѩ}]��N�'�љu{��@J��ŋ��J!8������,a�3q��Y�w({m)�g�������ֱ.,���%l��EQU�곥Q�x�V�La���v����؂��EQ�*hk��Cr@ԚM����deb���+7U�W��|߬�/��̠2�Z�V>]νdD��孆��&O(��u����ɆOL���u��4k/��"fI����%���V��޳���a�}��{��ܷ�#�XҳABZ�>=�raJr8=�.���%Q��o ���y�~W���U2'�P�.��E3q�Q������W�~�)�i]���E��2]�%���F=�Y���$�}a/�c^�rE�����"�Ќ$]��$���Ȩ��p��_y�P�LA��*%����֬Ý�a�y�#A�V�i��/uM�7�0զ)������AN�8��1�Y�ARV��r�~�ڲ��[M��]
/)��%
:��C�3W{e29��G�m���y-���{��k}���__��%"_V��rT��M�2Y�X�،��v:C����=vCS���5�t����7�����M��h��Y���F����+p��Զٓ[V&��P�0�U.�|Yaŕ�����,�y;�z`8e���:k,s:�U��VE��`��E��ƮZ��h׮Cks���K5��������W���`�5��D�QU�4O��e���'ȧ��B�a����Aׂ�JW ��o`�@P�}�VYe�X�i��~g\�x�v����%�б��8�����HA��ls~W���8�I7�>\�cB1�z��Q=��5��8$���,�����f���]���~�Z�CZl��'*�Q'Z�,����־���i������Z�Em]���AC�M����,(~���d|B�6�5� ��Α��=��b�W��-|�~���Sh�E0|��e�g��Ҧ�Ӛ&[,fe���%�i,��!4i��s?C���-���9r`��r�8W����^�'�������X����-F��/�k9��"�FΤ�(:�I`eCTR�Z	�����@F0�CSK3�߿�4�/�JB;*y��=wr|���d�����s����"\���������Jx����*v���.W"(��b���2ڵ���	a��x��Qt/_�/?xH��P�BG�al^s��K9��4�jLg����U.$�2c+X�����x��!G�v;(��]X{������Υ�x���o������~�{xp��8~�c�kF��W,_I�c38���R�F�ϙ�sq��*)?:3.ZW���WR����0�s���
�ڦ��`�4�Ơ\%��
6Aq���$f�\��}[v#@c�E��Q ���g�6/�IJ{uě�37��.�%êPl
�q��ΊW|��@��E�YX��-i�Ei�NL@��+�;F�_��Ew�2��8(+�˃����}��w�и��;��Ѧ���'���쨉j�ʽ�w�g�Sէ|��_��N�-�vͽ���U�^�{4ۚ��Tk ����sX��@�ݣ�1��9��rJ;u���cX�u��-W�u��FxC!0��Þ�'���	�f�M��s�,�SH�� a��zl�����q�)�U��a��]����!2���Ν"db�cҦxȼ(e$�Z�Z����ic딥K���A�6s)ӎ���eB1��t������5�pЌ#�%K�V��B��lr3�ū/b}�bĬn�=�;�N���^:B�"/F���6�G��lх��5u$%t^��E��.��	di-����!4�@�.*��9z��'�������Nݚ�*<��p	�˙�K� d�O?N\��9���/�˖f-c��D���'�:���1��4r>)tQs�d�&5�^� K�ϧ�,mb"!L���&_��A��C���Ճ�K�ҟ���]Tr���֘��#�'/���������@Z:�R5���5k|�:��ؕ�**�%�e����6+������\>�|�' �3�
��*��[Sq`���Ң��1��04������p� <���Pt�w���w�����ڿ�����$Jt��n�B~k
��Og
�~-��2�9��2�����tƂ�p�߮�;sV�R�+���Z��^E(/p{j���?�ɨ2*m�lL���4�UO�vF�<1Nca���4�5�si!���0���?�Hpqr���$Q�rs�'QGhCr}>��!�Z$S�Y�|�П�_��*s�d�<]��4t��k��E\?�)B~z��6+�O6[�
�/�M�TA�+�d�Ӂ���H�+|T��M,*� !'e��<:ڻ�7b.����!!ǉ�6�`�����2+&���h�w��WvJ���_��N��s�m��az�xw��)(v��
S�q)���	��W��B����fs�S��gT�A�RI��m��yG�U�mK��+|�$Hǲ�����'Ϟƞm`���d�Ɣ��ST��Ql,.��ˮ�Qf2s�2t�m1�$�b;(֨�����׺�>ј���O��kd4��Jn|)\��(���Х��!��c%)�c-�U]��]@,�M^黉��|���=%AR*��ǖ4j�U9�@MΪ���
+k�n�1�J���@�<ڝ�����'G�ӗ^�o?�mD8�Y�	��/ȕ��dz����v?e�:�V��y;�P�-�޸��H�Z%.�W��ކb$�qNON�O<��'>�����8����T^[��+�.޺���L�>Kw�Ђ_�j�"9��ݕ�	Z���(w���.�W�[�(TGJ��\�������K���	ޕ��5XGؕ�Q�0�е �cn�"����ML�ڍkh7���uܷq&G'�J���Gg�"L�c�����a?�� ����`���H)_(.��PZ�~F�\�\)�|>	�4x�+��4cIYv#��ѿ!T ����SM�N�+Ҡ�jɦːf�\��E�7��qZ٢��J$�ȗ9:1e� �����'p�� �z6��c�x|v�=����F�Py�.��al�a`dd�1�&�ͤ1N�X�KP��t��7V_�щq\�qU�M)�D��Z�"܃�����0*BK��ݪР`�
�<Y�?�O{ϡ��m�-�����°DQ���~hAQ���D9`HɩӮ�br5đF�._��U��@;�@R�f��~7�rh41�#�>E����]G�-aK�0�$�4W�ŧp��Y��13�o�����2_5s��<t�\���wC�*c�S%��}7��|o���P���+~��_`����-�#�J�A8	�*ٜ��l]� �+�p�N/rfQ,DqYh���mv-��]���B
P���\��C�3�ĩ��r�_��&��؉�3p��5t�,#�W�:2Jg���?� �#(�8�ِ�<�G�8��*��-�:.��a�h|>�Um��g�Ԗ��%���<kkL��3�w��J�W�Ĩ?��~���D�K��oêy��Y��˭�/[*�T�<��T�������BBq��K�T:�E�XJ�r3�}S��RZȔpY�h%���<���#��I�CX������i�<He�H�cI�"�>��U�*��dri	Z�h�3)B��<y�h��2�xb����#�õڒ�&|^���.=�8�
�]��X�N]'�ފ��v�?g�{�޹�^FT��I�Oaj:�4	�x|	B�h��H��1C��MH��k#�j�I��3���KD�PR���*h��M_+�l�WTb���\�e����2w��*�>g�16zW���⛤ �*V
�lEק�]���[!����-�èj|���#�̅��I+�ZD��չ,��ϰ� �U����??�ϯ]�}�֢�֕���իeL��@��+�q�P��1Z_�����rA�#��=����E4ST-�2�f&P���u9�i�����ڍ��[��w�	Է���g��U��W5�l?/=��ef�:�oH��	#�j��9?s�w�$�{�T�Z�sV�Χ���J!�0.�����N�oz�Ʊ#t'�شr��Ju^���?9AJ��I��|Y*4.���	W��E��ru�g�v�ڂ�ι��٪
-��ue��\��?זI�j%�� }�s�犐u
,�N�Mh���e%I���ҵŮ�I8G�L��r����F�������+�s ����E�'��ͦ��ŢRI����'���&�.���ϡ��--�$A>Vߊ��	���m��9A^R%�*!O��:0���T�������g�{Č?$H�ɴIs��ׅ͓���M�r�I_�hr�:D�>֯!tv�Dp�tw�Ĳek wu�
�*�4��������7%5�K�n|���/'����y���~L��º4��Ƶ�[H�`�Y��Ջq/$X+��YQ�V�AN.'7��#��c����" ����+��P����r�2Y�A�9L�aTMG��U爅��{�dk���è�]����m���L����4�C�t���HH��@�K���k��LqY%�c�T����W���Z�#��\
ʰ�֕EE�D�?���Ԙ���Tn�f�x鈫�5���`��YN^��S�Y��ρ/�.]l�%[�S���k�b|�y�k>�]i��x	]�L��KS�r����:�����i+��}��h�zB�Y:�S$&�3�<y��,ə� {N��N=�����B��e�5j�zj5�4��斮M'h����Ϙ����|��_�'�(��㵪�R��n�����q�*��>"i������v�����M̐������Ё�%M�ʵ+b~��o>�Bb��^�.��#�-x�.���װ}�NYlR�hj�B��U8{�n��!C�q��2z�l��$
z}����굫I�$�<L��k|rR[�����W��a�ǥŉ'H&i|Vj�M!i.��	c��-��C_%�'�Z�Tw1N�I��b��?2���5���`��͸x�<��	c6�A6τ��5�DO�x8�1#0�B�)Z���XPE��<��-� �C�c2[u�P,�dy͹t�$"�.�G�.C*�R�
n�C��+�q*��6T�����EXp�+��v�6���㯼��䲰��ݸ,[�NB�B/����xzZ^瘀|t�d��s�%)���M�^G��)�W,{>/�]6�~�/��2VM�!�p;p�f.�6h.\B���Ec��$}�tu���Լ\Ps`j1]u��ײ��������V�V{�\����TX���q�x���[�m��;I�*���
��� �Ɲ����i��:�EG�x����B��t._B��8z,�)��vo���wL���YT�g��6��Ҟ0{� W�3��[��rU*��!o��㻨H���΃�:�� ���p�L~�b���C�;��3c��̧hnh&�5J'�Z]Ӓ�ʄ8-�f!?�r~$R)B�%��*�0��qn,߰�H(|�Y&�G�v�0�LK]�H"�$���/��������d��+�4[�H�d�fQ�x̠vM|~��>�<rE
��sy)��hv,\�][w��~��I���HI [8�ȄS3S��_����}=��i�IQXҔ�.U&��0�޺us��S��g�1[H�&%S�+de�� �s�]s@j�T�Yi�j?9�O�	a{h.Q/�Y�Mh�������(Bሔ�NM���ށG:��7o���u[���fE�������9ޖ]U�&�s0U��1�R�5&vU�C���,��	01	LN�^�܎:H 1�!��s\!�T�MK�~�Z��:0���Aa�*i���RȌ����UcQWW[Oɚ��4�r��V��V?���Z�Q+'ړ ��p�,�@{�"�x]��+�_\~���&t{[;V,[����ݺ�D.��,�3+���L-`�.Y�W�����5߿?�c�"@��{�(��Gw,���BH�AH�j�ڔ˞��Cɯ\t���yŅ�d6-��5#H��iR(É9\�� &pl!�pzn��IN��ո;*ယ��X��q��rv�kv�r�Jи˜���^lq�n5��Il��E&6.��Ga�������O�#�js�+���c��*��[qh��O�'Y9��:_�:F���D�.)�{�f�	z�A�hs�$�d�ee	U����Ӹ��O���%�o3�1l����Y�s9$3���=�p��z��P^�W�oe���dnAoL�@����5lBH+� ��";;C�X!#@6���V*݋�;���U�q2k8X��Ё'��?�E���2��,��#e��%U	�"���q�iܷ�o"P���0�Ma23�$!��i�g�Ad"	�v�����-�])�����#� �wk(��Vn¾�{��{9��:��i\�y�.��dÅ�E�E���"><�}[�����A*��Z�S���1<=!��A׀ր9$��F�:��V��9���R�0�c��N,�3�i�}5�F1U���.Bck��ي�w?�����aln��?btrPރs�q��G煫�v�݌U�V!�c�*�:�>���a:�D���&]�%�M�IK8Hip�Mf�V����aT�}m��\҈��R�8㍓؅��i~M�zt/����k����hmmb��dݹՏ��6��R����c�}x��Ct��#��bo/�'G�;؇��I�C%��^E=�R��9]Q�f8ЧyT���Z2XGV� �-�ai�j	���Rf$Mg���h�{Za疭c�t�K׮���,H����A�H���Waώ��'�8{�3��$���_C��3�i�|��::q��cƮv���TlkAe;Ӱ���E�R�*���@���lu����qU�P�K��,x�����`W}�����j��H~�O�f�+&�ᘂv�TꇕZ�)��.L���E�5�fP��_,��Ğ 4�������Hg���a2a�*>�z��/�/4�ꄡKDHIUqz���y��>�D/~�~�>^8�V%�	��+�H�C(h�����p(�x~9]b�����9|r�"U'`Je���g'�	3'��ڹ-�ٹ	�Bs>i(��y\9;A�Fď9���dqz��"�W���u�AY.�6���D(%�Df;�1�C�Gi-��voٌ�t�7�݂h�Ax59���ʍK��L�c�b�F���&E7=9��/��K����O|��oŒE��}�f<���;8���p{b�0X�n���X�2Iʓ`�CRRE�W��ǚm���G��
���O�բ%8�� V/_���V45�	Eޝ�!���K�sn�CtT�
�PHpݾ����3<���ز��پ��n d>���*��ꝛtf-x�P�T�s��F0jlC��E;5h��R�qd6eUB��a�%Z���߇��?J��X3����o�w^��W	���}K�t5��~��qp�oَ������I�y����52�_��U\軆��&��t.�$����mW��SN</1�6GK6�-�\��&<��y`j�MkVce�JZ��t>��>0D������s<�0I�h�&&�'`�e�}�F�ixd��W�L�:̒�dw��
qR�Ȱ !1�3�Yqq{˥���b�\.J���+Ō�о�U$\�l�%h�J,J��t������>ٻ>j]��n��X!U�pC���UÈ�K:9�4ms��)���Ӄ،�!�'�,�,uD��V�����	B�c��"	15����$�;}���}U�
9k�L�*jd(�MB,S�,�J�BS��)�_�i�����S.ݮ��<!(�t��'�l.�H����� @;�d1;Gd���E+�\��~�g#!�p�굅��x\���� �X3�ݢ�;v����m�V	��qdh��>=����Lv���y�i��xٕS�q)��&d�ӟ?��t�w�E�����˱�c)�l�M��	��՗q'5���Y@rd��XeG�.�@U���RpjWm�mR\~�Y)胻�aߎh����D}:��ǟ�����ӣ�$Ę8,��l^f�9A��q���$ &�O}8�fB��,Ǯ�p��8���G���k�����KS���I�s���D��>�T�Ps��sX��۲�����e���FL�vl������{�Bbv����eD�AX���L�M����y�W�#�Cch6��5�%A����d��Ӝ�� E�J:�Ґ��;�D9��U��5.�ܔ��q����`+/Á�`��M�����Iq����w08���7�>��X�J�Vޓ#�x���ok/�i,]�Wl�#;��r;q����3c��16�>v��m�*�˛`�U�9�aT\�g�T1�*c�}��]�~����vWV,1K�"��������Ul�{mŋP#d�MQ�+S�1R��-�=H���*KA���e�L+qk[I�
��z�J��2�$) veA����+_H����gåM��ڴ�\��N$�\�vj:�QPR̭����� \H=��R���1�3kV�'G�]n�G+2�e�$�8�&y(�gqX��S��
���N�rH���2�i&�@���ֶ*��K��tac^7�v.�#�û"+""��S�B�G>9�7��%�K!2��bh���業:w��F��:�H:���9����ȥSx�����Y�܁�?�4֭؀�x��p��E2Uu_hN+beh�k�UPe�rZ��<�z؆1�k �s�5x��/c3��\�Ϸ�]�S�x����滯!�N!ԅbB�.�U(FJ�]QR�gI��Iٝ9�9�i<�����JB�G�o�S_zWm�+o��?;J��m���ՠ��W�Pu�j2��ξ��8�a"_B�Ʋe�|�k����؝�*i��	ͷ>x/��r���+%IQ�ْ��d�Y	�1q<+.��R���$~���=��o�ޠp��Z�?����	���?�-.ܼw,�D.���y�k(���OՔ[��*[�-N,�I	.k�ēǗ�����b�Y2$S�Wo���I�n&m2�r2���O�"���+z�Hg��~�*���7��t�w��Ģ�.|��.��/�q�|򡌓���^�X��]��;w�kmz��f5eK� �UsW��T��&��0��VhZ/���!�Z�¥[(8�FE�����	"t�4tZ5u��|_��6w��	ȅ+YE	@�t)�s3FSO@_��c-乆"͖�R�r��S����+��[gA�����h>�~z��_���q�˩�%d��q�uQ5����>���sk!���E�**�v-�<c_!�)r|C�ͬ���u�P�Zz*7�a���M@f�W��$(�����u��o}�ݤ \$XmN��r�E\�p
ׯ]@��@GS[�<����
!Ivn��9�7Q� 䡋1��\�|�LNN`ߞ�ty"d�r{��������~������Y;+�&,-[����8��NzN�>P�٦Ҳ�����xt�~|��W��P3�p��+7.���q��e�&�h|ZcA4�7!=���!�K���٭�mQ̑UAVF�?F�3�Df
���1F&��c)��X��@�;��?�C�ޱ�/����ۄ�~�*�`7�}Y�ٖ��t�e*fPVݖ��aBg��'��b"�M�-�7���[�č��:� �z�������gV�U8�%DY���L}�� �J�W~���<L�<�
��>l�Y����3����׎} �Iil(�T�����	3��str_Lfĳ&�Z����_y����F��@2o�y��{������x}��loSE64�t2��n����7bbjqB�EZ�_��<���S�Z�/͓o]������M;��/�r�5d�K��"ʥ����K��8-0�+�厕k�}rV�+���� ��>r�t=@Y�:��]�!9���IjX�^�Cޠ"���ui�:
Y�ɇ��.*������V&��}Vlnq;�W�T[m�UdAK�W�����**7&�`��bD�y�,`3��[�,Xw_��tj��34c���:Cf�9t�Gł0��"i���&�eeB��\Z^�R�iii�g�q����������ښX袱U�>��29��n��l"a���~_%3��rEBK�"�;ro��&&F��h���V_���FBF6R3)L'���\��t��9y�B��s��֚K|n��>:�	��M�F��7��5�V���<�[�*��/?��|RRØ��hݦ�İ�h�a.�R3�I��P������_#AF:[B�^w��˄^_#a:���:S3!���ې�ț(0M���Otf�HJ����vs�M�������u����C$�W�,g7vm�NB+���o�+n� M�����^�T\�����pY�rI/�c���|h�.����A]�Q
`f�Y���Gx�臘�#��C,`����u�g�M�Z�f�]	�JP��\��d��&s3d�����ŅWQG�y�f�o	�:��?���?~��	9r�6>�>�3G���+��w�����Q�>��C;&3�/ ]�G��p��g8~�fg����Ѐ !ҩ���U����9����!D{�C@�}���$��'?�ν�c���떯��.��՛��މ��q��g(xX���g���X�P��^M~�Ӷ�!|qX���۵�_˃
��QS�V,+Yڂ�/d�h����?�w[:XfW���Z�9@>
r����SiPAB�(2M&�$�)Mfk���R�!M�
,D%��!!юj�1�r�Ň�Q��7S�ɉ0* ����WTTGe*%����>�Tn"��%<" M�� *n�Wk � �y呦��"�6+([�C'~��]����s�	A&#���@�w~�x�����;g����^zG�B{�E4�����Gc8"-���D�����ˉ��ȇ�6s.� L�^�J~B�a�����dr_��_�wܿ�~<��t>=�{���'�_�d*!�Y�d����R����RQBL�H���;��������9���Wq��5�G� c5������'15KJ;�	K.L�:By�� �H<���/{�����ۣ#��1<<�K/���G���O���潒~��~���7�:r&	si�c+wͼ�	�.�ݑ/�����O|��2|��	a^�zϿ�<.�^""
/W:�� )�EM��[��h�8+�������DI���RP���%EB"HVG�D��<���3�R���k8�{?��̳�0V"D���̇@�������(UcĲX^�Q��+Q:H*�ǀ�(%��~�7l��
y���8��k8{�s�=�t�@�HY�P�d�a�K��-	�Y05"3�-07G8���6�P�H
�K��'El`��H�>����J�<��4��w��������"�S!}˺�/�^�֩�3M�aAտ�Ȏ�e]��r�L,[h9�G�����Q):�٪������)V@ŵ��n�`;�l���T�^����P�L�2w��nS������.S*k�4�3�eS���[]ڌ����Tണ�N<W�]!BK3�U��Z�?�+�sЛPI���Z(�;X#`��g���t��Y��q����{����-�����JqRm-����"r���M�J�H�jP�>L�l�Ғ��OOz����,]�ׯ�_��ϟB}��b��no���X� �T2!��[6�BK}�ϟ��3�C���E�b1c.d�'�_���s1::��TϽ�s���/1=3����G=	�6l�ˑ�Ko����q�j��	���K6��n؂m��#�*b���'�᭣�b��IC8(9�A��%����c{%�]0����B�O�Kg�L\n��f(���t����]��3�<f�IL����~�;c�x`�twt��u~�������b >N�w�UUr��ڎ�G�2�h��a˪5X�l=2Y�3c������"��D[�\�B��$������Ȝ��n�����F�AO=Y'A!V�J���[�}p�S��L ��\
oy�^����=��0�L�nۃ��I���_b�0'y�0��7E� ���r�e�����cՒ��-͎���cx�Wh����Z?A� =�9֌�/H�����nC�?�K9t� ���VL��s�	�u��	5b�\`pyKx�͟���x����h�D���?������}����4;�]�����@�:.�*����>��]�oއ����^H_���)\Ј��:Rj)����cPBV�W�����2D�x=L�ͭ0rR���O�''��.�F����/� !؟aJA�x��WY��P�u��]��,����WS�Y�,9�/i"P�SY�Z��	�v�M�)��-]���\���I?��aB��pI�R*d-P�A9�R"��A��GY*\\����l:�,�D�Y�H�o��r�9�iIr�;�N5�̉��Жz�~���x��!����|�������~0�sO{V/�T��bA��²�=+�%�������
�������l߹�����&l$��9y�c�ę��Ǽq�6�?�G>>�㧏K��C>$���Y/�ʫ���tB|�rn�+���%8Y=@����k��@|&�����9���J&��+���K�C{C��!�VHd��/�~�$�#���J�Aʞe=���Jua������	�v]�׹�����t���M|r�c��U���-%S��G���^;�2k�����U2*�!�."/!Ff�nܿi!m?&F�x���q��c���x�d�5br�h&�b� �ˌ�3�}.+�������r~&Gȷ��W�.B�3���<�h���;�FV�DbN�7�q<��O�b��;��ص7�p��Ii,ɩ�FE�8`�;D���.	��׮��e��K��w����\9�Bq��1����Ҷ6���B�_����{Q#�'�$�MխĈ�M!�E�������$F�h=�m���%�	��|�*\�ҋ������}�7���{���׾�9R&��<~���b���]�_6� r���&�ei߬tfv�%�+��B;��N�BS�O��L��5BVi/����$�j}8`[�Apb0�{��[0�����ӥ
Z�����2��4��H���!�Q���V�	�"A��G���R��d>/M՘UK�Y���u���X�q82���E�┩��A���M,���tᴡ�;jlo�nC��K�=��ż8�͂�5pI�mUz4�S�#�)�n� ŲZ�2�9�����~��8}�m(� ��V"��PֽޅÖDr1R�ð��R)inS�ڹ��s?�y�q2�ct�ܸ~���_~DwP����MX�сB&/m�c��v��A�.��	:�	quHR6���Bo���ܪܥ9����7	U��ڵhM���ix��i�|�m$���;qkhs�sA)3�F|d=�O����R"N���8I&|����y�E:Gt�����$�`?	w�ҥd�^<Z���<�S�/G�GƦŧ�z��f��+<�'.�f%�֒7���Y�����G�C�ֶ��]"��/\ �>+V���35x��� ��*Rf��n@,Ҁ��7�'{�:3ID�B(�t<A@�$�tY����u��T(�8��:M�^��ŝB�
�ᣵ��R���el�rh�#��]�v�S��/��>���E
�O>�8��b8>D�-�J#D�f�<�t����ۼi����ч�g/���B��M�ҝh�o���6����P�J�x<�	�x_[[ŒP�Vn�KvW�������#5�&��G]c�#���۱��}�o����o=��ھ���}�w0M{w��yD.����tj����xLU�-*�Өp�Z��N�1�
JuL\[w�q5:����-O�&AE���B �%hK8�0S�*��Q��t���iTO�aYZN�q"����t[W�D���H(%Ix$�06���O籤�EZx{iӊt��&��d���C��u�A�n��J.i�h*
��UqI��S�z�[]�4&s�Q�aq~%�³@̑ ̊�u��A�n!є���B ��M0��+�$��"Y�2�oU��.{$���ׂ�' ���_ؚ���[ZY���C�`�����������v���cc��?�k�\'o����{�r�yFK[;�E1i}��H�3���Fe�|NaU)��T\~�mr<^&�b������c�0>5� ����V���m�=��y�a��|�LJ��S4��b�J��I'��;�ۂE�FF�z�:�\>�l.E���
hij@'	r�B�b1���bu����ɤŔ+��(N$��CBv.��1�E$��ǜӡ�LD����z�M��rsˠ׏�Am�p��O�)~�/clt�ǆ$gS|�P]F��rIK;��y=��I�����8��1z�׃663��"��,���x}�<�`��L:+��c\M'A:��RPư�G¦�-C:��3bA=�c'�''Es?�A^z�5qc�߹=����o|���lV��R���A!�%˰j�jIAZ�>��ֹ3t/��}�}XL���aoH�~p���?�,Z�.�������%��ꯉ�)A}��8�mۊ��.\8AJ�'����n$��͢�����ϣmQzZ��Js������č�Q��f7\ٮ2�Jꠥ �Z��jY�|T\�*���L3̅�/�"h*L��m�*�֬u�����s�辴���A�!-+�3d�v����{� 79#�X���`~6GՅ�]�c��p�9��|ɹM��n�w��|���҅`�.�_��006*��:��w�vl��WHUfɌ,ꨢ�S��� Y���18�N�ٍ�-i�kQ!�	�	�I�F�	�p�!2U��(m���j�̫���	2%�
��
�9����CڡR��]~���i_�"�,��>e~��ͪD1]� 8c�7��mB%�} �[Kg��T�ÿ��i����s,�9j��h"���Ԃ�a�-�ϸJ��y��ѥ	�fg�� lKJ�}� b�R=Ӥ�������x�Gp��U\�x�K���D�$e�����ކw�A��^���s���LB������_T׀-+�c����=q
'ϝ���4)@�;����"��&��r��B�i��++�Y@¡Ü�ܡ�P!IU	���B0G�v�^Ǽ��^;@�gN�6]�Ka�p�<!"Z�X$� )<�Tq���������}�,[ԉ|�������HO�J&�Wم�[va���`��|��||��BMa���l_Bc�a��m4��҉9L�NД����L�ˊ������jGV�M�-4~��qQ@�+GGF�l�hN�x��A�w�c\��bV��EK�A�ב�ݽ�~�q�C��Jl���gx�@�{��Үt��x��Op��<��$)Z��~kIv����
HL̢1JkJ��.$���uR3�z�a�0#��E+�u��"����S�@�ҥX�l��_�r}7o�$K��CssJf	7�J�������ϰ�!��͋��Ǿ��z�1����ɝ<,A�:��vʡ�%4횯�uIk��Q$hmW�!A~ܕ]P�'9~[;�$]ef;�D��@]����؇)Tx�R!�FnLh���c8�+Jd��"��3�3���K��ʌ��"m5��E:�f'�U�]OH(`q"w �z��KDX�����؉���s2n7r�'7Z��^c#����1L&R(�xS�LJ$���VN&S=�kS$���,!��iBG��L��/��Ҽ9������e�;��8Ahiݪ��^�S������B�ܸ���gy�38��i�Rq�F'���:�C՜;�^)x��a���渡{%�Gʇ�f�B�����̕ �/ ۣ$9���+�v7ã�#���EȊ��&����xB�
�᥈�0������9Z�H(��_B|r�N~��_ڏvRPsl㽏>�Ԯe]=ط�~����ŷ^W��$��MKW�G��?R�qB�l�N�ĥ���.������K����ut.� ��mAzY\�t�;W�~qv��X�.y��_��b��=LcL�$$��M>O�:%���Q�H�>�ю;��8y��e���AlY�����gΐ`+�\|t��.Y���ף>ڌ	,0�O���l)Қ���у�N���FB�y$�	�gfS���-]��dDI`�O�;B�d>y�2�[G���T2/	� 	j�?"{=x{@�����8����Yc��y��\�!ËC{��˸39Hg[sV�?&�>o�Wm�l��O��QB�3��`I�/nh@#�t�xI\bnMIȎ�p(F��K
��p��ΉW�X����FQt)�<f���%�y��-�ݸ���zlܰAZ�KW{iZ�/^�)�^Rz���%���o�ЀC�å�+x��di��'+p�Q�vM�� F}���?E�$�R�N�����U�yU�ڦDt�RQ���K%��6W��4u����gb�r�}A	]�ͣ��d�J�bJ.(3:�RE)!��׋P�
h.J�`�&S�b�4s<���M'�����k%Z��0Nf���|17\E[J�<��İW��I��f�y�Ȓ��O� �\SW��1�Еt�2������q$�,���h��O��^���}ŸD��n���8�����-r�������IP�>G�!4�ZE�u`�&%���𜜋Y�x
CQ�'������)��������ڣO!��1:=�O/�&%U �nc!�.&��w@�W�_$�1���p�-� �n�PE��j�*�(|v�"e�)B-dbӅf�Y2Os��QO?�^~�0��6ף��N!��	||�!�Eh��㉇���>�HrR�H[���-��a��m�y��s]�5=����܊��q�s�JZOva�1dַ�\Z1m���#VD�l9;O��։��@g�KȈ91�!>r��O������w���K���е|)Ŭd ���p��El޸KI ���� w��)�qR�sXҺ�<�-������������t�KB���֍'�:�"�.�Mc���عu+N�8.�z,Z�KWJ|�]Z7����Ĩ(�n��>d�0u��W�'���OI��pޛ�W����'F����0EJk29�[#C8������,·�x�ҏ1=7#e����5��c_AKk���9���	'�5��c��]O��OJ����A{c��Y��0|�������h^�E�7�|&)Ap����h�|��-����krb��c��v+h-�e��[7��k��$wmہx"��?|�,��ؾv+�Cux���S��`�4'V��4���=��,�����|	߃�p\ �X�V�Vk*r'�^���.�+~�NbK��\yϦ�A~���"l@s�a_D�:G��t9�ed��� M��FF&�Ȍ
�����Uk�`��D�v�5:9�CtY��$
.!�f��-��	Y��)B�,,	�L�佘!�%�GwK�Y�t�$��+�v�d��4�|�_0Ȇ���gHk,�b���#���ǐ��3��t�":K��A$�<�V�_H�r��<	�hSD����D�����N#��B�ۏKJ�+K'3}	S	m?����% P*q�����bhb��Z�$�;i��0=1-B�[~\�|U�<�;��J�˺'�Jh���
g40o)�y$h�oG.�%���%�[ D��3O��O��^u�-�@`r:AH�8:u��G���˖	����H�a7voނ��m���52u?"!�.����b��LD|��4m�4���)�e�Έ\bL~b	៴br� YM��T��Qd��Js��g�2��8`bof]��\���ML�`ZA�M��Hp���C?	�%�=��X���<��?'��-�7�aRA���&qⳓd1��;�����q�L�ׯc��U�ʣ����ӂb9�f��ho������,	gW�ٔ��
�s�rϙ���O��g�9ګ��%�\����]�"����!�����Շк�·b��-.�x��]x��w�#�̈ Lw�5�����������������#X���zV`||��<A
��Э��)٫��V2�W�}XA��� Y�C�b�Y�ӹ�8 [D����y`t_��J��z��ٚ��w/YJr����;�L�v`zv��I�.�q�{hUw7Y�q��)X\�� ���eּ�mx��|��I�� �i�"��2��y�Ǘ�L_U.�!uE��~���D.Ku�$�HR2W�0�t��x`�.,�X����t)2"Ӌ�;*9�����s�����.��T.E�@��÷/c��
]�BN��L��mn��"��	`�bѥX�z��gG�$� TK]H�0��%^(�$X������P-����/� �L���,H@�&a�cJ�٤�@���	�p%��l���Y�JoJ�\���qR<>a����p4�h]X����s���qә�0q�[]%��NK����6PvaזD01ʽI�ӥ+���qa����I��0r�B�0�@Y��㔮�
tZ*�&���*Ō���	
o��\H�"	�0w������߼A�҃=���O�cQc��1<1�>��w�o��8�]L/���Kh����Kh+���R\�/�ӟ)�|��c(F.�Y�*��<Ü�/
�M(N0�@��Ę}??;��(�0��N�+dr��T !�E%���O�:����}7��V+��|hoߺ�c�Nb��d���g�ŧ�!���}�>�D�ݏw�H�#��P=��-�t"N�ٌ'~C�#��z�j��~�0�S��t�D2���U֤������	K� ���Jd�|��m���Iy��%��%$�s�JaӲ58{���p�������a��?�s�����}��0�Ź���D��,����kFcK#�����PO���������a'	����}�=91�`\�B�1�p�4W�2C
����=��7����1ff1F�K{��~ϐRO�k{�m�FL����¥���҈����4��;d�ޘ^��us̚���?>L]��ڄ�zA���òe�L�'�c�z4:wl�H�[�*k��7���s��q!�U����}X���Ϟ�d|R̓��$2�9�m̑6fA���p}"$<�6_� n�^�1:��iuB9\v�hL��Yb����D����>sR��tQz����: ���%�a�,KJ:3-��Z_
��
]�b�+y��3�I�̝[� �O'�9:�ܶ�D�9C㟙��MjzR���a�o��##�]`rਭ�+H�pO/Ι�c�����ނ��7pm�OȰ9�M�Ĭf$n:Z�(�ݼ���v�z/�sq�t����P�gn9�e����)"�/Х�K&��As4��d�e���{Ŭ�=�?�Z7��I�%B�}7n��������e�Z�B�ٸd�����b�I�0�F]�B>k��E�l�
I7�>�(�X�[u��?��W�d�u%��o2#�Ϭ̪,oQ @ �!	$A�ˌ$��zM���gzz�׬5_�1k>fuO�FӔ�$RC#R") �U�{��{&#2ܛ�Ͻ/2���T�P���{�9����>��&��&�J��G"����+k�fS%7n�`(lԝ�V�33�9HV��wL�ù��8sr+�B �tK�8�oO_�A�٬D'Il`�8p�����A\�rQP�q�1$�pxx?Z��8~�6:L/-��wޔg��&(F�Q�{VW�do�O}Z�{	��\T�-��t�E���;���<�K'�N��ß��UL=S<���g
���Xz=-N=�?�֤��/�#��Ȯ��7���&����p��y\�vOH��� ў8�s.�ܥ��Td710؍��N1�-�;3�bkݲFSSZg��ʾ�A9�8�Ϳ�Z�)�c)����ܢ��67�Z�e��ۘ���d$�Js�I�q�#'O���~�SMXK��?�?��?ǩS�q��	�8(���aL��k�y�N��7}�7Hѫ3����Z����o�2��]#��A��BRP��8��1��Fִ��-�J���n*H��\Q�G�L=��'�h�+_�����4g9=5���%Td��s��^�!�C�k���DJ�X���skp�A6����mAbt�������J��v��-��Jmrt�-=��켆��`D�-��L�C5d=50��B	�3+��zf��jT�>����?L'WUmH�oOK�גQX�u���)�w��}(��������3R�|"&��U>�$�< �]�����a9��m�G��ٚ���wK�IђB��S�N�"F#C�ہ�X
9A!-��9�,ϐ���*���VYG�6�n��FfA��)((."���T����yc�RE[`�G��v� �ՂbZ�V�g��30����X�[������(R[�a�۲��D���T7����KdR@D�A��vA�-b�V�7�h�����ƴ��3-�0M$��,Z�a��qD�bI��;ǌѓ�ɏ��G���A%����+�56���U��T�D&�H��%
/f~�Y�Λ׮�1A|�bh�����.F&�c�/��z��)�͂Ҏޭyxw,�#�N�������1���zwn�ñm:�EU�R�
NV�4F�Jق�� h�G*��j]��w<���jT�z�\WF�e��>tv����C8{�F��ý۷��ѫNg��Ӛ8AJD��<'��;qw�$2�g'���i;UY�n��s�t��a9�F�*{`nzAMIL�E��ދ��vU �6�,�V�{�3�#3]:ڮ�T�n��5%F9/�ae"$v����ı]�q#�F��H�|V�?�S%�KYͻ��S��L>��j���h��j3 ���Q���Ӵ!��Vj�е�,|�1����!`�Ú���`��x52�
�&�
��<a��^��XR���n�(�#�[Z[䠵"*F��-�Q��NYߛ4�p&�������#�C�"a�䨈*iP�?(��p6��K���V��%Tkհ�.#媴#�f56�rpsb�z���_���̒��=*6�E��	ŢXʭ��|���r�I����c�d���}A.�l���D�]�C�{5�0'(g||B�SZǁ_����>���gf���K�*w��cO���],^=g�Ys����4π�tF���<���,�MadiS�W$����l6�퍍�1<lk��/U�Q���g����ƪ.��{�c4�)��9F,�t�f1�]��(��M�1������5A��|k	7�@<��g� s��MW���f��5�����J%4�~�g���=�\����V9�E�Rp�0��Q��.;Θb�Q;��9��AB�y�T���d{��_�L��!Ē�)�C�K� � �XxS�q^~�ŻO��iA{�*�}��-y~�GZ���c~a^+�Q���7��bX�@�8��:���uE�O=���'��������$}ŦiXa��yr<EL�艣��jŋ̴����t�+*�Y���AAñ��BH�$�����'?��W.i�ߚQ��a��9���w뵲�t��5�8�KH5��o�tL�=��gmz�Q�Q�TU�ͮig]Ti���Ҷmz0t4���}V� ֠k4_m!�A{O�\[6�95�6cX>gaqA#V� ?��Gq��-��9z\�5����G���� �@��f�_���d����~�O���v
� ��zz�[�
�%��t�ڻm;�����K�LSp�k�FD�)�1���;,�A��D\�rd�KSb�dA�KP3�s�s[U����R94�R�L��<o�ׯʁ�Թ^�.4�:H���c�6\~�}��&�,�����K�1\:9�O|�i,.�p��#(�Ɂ���.B��r�]�8�'��[o����P>�zB*�%R�T؞��q��'	6댣-��^^������J�2M{g;wi���+��n������(V�k�4<(db���f���y���5E7C]�8$�;~���z�0Ҁ�tW���ss�L.�S�R~�x��f�]���=���C��B0H�[V�;�;(��HF�K��zݝ���@�5v�C�?�n\�)�vG��c'�Ʌ9�S���cŨ������!A�3�:��9G,#g��Y���)�����cE='�H�Y�!�0!��5ܓ�ĵi�}�ܘ��6��8ʨj�yd�P-.,*���4+a���Hw��kJ$�J)L����Ȕp\ֹO��.���l{���k;��{��X$�3oݾ�Ǝi��L'��=j�&�#Ҽy�l�6�" �	���0��g���p2-�-�016&�ۋ��BoO�8�Qu�\㼬�7?;��aG����(�'F�6!�A�|��ǣXY�@A��O?�y�Y�|��EY6�4ɟ�e,�/h�K�S6���rYK�tk�'�;��T�N�WU��q��X]��"�����n8q�F�lp��+�$����4/Z��mp`�M�6*�˪6k�����Η��w~����x� #����zGô��o'U[���e{�.�#9F��	nnh��Q�"V���_a�d{3[Z��� �:��/hFB�� ��|�ܞ�ET^��.QP��3�g��L�7墚>֠x�*⭭>َw~�R��0��^`�#:v=���S8�³X)�07uO<pE�YF��
i��ʍ6
����f!�;����z�Z����������lmg������9��l�D�Q�i�؁�70��+l�mL5iVmYU.%�S�$�#^�|���+�hk�P��r���M	�����x��'y��R0�l��4g&���!��&�䘷$2st�-��c_ǹookE��(q�D-�"���kXYZ�A���O	�[�_Ķ���X*q��򓟿�)I	�'��`�n_�#�4f�:F��U��Ub��fP�=��.1"�F�\6�@=� QbX��r�l��uw�s"��2��T�|F	w����8!��6�S6���9�ۓ�b+C��8�eq��O�Q�
*F��{ �r���->rL��u��5SPd�ʂ>R�hH����AȎd��'�Nӱ��x�nU��Z3�|����k�U������g�V#;��������<��>aj���+"̀F������ݍ�;�)ۇkJ�O5=r\���5�+Ə��YY���u�;�,�h,�-�e�'T���iQ7(�!��P$�`�Ȝ#j*%�LH��Dw� +�{X��իה��Ԯ�K�ʩfV��H�����t?��7��,kF�A�}.�V�5��C�lCB��7�昚�D$��q�&�PUcݔ�����ȑF��H5!Vw��6d�g��5|V�� ��4�$�&�?���i�n9'�`Z>����`��U,�����/9W���4Ju.���5AX\��T�g�\a4����;��ֵ�h�x�%'gd���RY쑩9�r�e��-����!f<�Ķ��Ř�4K���*�׳�]uM޷AHC\ǻo����E��� "޻j%���vXɳ��r=�w�Gөb'E�s�}���� D
���{v�Ɗ�	洌PJX�w��ip�mp@ך�z�j�N���1AZ��r�Y�Z[S�P�	DQ�D J�������DGlItOt1'��{��-VulNE�Q*�#��St����.��&:ь ��Җ\k9~�:��V�Ibomm��X������v���L)}���%3�(��w�����(�:��fma��T+N�e�{Z�c�#m�F��n���h1EA�yGK�
:#o�~d�Y��f6���(�ΖO�x��]gW�2QwҶ\�Ú:�S19i�1����$2�}�޼qQ�k��#�m�[�F'N��k��D>�Իm��&q���V�����
!�ı�q��1��^A�}ؿoXSB���7���lmD�,VŐ�h�?d[�7$��c��kU�
y����
#���v�޻_�i�̦�^ȡ������}��g�TưD���Rۡ�]U�G0��"�P'��/_��~D����!����`&���E��|�SO�ҙ7>B}�r��4�3߇=�9]+v����&U{arJl�C3:;%���&�B[2Um�Qm�s���e�:b"l���L�,'m:�i��}���W��(�ܽ;��ƒ�^���g0%�PWT�s�8�Y+�9	���lxh�Vn�{j�<�x*��j���
d��G�ML�L`�7%�-�Y�)G-L�de�P����[�41:��m��aw�[���֭�܍�h��Fx���'�I�;H�M��ƃ�ȱ87'#/�q�]��ˋ׍NH�<#�^yM[k�CU+�\絥e�t��!x�C�j�r+�V�g{w'����2��J���{tcl�f8�]2�M"
h�F#H^jE-%H#���������%�Z� m�!�'S�f_;� QCg�zJB��Ck�EN&��[K�ixp]=b�%�>��̖v"�9�Q�7(k�N��u���K�9�`eeIܚ"��v��}nz�M�3�/�\(����+��g�61S���LH�=4,�]P�|�.\�r�l���1L�0u�˼�.q0���^'��C֍�~�H�� 0��I�פʲ'X�Sc��nPVŜ;/hϳg�"V��uj��=�S#\�\.��>*�Q���cG������ݺ��cL
6:{���p�c[+N�J�R8~���e�$Bu5�R�+�	NH�� M�9��y׈a�����̏h4�yYQG�[P����D7���yf� M�L�C$�&0�ajvVS"��gf���g3P8���Z3ەE��T�����Z[
�U.k^�iZu��+V�O�Y�.k�>(%���ܱ�i:�$��>bG�yY^�'�se14��Gp���8���Z���qS4IX2?;o���۬㴃��`Ŏ6:�U��Ż8*�uP���&�)(�j�PI,߷d{�3���Y68�0KY�S,���N�l���I`j��
y���sI�7̠R�ac.�F%���w��r|7�
���Y5��" ٌ�N�	4����@���ݠ����C:�� ��W����Q�k���Ȃ3���~S�����4����>.S�l�����!�����wiX�F�ݿ7�^GR��$Ԣ���:>>)(���;,��͹����s��kH&4,'M+&�'?�+.(ReH�.���!2Ԥ��Ɵ!}Z�pzsCy�a'����U,���.�7��/�C;���f1Ђ��&��WiœR���쌶ò�F��]�B&''ĉD��֪��X��*]G��{�_�������S�#�������d��SO>�9ErY�_�V��d�����3��M��i��KM;<�OC��U$Iun�*�LNjaҳbL����_�?tN�����r߰֜���ls�2|$k^��cd��C��?j�k����8�444Y�i�wM��X�d����[�n��_\�Q����QUw��ϓy]���D!�DJQ3�]�o�z�HL&�SD673�y��l�!F#Qtt�ɟN��+�eC~/��A��*ڱiI�c��˚8Z�G�y��H�A��H\Sd�E,�>�f���^���ܺi%6�X?Wπ���@p��ݶ-n�������F�쪙��#�Y��l 7�jM�n��UlH(��z��059�C���ы!����yP��q	e��S�� ;4X1�v� <mLx��)�xh�=l.O��3�"��i"p*F���y=�;� �5�\'V�3YѼ'�-GŔ٭W�Z�dAˈ6F���Ωl R�`�}�����O�>GP:��rFca��b�#ޔD@<t�^�Q�P
2�-��W�6k$c�s��Y�('*=���E��!d�Zѡ�;o�F�4USN+�e]�9<\��2�4H��J;��Ѹ�4����#�������%2���2ʎ�TF�����H�2	RMͺ)W�W01:*d�)q(�ul����B��c�d՜i�b��Ҷр���	�J�AS4��I+)(2��͜��������e2?��.�9EW�9PTћ�I�U+��T�@ѐ��4�!94M�j��0�Ïqԉ1����c��)�%�L�fYC]G#��\#Q����1���Ѩ�JyH��O63�W��'�i�f��;Nm3�9*�E3�_?�X_�v,C���xL�A�d���<��-m���2}����d4�87��!D��(g�+����3�8y-�1:�����'EóML��e���)s�TÚ�"`�Bc'D:��^���&"%�VMڃ�ڢF�!M�����-V	dhp�S^qzr�4�D�̳��Qg0�Z�Oذ_S�����p��Tn-���p�VY�?LǂQ�WDj��/��n+r�d����nV��j�P�@��gKs1X��^C��9\�z=-=޵W�/8Lb��"��b �F��z�b��I�XbXם޾q�K8���W���PT'�f�	�z����"�l ��?�C,�L{hF�e�,v1ɵ�͜�v�8�e5G6{4��������H	�	P�E��Ym&��ؕ©�	s�4�0�����wP��jkA�l��ZZ�uT�<s٬>�\�4���\��
|�Z�!'FvK��Z9�cH*�;���M��QwTB^#��h���"
��������$
Y��/�z6���{ M��вU4�#h���4���$7�,+fj�ڟT!#�^�"��D$S��7sy�w��%_R�.�$(�B���ю��dŉ�EU�Jx�fJ�<�B!��g�\J9T뛛����C����}�JԖI���k����b�.-�C-X|�j����ye�PʏT(?]���zUR����fs�ʀ���4K�٦��Ui��DU�YXXԢ[��zɾ���V6�C��*
�,-.
���޽Q<��bDbA1��&�y�SN	��Ю;��-?�yqD��ł��G���\?�4�[X�PH�H������,k��{+j�A��-j�e�)B�Dw�eV��'"{�p�Seg�;(���5�G0u�6����Ygx��+�iO[Y��Ut��BNv2QTD�k,睼qW�Y�D��ig�BV�ޔE��#�!J'FCL����f���|aUӑ�o4�%C��X�0�C뾰��ikA� ^U:&�,��f���Ng���7�X��_�r�H�}m����?g'��[q"&zӲ��A�;�w�]��a#�oC؂ ��T�Չ�)L���vAc2����Jg���A�����haK�x�d�������w��ǟ�؛?��(�+��,a;�3�g�����[�0��YF!A�A,��3�����b�X���xeq
^X�U��X�����L�g�[Og9�^6��]C{q�ģr����r�tζZ�WN���j	�K���6Q��ء9'�b
|�QN �EbT��n Ƕ�xyy��-�88Ҟ+=PD�e��`~�O���eU��gμ&�l�EԦ]{��N��G��DC������T=��}�H���:f���DB�:P���'?�dK���g$R��w]�!��`��Bل˫K��d�hj����-�9QS1h�D���Kv8%y�$�id�A�YJRKH��P�Ё�8v䰦�VE_�qK�2y�V�F(`Q���r/aq5�5���Se+5B����E����#��$�`�i.�JE�A�F�C 5��L6���Mi0���<b���Y�wu�W)HD�ҥ�>��T��-}�d鄢!wu���Ĵ##�#v�b�D(YYCrdW�PƓ)
�i�dX,�h�I1TT��m�Z�Ø�l�R�D�d��,.�be}��XF��6��!��BZD��4Y(�}��_����4~��)ڑ�ѱ%e{mJ�>SVLQ�&�I}�ܛ�\�6aֵyҀ�DBm4�ca~�g��JI,��H\�E�E}��}��v�Y��>��h��j3aS�N���e��(\Ơ����|9��oB�֥<�=������Fo��\6�*'Jf7�K�B� �"0���Ǽ5�U}豎� 5�ng�	ZI�Aa�eI���Z=�:��54�ܝ�r #:�ӣ4��*| �Eҏ�����������4!���򕫶Pc��-�÷������1�)j��ϛ�����W�{�|#Fe�v�ЋjSq����,�5����ʅ�
N^7z(��j\	lf���V$t+�njFj !�V��z!/��E/φ����ʁܐ��.���3�E,O6���4:[:�M�����(a[ދaQ��=rй��<�t�fgg�07�m�͂��Mx
�xn=�Fڍ����6���������X�Ѻ���=��(�1Ϝ����}�$����f�lWB0)Ws��)�,�,봂�����T�1ǑgJDg_o~�Q�����;��ޝ���u
�Ya����)e�oy���Mr0S��Ǔ*�^�7���u���`iyQ7L��1e�y�`P�>�"~����<���(ttu��[�*Sղ��8=�[�4���,Ƥŧ>�i�<b�Y�b�'�&%2)Yc�5q8;Ӗ�gn�Z�zI��v��7���^7Z�l𡴥�OZ��TB��2D<3�^���J��*�0��ᓝ�?w���ռuy��ū͍u5��+4� 
�[�����)����^�g	���er�ᘉ��o���X�^���(ȭ͘1_\���m��=�f
��NP�	PS��C��c��7�6;`�<|�[$� u�3�hݑ:�$���꒼5�o?ͫ7�;�c�k׈YT,�]�Tt�!OS0�־��P\��k���!1�-���d�Ġ�.	��r�xh�DC�������\	ݔ\#퇟4"l��ܙ_D\¿%��p����x零	��O䣡��l G�<��/e�R	���51��*a{�YDc���g?��W��(�7բIzv��O����KJ�v��Hcʅ�� )G��⩚7F$�����`�H@E�s��se����@�)p� i��F���F��.�Q^�i���tt[j�i3e˫��C$C��]��Ě����9��{�)U��L2���ïhs�<Ф�0,����cc�@3�WCOZ����{;�Ko`uqA�&���,�U�9��9�C,b4+��b�<�rh�?w��bxp�8ҐR�x�%Ax��o�5a����12>%�,��N,�4���"@Mw��<���c��MC	�_چ3J��������r>�,�ș�����TJY�	A���D��G.	�"���*_[j\f���5��f����R�mhikUg�٥�9�lQ�4���7:���z��9�]����>q�$�We��D��x$�kHcX�2��Y��n�D$b���?\�xԬ����(�s�����(vaF����<�5�ca�$٘ԳO�#���vCC���1׋Ə���)����s�}}���3i���t�YH���[R��
 �/b��gp��v4��L��j��	�/?ZoX}MX[��Ӯ�Cɚږc��|�	�:�2;삺bWM����T.d�ϻZJ��wu�g�u^B����0C�϶ AU�֓t�$�I2���H�ڔ��O̅��VPzC9���5,d�p}~L7�4���b1���*���h���<���Wϫ��]$LaC)Pv��6R(SPg�n�[٬*^����Xmp���W~�-���OB�'!�����8�Wj>$0�!�*�-� ��	�HX(���
���qtv�_T_�j�Il�A\d�Ԫ��~A��_�C$�ҍ+8,H3N.����f $�UcrP��:�jC�C����E�;e�rcm*�.a+�SC��h��������=��r:�gtlW.]�����E�=�P�����~-G�L�Qikm�'>�">����c�S�~���)t�`x�\�{UהHkfaFյ�\F�)���Ѯb-�t�氪s�ȿ��'$d����i0�
�_8�^�&�i�7�jo���bT���{�E��}%���"_sbb\�Z�b��s�ڦLJ^L�^�Ա�:��֙����gd	Y�%JZ��M�c��9t�����c�Y7Aҝ
�hWT׀ΐўg9���hV�}@�{��Xu)$�8�w��F�0[�j�6g�Z[ZZ����٩��ajz
�}����z�m�CA5���1yV
:�Q�x��)���9���F��-�+Ӄ Eօi(��Q搓k#Jg��l`׀^�8Lq0��(PUGE0�b�(%��-���t�[Q�k*:�_{�ԋ�9�j�|�Xml&	BL��qM*�-��``GK�t`DQ�?��a���?�0N}����ja�5ήc���5��Z�I҂43�خI(�2�%A�ƅ��)0צBjʗ�n�\}?�K阎3�;��U����f�-ÿ�,�ge�L�̜τ*1Y1I~�?����fv�g�l5��nR��7���L�4ED��"E#�|�S�%_�##� V	!�9�ۂԱ�xj�6�g��}���"��������?�D�	�>�4~��+ؐ�y���ڽ'�g�<��_�~��uܽ{O�a҆�1�b<��FTy�Fʱl��jlä'�q��Qݰ�##�_^V�9�2� ���LAL��c׮]��X���K��1"T�b����⭷��`�6������Pg� �'IB��ДE�������K�/c��~	÷��믡 6�2�D�t;�a��2|��R�amcM'�F9������̊r�Y�Q��:t�"��T�"v��ۣw�	}��q��w����x��9M뜻x/<���(ޔНU	"gy�۷nj?>?k��A�T�jhj�������\���kOs��fxv�^E�[�sb`�ݹ�{1"jR�����U�����{z�a�xHևF������f$"�%��蛼gA"�[��`߁��Ȅ\����0��t0���*P��'�K��5Ȥ3��0�����r��Hoe�����t�pԤ~xX(��(G��i�)ۧO�<��O�Td�%rB�@�9��AJ[@IU��ʖ���5����exuF���\5�Xnp��R�*L���)>hh�_��s�>]��`�vU��_��6ݴ����)�Nͨ�� _I큢I�W|���MY,��͗�`�� ٧�p/#`���c&V�$�]ߟ�q�ldp������� L�ϴ����am&w��%�V���LB%/滪V��(�0��"�gϟ�a�������Y��I��X��c��c[�� �Ÿ��s�\]��[W��n��/�ԡv��.J����6ŀ�1���Z9dEGu�RH�+Fc�����k!"e�X�)�.��-��bKPs�}�p��Ax�����C-���X:L ��ݚ�.*�`R����BY�l�>eqB��IF�Z0�,dD'E����|��f�n����+m!��4��Q4J����V���u�8��k||\[yc��/�=�k��c��a��TA�4�\���U�<�m��1#�8������]Z^����i#AK�A����F�����q<&��\�k������o�^]�1�g�(ly}덷4�MU���5-~�*��4���՝�t����9[��n�RCh"�R~�(α�O��{��w�"*�oais���5�Ԟ��,�������DƉ�&FƱgz��8�;���Р}4Z������J�(ƞ�ڲm�(�4S:��s$��) �����i��Q*���{�iK�d�I{dC��m%�/�c)왱vK�"����l��A��m�����YdƐ�޳�8[ �$�\]��;����6�����*cNK�3�|4�Xzm�oF��>L�	�75.�d��/�M
"hnV����c���@Bm�U��G��l>T���݀�Wf��3��j��E���N����3���)�~�����6�1�BCV$��i����ҩ���A�}���
��ڼ�ks�N� �MO�΍�7�O#.ޞ)���b(˸r��	���8`�*�^ryض�Mz��/I���&���>9���@-����Ɔi��(�h�ac��I���}D'Y�m�u@n��4$�3�����l��_�K�99=��5�;�{`�o�������	�?�0��uh�xnvA�3�d_	��[U�w�,����j�m3�sf>A�yZҶ��%mq~fJ�K�DJ=�-:~;kTܤ��n
�L�1�w����{��.({#�)d(��a��o�#�b��ﾃ��U}/��Q�$�UE��*�5�~�t������mw�
Ce��<��΃�) S*(R,���a���+)����b\9���I���;Y9T#H��tnw��U���ގ��A���U�����3ￏD8���%�>��
z�#'��ld�ư|�l҉��E�ժDM�\�\����Z�kς/�[��L%��NG �S���u	Ũ�:TrjzL���4½.�C]b�%`�j4=c`=nx.�(�էf��D}��Wͽzv���(*���F�{�>�U�q�c;���3τ�~᫖k��6�G�XU�����8t:��V�=�O.�	f�P��П�4B�7� E�[����m]4T�G]��|n̢y6�'�u�"]դv8�����Ni+������'���[�#(�O�8U?ש9��-g��}�����	�S8t|Y����N����*�[^����C�O"i��>�"^�� �M,o�blv��-���Vu4EC#ċ�)�rH�bۗ�!d[rT0�����;jH�&x�l-�>�@2�c9��Ϸ�o@��l�
�=sJ��,�.�xN~Xˈ�lK��rgǦ���������Yt
R������HA�D«���M���M��6��8���v��T?�.�4�Y1N,Tiq.��K��i��ŢYȨ���O�xƖW�J�oD�D��?���1�2A�72>��diH�׳���f�JK�e4,&!�Ʊ����w�Ʋ��#b�:��)������K��S�K�4��9B��G�j�]dE��֔���M�n�ҌT�T�v1>3���G��ϡ�Н��hxajａ]��qx�A��������v���hYmDcsڛ�06DIP)e:��#E̮/"%�9R=,No
��JU��"I������e��r�
�d���i8��'bߴ��L��,p>ׇ���8r���j����a��u�̎�g�[�Ж<��L���v=U^ �(a��Y���:��Z���L>�v #lA:�VL�Ts� �کu��Ր�1� +tM�R���yG�f�k�LmF��z��(����m���v�UZ��SQM�� <6g�P�^$�V�F����ذY����@|P>��7F*�k�~K.���_�3���J;&�=�d6�m;���ǃ_�5�~>�7���x6^�Q��z���Yڌ��3׿M$��G�Ù+��{��2�
Yt�q�n���ZA'�.�-"$Ϋ%�@��lU�2">t&�@U�ޜL��`��LM������ˤ�����Bխ�:�<��]Cp#1�;��?�(b+SPq���%5��{w�{Dؼ%vI[-�lJȼU̡7¾�!	�GqwyB|Y�K��VS����(��g�#��C9Y�خ<}H�gS���;G0Q�
�˿�:��*��q2򝕅9�S8{�
�&��%!,�yLc����p�Y7'F�!�W�r_�R�Ǯ|':[�tl��Љ�9�.L��JO�#���"l^	��N��y��Q��5��jN� /?��7VhJ�dʔc�Iv�,Z:V��1ȍ�Y����V��И��&����]u���ЕmV��p?a17�U*�Q艍�
�W����E`���|I�%����6�)��(�
Y�0mj�}���͕�|y�����9udu2frE������X�	����ò���M� �
#��c�(%:���2'��:���V���ϳQb�����k��NNְLT�M���kq��xf|�9�;ů��j�=�v�������N+Y����_p�p��v�����f��q{յ�T� ��h��������*��F�W��s���՗�ޭI��R�^�����u~�W����W_�?��o����g��-���������l�����ŴF��j�{��3K�b���=���F��羈�}篰&ޝF�-�R�O� �����=p�lb_	����i����Dt:�T]�=jv�ҥ˂(���مCG��!~��WpE�ݼ A��y���YܛEW[+���U������:�f)��������´�{oNjuz3���(`��,�-�X[�d�����lGu�m�	1�A�BCNb=s��*UՎ���dU9L�kv�����X$��ۘ�-p�� �t6��9DyAQ�g��xp�>㾸�&a��<W3&��eХ|�CG�aqe�x��E��V�H�(,�[:z�mH��&i�R)�Zh�4�Z�e�]���3�S�0HJ�O�;�ƙ�(m��Uz���'�?d=evw���ynq	�*4�������H:Շ�13��S76�򶱲����{њj��ǔ8���T&e��r�3� ��Z3b��6�룴%���-���M�� іL����w��P\Z��Mɨ�,J����O Mj���g�㿠Q��+�Xd[����Ӡ�O�d	ktZ�H����?}�cs�~ܱ6�O��~#[�W��c;<��tme�7���s}�|_�5If�w�b�������J�+_V��r/�F/��>@�����ש�Y���/�S����3�T�M/�����3�6$�������g���{����e�s�{����Z,���<������𢡄r"��=��������IgT�-�"�уH�I���c�ib\{P]�][��l�c7��ɦ݈�bX��Ez#-����ն�����v��9a�A�𥈃�9讄χ���_KQ��<6�[@,������55I|��0�2��W/��an��o�r Ux��UU�hy�:� �c��@��cw���k��]\DI�t-��������*�����6�ah>v}}�v�CW{��M��.!�v���@�L7m!���?��ߺ�����RH>�G5_����٨s��*����UuDP��`�6�f e�
{Z �����m�]*֜	��
ח�nc�#*�rh����+G��Ԥ8�--�-������GO`����ø=vy���s�Z�^^�ݑ4��!�F�*jyaQ��m�7�+6����Ց�<�l�`���,�Rs�*Gi#)~/o�<��R!L.M�ڵ+��F[��w�&?s�<r��!Os�&�i��W�@U�JY�6�X��4�S���"�������S����_ٱEjN;��A5X��<";�j��Θy��׺�u?7t*��pO���!��͟O��A��P�ը��U1H�G�N=�����8�^�~ԩ�+�b
0Csվ����zP���A���[��_�y�=|1��`d�˽�g飿Ϩ��_���7d)����(���w?�%4����翂	�.O��|zM�Q"
��3��%��aFxF[45��Z��#X�fH!_:+�f�r�U%�=zDf�/�ǂ���V���@��Q� � o�.���8��0��۱���� ��RVS�=�V҉�Y��|��Ǿ=C��'_���4��@�.��1:�O<�,�b�����$�]N&�o*Y^�78FR�*g�d����P����;�x�hH��Z���G�/�~Yͤu�dJ�5�X��4�w�C�<"(�k�S��{&w#�y��f�&h��]��x������X㨚XLXJ�/,S�  S�IDAT���ͷ��g\rTH�����Lqة�2���9fj���?QX�ILH�C�U���23�� �g{�X�,�`\�-��s8`Z����$��u�`�|�c*�����[�u.���эFJrJ�@����G�37�	�ʊ�Ӵ5H�Q�ye"s�T-K'�G^.�`���T�!z
�PՋ���(��fO>�<���q��{ʣ/��t�X��^Yu1*��.SN4�|C
�ƈ���:�8�H5���um͵�A�������~;�/~@ŧ/XZ�^ygc:V�_�`��2MSZi��-�i,�F��Z����Z�L�u*�I�J�����p��=*~a���0�`�joǲ��1���ͳ�;�ў�Z~�7�Z~�7}i����tj���7�5{�N�M���3~��?�s��j�E��.���������'���=�C��������&����0uxhђ���hXS*:^.�o(���Ϊu,zJo��!-U��^ ��hii�R
�s����r��v�RŲ��U�����ѓx�'��ݏ��37�`bu�P��b`����Źk��_D_������_�|�{�����!_���H�����ަ{i���+�s�U��rT�3�םc�� 8]!`�*�,�Sk�Is��l�<��G�*�bS�qd��MA�0{ԡb������(�|�)m���/��-�So+��l�H,�m1v��Xn�o��*�� ij.��kS�ډ���b�͕����3d!X��j"#�PCL��)�H����x��g��ԆiY��o �Q	��g@Ԋ8��W���ǟD��O��"Ff'���oj޳-�@�rd��eR�p��*�(6�h�4��8�P�(���]x~�õ]x�����������Iq�R���~��G<�����Wϼ���M����m�S��0���L�0�Og�5N�rh)�S;y��/`�{5�W{T���Z��;5����55s�Jq��q�_��Y�L�y�c���e�O�6�AP��~/�Շ�NM
M�zצoM���m㘰B��lnӳ:
�o����TT�l�#��V�7P~���}����r�kl��A�c}lk����n��k�Ӛ���ACoG����I�F1_���������&�<t�����XO��^e
�=�ԓ/���k� �7D�!1"�t�5�P'�ϲj�ZHY4��K�>U��Ȧg&����MkgSϮ��.���{{��Y12�w�O�{o]G R㮵I�t��eM6W�֙S8����>��Z������e�/�a��� Fd��[S�Ӎ��P3����V�y���	�l�3�EfZ+���Y��5�P!�|i[߻���%toK���?�ށ!q~��O127e�N���X��}x��5�z�}�i�E��ǿ�G����w }��7�����{i������H
���Y���uO͎t}�Ϧ��OY��=�x�'�g1;+{��_��o��K."��O.�����2,�Ʈ���k����k）�y�Kh�����;�=�r�&��S:sh`�ݸ��Ξ��?����K�A�>�%�c�{F�}�c緋���&���x�\�#�Ke�Du���tv�������#�U$� 덷_���JayO�A	��� �;����Xv���fR��h�9&�`��1��S�p�6�r�ն� M�~�:��⾜,�T4JoR)���!e�F����@e�|�a��1�!m�3�_�$*�;;B���McMK��S�W�Ö������P�l�@"�;Ƨ�W�Q�Q?���+����Mh�����P�˫��C��,�~d{��|�3������۫{m-���ג��G4�;#�_�1~�S_DSC#^~�E�]��o��x����i�3[�N��B&S�nft�65x� 6�l��l%��rXc��r��HS�<���Q@��Mb�b�8?3�c���/��A(ތc��֏~$(�@��}���#K� ��͟c�� ^z����A�쳟@wk;��7�&hl��^=ê����5�I���V����� �`�\Y~����e�&���$_(��8���UqJ�H5'5�������<���ڵU���n�s~E%/��W$��#�ۉ7V���~[~w��Eok���m�;u���ލ�b	��9l�ªN�&4BȄ�t�%�ɏ;*8�ۥ�M�����|\��;��R�������7����/`@�ɋ$���O~��{��6�BS�!�����F���x��c�78��������u8��T�8k��Ņ9�#N��O�c�=551�c�(HΜ�W(*/���vp>7uzjXLJ�Βч_�f	�uݸf�xk|�}�8r��<�(�b~)�⇿|YW�W�P�L��*u��3�pDS�kЫ�к�s�2	j��>��Ca�x��S�ɔ��q�����z�6#8�1�I]wGy����6�k�1�������Z�NH�D����4]���F��4�Q��ر��Z7�mT�R�$�a{�����\�^s��N��O#[�~�֣Jc��{�n`ڃF��%<�U{�Wo"�����|�}O�B���L�7����|��~�F�~��;�p�� *(+�{���C�����A�/<����[!!�8.߾���ݪRU�ʣ��	QꢺF`�tVUz�mH�n�YW��i�!���E	�gfTm��������i<r�!|��>��C���%TO�Go��	�Y��L���b�ڲX�|^�\�׿�m4�;��#Oʽ����GLF��_����+�)`O�G�(d�
�YN~u��^C*��	�W�` ���ek�|���6�������f4��*���ݏ�����H��������B�~�u���Tm"}K�bfc������=m��hnǿ��Cs��tN�a�cniE{G0:2�d�It���-I���:�=o6�k�&5F�":-lf�4$p��%�8~�~�+_���K�������[nE�I��Xcg��gK� �|����=��9��{�����ox8+h�;������E��}��طw�ʟ�Dk�<˓����*�/1�쫡*JA�a�,e$�9��fbk�Af%9*gtjR�?xPl��:�g�]�����KI�VUk@�ju^�Sw�!�PR�\a�Y�k�|�v��Hh�X�l�ô�u
���i@���)�,4lV�����F��8>9�t���c�S�*��&�I��
��(g��#i��۶��4 }_h��N���d�3�b�B�
��0|H.����+U�$o�֖-��|�����Qq9��U�U��Z��|#Q�����!藭`���������ߨ�]s����Ϳ��Sg0����>!�ܟ��/��Z����V-�S]�j8���&����D��8����<q�Ch��$���Ĺ�gq��-ݤÂl�9e ��Um
�4r��Nw����ֆ)򹄂�h!�Q6~��G��G[g��ᦠ@��?��'��3/`�{@n/��|��������Q�@'���?��7����=�O�/���눛�GO謭�O�?������wpw��rj��߇8�e]L�{F�QDq�/Ķ�*M�G�'%��N����J:�-J����&�E���C'��Sϣ��W�AS����o~C�4�N^���Z��݇�)r��U9�.޾}�������c�+�����7�3����믿���Q�+��`Q�'EStD'�F̔ �e�L�5۵U�Č#"י��R���h4��2����~O|�)��Ƶ��������Ť8ȼ ?'�Y1k�rS�d+�e1~���[?�����:��ػk����;�����[o X���Z�B:�C�8���˴�io/������m��耔]N))�1� ��Q��m��׊�56*N3�b��NX�-�7Ͼ�o��
���c�l�A�ac09�đh�c�Kh��(��!�����0�r=t��#:>JLŬ
bS�r=yF����B}�{�)΢>����$�$��Z�.�E����C�<a=�tբ�bSVٰ���|X��7n9Ivɯp�}$�R���@z���ʴlP���o�f,G�a�6{�iˊv�s��0�\Bu��x�Ns�'��ir���9>��L��qw� d���ҳ����}� ���o ���-Z~ �GML�7�}�}��D ��B��o/O���������ٓOho�C������/>���NcvlM]x�䣸{�֖V��S5��`D�AM�¶����u�����-ETI�qΥ:�'�xR�aW66BX�e�_�����_ �tF��b��>���ԕ���<��7�+���KA�'9�O<��^�{�=���[X�YA���ʘ(p�a&���]jq9����Z�<���[���E�m��[P��#��+7��N�sٿ�0�<�F�g���/p��e�Beq^!m��a3<q?wjS^D�ˊ���_|W;����-�Z�I|�˿������ϱ�2'�˕��Wű��2w%��dt
�@o/6�4��X�����Ġ�Z�R&S߈ ���%��=��GRyΊ������(��U��FCW��TM����-�,k��7/������Йl�Po?���k�����4޿rǏDGG�MM�s`��#j����0�|	ꈼ�]�mhZ���SI�ӱ�E|L"�t&�����i(Tۻp�&��Ə1�^@!X�n�PD� %8J\cP��G!rY�8u�#�%�n����`c����{W5TJ�l9i�R�Vri��/����I�#'Z_�L�Sq�tD�6u�vГ�����Z(B4�f<���X��U���Bj�$J�&3U�G;1�Ӆ�T+R�(��!���� }%'�kikc�Leװ��u	�2l���T!�Z*��8nY=[U�[1�5�}�,�7{ۈ���異Su-[Z�+��W���_G�}קo<X����W�;G����HL:��_��k��Ʃx�0?�t2������aia/=�q�T�p��g_ĉ}�0>2���1���i�55kΪ���wj�:�B(�L9?���Am��{�n�P�Ι�0�?��?~P[6�w�EK�EKa��ɥE|����O�}]�����5:"���3�����UG%����$��_�?��O}	/~�9qa��B_O/^x����cZB��մ�Rklf[eI��ᐉ�6�6Q�Hw�}#mH�7�`5���!��u'�?�S-����jB�	Q]Q�[7��}�]C9^��1v��ı.y�j�֖��5p�{:X�k�Q���/�6��;U��#~���\�tV�7��el�3j�ʥe��-	�fȝ�z�v.V�	R���M�Ȭ�q0�|�3��̦��jjH)�$��������.M�B!$F-$O��jځ�+����U�T6�t�϶d����ϔ�/>�����qa��g����~����d-�QΖpb�A�v���WU�%&�E\��+�I5�I�@[8��VN�͋��mo� ΞET�=�^�Rͪ˻%����g���I䶂<�V������$M�iE�SZ�mM1ٻb�;�k߅�p
=�mH��"Q��k��K��&:�
dEW�[��o�� �����א���#����T\N�`��#��(\6kY��N��Q�g��m��T��������D�p�78�;�=-]�6�)��Ƣ��T��x�lE[�p��{z�X����2���Yټa�����f�<Y*�l��[�����W�}�_l�v��]mzݳ�sv�:ne͸=` lF���+�������7464x�[oE�;�٫q[��ǘ�������W�������/����#"n�wz{�=��aj|a��r0G��T����-�V5��FZL��h��m��j�~�g�{ϰ́�y�~g�˳�������e��H����PX��+
��xە�)l|}_��_+{�^���-A:r8�z���=�C�O���]ܹsK'@���ؽF&D��L��*��/��?�Fvt|\�n�Q˶���2���]7��ë���x�r���|�V��c�+�������6�nӂ<+:�37/"'φ�v�oH6W��8��:�rYP���.#%מH&4�^^]Ո0��A��/9�M�:�:�h5�����sOah�^&!��Ģ(�=�_�����?���]� �:��$�+�L�A3D���0�Mc�ܶR��<RŏO����?�wd`Bb>��c8|� ���aanN��:;{��E����gW9]b���� ��FX:��%u�d$��98�q�L��X4�ϔzɿ�t�
�ݜGI���D
1�D�4�Q���\�D[9�&�i�ކ�Drh���M�#k�����Lqjz=`r�q!r�B��܀��v�l.���=\��bY>#2@T�O)`N~�[_��y��E��7`$R<��W�l��ll���oAk%��h+�ۏ��{�;�+�F���M������l�̬ؠx��X34v���s#8-~+����Uےk�����=e2h7ϾHve���Ϭ�b�����G���L~=hd������ox�}F��ۿBY0(���w��%�C����f[*z��a`�+��;�0�8��=�)<���r@�e��l�Ǟ@����Ξ�	��0�xD5-V�ٳ��dx�M���ցT{����=�nհD6%�z�6^{�m���)l���b�"%e�hޏ�р���=�W����6�/ߙ/��W?�..���������� ���".��?�z�����*J5ڑ�ca~.���zZ[�����)	��9t��i�F^,OG�
R˫��+��'l�0���mM��V	�� '�Q�?!ʵ5\��ʟ�W��ƌ8�e�"Ab�N��#��1���v�=}
3ӓp�1�O�<����N"��x\YcCR	�caJ䩧�C�����FA���̣�x��Y��/_ǜD���(k%�z��Ҭ\�V�
��d�rp�L2�!�{�"fĘ~����G�B��	��vkF�hY%Ϟ;��A��4����X���6�Jb��51E��:	�eM>��'UT��*UOE�Y�������㽻�VJ���TW6B)Q�}�Cej ����r����L�Â^;���hooQ���&�
 Q��m}��5`�D�b��
[���D�L�m&�S�c��K�GZ� ����Dl�Q�j�y5D�oGĚ�b7t%��j'���އ���W�kB=i��43oȼ��Up�(G�3)�������܄��n�z��.�cUB���<P2m����Nӄ��m�@i���P7�
�����3��1��ڑ0{���W����������;\<���q�s�~��GL��8\3V��(�M"��Z�w^�!F&���C���`� �hQ"�)�3����F%�
k�(����0��[7��ÂXN>�%4Wz���0*ɩ���w�����0�4o�U�3U�AEY&a��oZL� J�T��������[8���:�a<v�am_e=<<���W����LfK�]�K˪��� ���Q�����a��}x�gŀ���XA�����{��x��{c�J��*�3t$e���+������������oh�	T�˻���_��K7�L��O|O>����dR�-����̙S�{���(��h���TBg������1�o?��8����=�9/��(bs��%����0����J�qF�E��L�-���Z\U��Y�:���/�Sl}��;_WJ�g_�4�t�#���b'8C��._��A��R�+kX[_Wu1vxQ;#ݔB��}�߲=��?�2�F���ϯ,����\����w��n���W=��$Q�+�'m��#�R�cMx~�z�D2Ԁ��A�c	�Vߧ~ڂ�]]���t�y����/o���;�����Y��EQ\D�T�ݴ,Yv�r;����#�*��S��R�T*���q�؉%��bʒ(R�D
 $@��`�����{���~3 �3��������j�,�؃�Y|�k��}��y�l0��O�HW��Ը��֪��;��}L�l�U9Zv����|�K���Qϡ��*Y!.F�PDT}wl�B�*%@~�tLϫ��햰��o{ժ?��>��2���$V�3��9��(�UI��eE/n<���7�LM)�s���P����b>�	=�y[�x��Iw��`-���#�R	�I�sמ��6�����7��g���o|���/�HhQN����?��7ހo�巸b�xV�d�H��y��?����W_����7�ܥw�������:��o�]�� z��D\])���MC	w�e��Y0R�Ip�����]�������s������S���g�'������_�x�W��ٟx�5+4q�n#�om��������WU�ǻp����r޸pΏ�pu��E/���x8��ab�mK�j�<�LV/�&�L\��a?����5� �G��_�����~�~�x�s/§N`��"��[/C{mΝ;\� �NEIS��x!	.u��_�*<�%z*W� b���D��o���Y��q�^�F,�	�
�����ʞ٩+Ä�q�lV���@�3a"K^�����_��y�������8v�(���#�����'p��wa��	h��y�0�:�nl��˿�����^����^�.|����y/���O�꽛0D:�G/F)u|���z-l���������L�_��s��SЫ�p��1� ��hQ��e�Y.��L5��N�`Ed-����~�y�\�������]�v��E��s[Z�C� 5䣷!
	��cf��	�=����1�	��Cp
�~���ERLUj�A��U!�9<G8�܆Us̋P�c���^MܡD��j	@���#�n���0������AW&96����4'��=��g�Ty^8�N@Lb.�4��5Ԉl�\�"L��@�+��=�a��cB&���U����V��-x�̧��/}N?�8��,\�e{�E`ޭ]CQ���*��~�]����m/]��4K����W�2���MSPjEUUW�A�Ό��^�X.<D�J��0C[�-pA�7n�o]��?��W��W>�ex��������R�f����/�܅��UA}��{�󳿂��MOxJ��e�
�c�Kh<�,�e���i�h��c��Px�_q�L˞�{�#!��l޺�^� �wOz��7�~�@c^��g�K��p��/��d�ᆗ�{p��	���~�9n�ý�-8w���֛�`݅a������O��&xy�<��(�#t<�%59ġ'�'���@#q��v�K�[^Z6�������{�����+߆k��~���˿�,w����۷>�W�{�j#�]�1����s�='��l��ks�ݼ��}^���pgwZ�.8Ē�뎒$:NI~�Lo���Ŀg��T��+<���>_>��'�Ga�oΕ�U�B
�N-é�<1�����!Ĳ�ҍƿǳ�Z4�4.��>�	J�ܾ7�`1jq�b �(]�o ��Fn�'ݒ:�垝A{V������I��~ά����f�����⧇_U(%2΅4x���^g��Ȟ���)����@��ynL��S�aX��/^~�Rr������oXt�H�{���L�)6WUS�AJ��!\�[/��k�1����.��������(]1P �D�d�C�K�����T��l^���Y�s��2����8��.;�͛��k�)d��"Ԫ110D� t�
�w��?���2ln���O�]i1���M=Q�	9R�U٦�-����&(i�bSh]��T8#��!����w� ��߷������'̾�i����f�`�`�h�y�o�/~�]�Vv=��]�]��cZQu�; �
'68�[�!���J�m*�T�����f�"��M/�9oC�0T�3�7����r�b6�qzu�1��1�m��������b�ݠ�UU�tCÈ
�EF��U��L|�� �
 �����
e���z��K;�����.�-��妰�q��?+����#�b?�&_�N)�����*/Lt����OvX���Z��-r�ּ ��5(�\<�L�od�$����.զ[�5Ӂ�n^<�4h�@Q����A�:dk����񴖠�"�(@�DI�u���Lե|��X��w.����窓�p{�ň��~!��Z�K��O.��7�}	N��t���'�K&�2դ�;�}�k`�,y��c�{�ȫo�͹~�(�`��+�*�(��E���@�T�W�PTڃ}=��}��H8X05�>훸�Q��������{_'oWad�0)~�Yq6�KSJ�*/��L%E�*p����X�*��Sa�+�b�d���5��T�Up1li�9�̶�	5G�&,"�"\hw�� �� m蔢�TƆ�ѣ,�g&�DTHTD�J�_Z��b%zڱ
*�?�Ѽ`1��"!@�>R�4�:��8:֠����đ(���bw���@r�D��G0�Ɍ�X۷(U�${������ͱ&Zk��@�r2
���LKV0�X4�\:g5���ʟ6�d�a��)FqDтb�5]KN�m�Zv֯�=�Lesf��a�B��n_����y�F��Xm�:Q�=�Gr�8�=SY�0��u���׬{��s�=�W��lk�=J�f3g���i�����ܛs�I{Q��J��q?�I8iݏ���,ŕ�/�5e���	9g�s�5��x�x��c�h{��	�k��G�L\d� L���p�����KоX�ݫ税��q�%��MC�m%:B+Ǌ�+4p �����:%�M�	�����CjXJ��D�������x� �@(�yG+�tn֒�Y���ID�G���F^}k$L*ǃ��>�� �tSJ��`׃���l�%�at����%)���H[.�N#�*	���f5�4�'W�=��`f%��t^��)��M�M�(�i`]ӡS�A\ْF�Έi%,b�5
�Y1^2��275�Ez�5*g��"Y���D�8$��R�J�.�͸G]�9�\��V�<��1�A���y0�v�e'����YaM.�+D7<����(W���["7�Z1��3j��R�9������AO>��S�Oª�����A�v���k��ϏJ�Ț- �Ҋ��hw>w�1����U$����j�p /q�E!]?�O����?	��w�e�	��y�g���;��� ^<r� �~z�]�ă�{KV��c͆{�
q��N�ʒT�Rt�Q��N�Y���U� ��*fU��� �g��}L��#[s��С�&�U�x��+F:����F��"(h�Ǹp�U���?W�z��K������g��Q�p��!{`�N��@�~�U��&�0�����+-|)dr洜�@��$,"�;�
�,��A�Ҷ�4{��q�3U�K��,�^IZ7Ľ�8h����V�c��̢��3F��*�^�>�D�J��� X�A{���J�1����m�Ugy/P�����@s����J94�t�$JЎ���!])Lw
h�&"�������x��*��CEf�C�\������0�-��<���u�`�;p
.n߆;f'�bQ�kz�����~>���N<�18�;K�7��M�xh� �5�d����t`i�j�/�'�<�w�®��s�P�Q͢�(gb$êm B�7���O&n�UP�=Ci����
=�8����7եg��C]9%��<(}"A ����f�[�\��H��PN�7�a�%�j�;9EB@����X*����H���:)����Y5�@�t�++�@�s����U�����F�kޱ��z(�TZ�"	Q��	f��n��q���:��$]������UEB��B�U��hchu�-�&L˾	`�_:�I�Pe]�[5���u�U�P��⬈���yT�]K^S\� c�x��4ٶ��%S�H� J�	4lg�K��7'(�+<a��i�~�ǽ$���nn�
"�GD���`��墝(~�P��Sq:���1��t� �@����CI�w�/�=�8�	�O���(F�1�>����DzA�
��F��C�+������Cn8�7�PN@�օ8W�(d3��1~V�MT�ssC*Z��A��|���(Y��Z��J/@Tں�g���J�B�����py�Q
$���� �B "���D��rY��i��_D�d<�q�A8ҧ
������Wb��I���Y�* �'*�qb��pvzp���LV�$�L+�V����BpPh�H����-���� ��A�B.�'��AH"�F/�	������$tx��4����eӾ�U|1�[i߰���g�5����iѺ�>�X�&�~�Hy�l��v)	�0K��ˌiݴt�'���:x�m�Ո/������j��ce-kaq6�Ǻk`F�#�Ţ03�<$�`�WD��
x��q8E��[$��Z���/�f�(�Q�Y��=�C��M�壢x��^�B�$����r�x�CL�]u��L�K�s��9����+|�֐�C(�Ȉ�S�K۴I��C����ϸ�!mL&5;�Ap�!�m�h��S�������:�T�T)'�H�)�"���%rn��7%�W��`1��!��$��xU킉"�ȅ��R�|��S�Ә]5�5$ve��l3����#2j���O�k���M���ԋaf���Dd��m�d!��|Z���Qˀ�ԯd��(I�tl�`�f�H�z	��S�k�\T���E��9vVIJ�$�`Y!��-.�ATt�N	�E�0�M���2���J��@Qe��-��9�ōP�a'0���6y�?p��6�B�\�gU��׽�%��H��^b�D��W�{�O� ���b��	�A�f�#T�5���nN�a���dF	nl}r�BU	V�tcۤN"9 ���sO+0��$� �n������ݔ!(�	?u3��pu����Ad�,�P����*uɶNU!P�@�wڎ	��B���Q�T��l���5�BU��&�*i�s&Zp m�>3a�0Aq�+6ِ[p | ����]P�
����Kn��;����^�Ui"qVS��0�o:�3���m���+T��J8�K� �����C�n�8JuL���H�N��Yy��8
Wd�3� �--��!!G�'� $(ȊC7+H͚.�,��W0���ь�)�H/ې�pY	�,VD��@ZLoF,���0�:0���$��7Nؑ�C���C)|�0L� (��l��ť��;���V� ��"��J$� 0���^�ҭN&�Mt�L!H���'R4�$LF'oR6�siay]���e(}+;�����!���6�9PUL��6����V_A��3N��M���0�>�`�dN�y��u�$�?n.gr�:����P�ǸtۈpVEo�Q�b�S
1w��le\ ��X��(��*��\?sq=x����M�p�֔J��T��9P���o$N,Z({��rO���bL�q�M���TgJ�Kz�s��*�	aşV!�Wrx��@T������(�yfԼ��lD���ڶ\pj�'�K�k���4�>;��_�ҙ3�$L �;Z����A�BdmR�Ō�"��.4�F$�c�re2��#��;p��X���'�cR�ڎMI�EI�8� rO�I�YJ%e��T-�Ń�/�4H��L&�Ĵ�:.�"^�'҅~̚ ���ʍ��� �E�]���B���?��焨[&bFD��ݹHD������\�ΘUmv&����fPV�Щ�[�e�?�F�؈���w����grl���z�D �����)�N�Km.tT���l~�Z�0�h�Lܱ��� ����ҭ�].�$k�Ղ "�)q�u������{:O<��7�����4nR�J� ���������"X(��o�:1IJ������A�;�ԅ��Tc�o�-�*)k������z�d&h�����X2N��W&h�&�D�Nɘܸw"�a�q����jy�m���������ژ��,�����.tW{\i�`�QAf$�	��`9i2�R#ZpQ�mؚ���ުBk:e�R��j��̎�LȞ(�d�Z[^C�r{�ih�d�����_��<�P?�6c7K�����?�"��m����z��UH���o*�p�a%�B�k&Y���K+>�5�U9��#if�d6I: PS=/�*0IF�~j�)���}����o-�.����A� �L�~Fp��qO$��:p끬�Gm���Na��䞤�\&8�N���g�Z�Zw�@�Z�sS��o��2*�;�Sq�a3��*֏6\�i�]ۂ�v��&���jva�cI�zp}������F���0B��"����@*�9$��-YqN:�aY�*��#�վ�j��q։C��;nȈ%( �L7^aCa�8�
7g(L��_�mJ��X6�r��و�O�XP���c���&Ң�7��-��C
T*���ƥD��������.&W���xn
�����N	�����G���p�~䜷��J�8�/f3!�f�P5�������i�A�7����o��1�K�WRR�%b��'<��e5��+c�X��s�#���.Z�2c)��Yz��O�	�:�sLGPbY�%I]�a�<`�=�"�ٌ$X
��0�s4gʂ
�n�r�al�OBl\��	2� ����Rd���d��8Im#���w ��䟋���3���f�: Q�*�KO�����Z��|dC>WQ�S)���rPMQH<&��on.�a�|�y�L6~(*����h:髕��v��)z.��f��\d
1�q��BA���Y�2��DBL��ȸ�J_�&��=��~��征��h8�V����t�`�n&{p�X�x3pX#i�:.q�QU׊�/#;dB�R��H	�G�b���hc�&�֢fc�ww��L�0�v���$XlU���j�rQ�M��)H�-\�Bǋv��W=����E�\�o�$/�@@����a����.�/*,�?���c��#;,3	���"�X�4�;,�5Q-R��r"��, ��Ñ^���sBSۼ'z�H;�F��'�7m�"Q��3����6��6�@.�9�j�J��̚�UU���g�U��׭?�i���%��K/��4���(���<)�3@�)9�[��`�eB�lb�*�CC����;%L6���p�D+���4j�D���Х��:�?�O��E�f)���a�mR�s��)͸�0�Z:gaڍ|ϱtX	�4��R3�,�RfTie�Ma�M)��$���}�WM���(nla*����ҍ�ڄfU��������<�vn�~BO"�?�
��x��l@A4�2lX���Md �D�FH���s�����Q�	271t�C���fn����K���.��(��M~���ߑy�%Y���$YiG��Ԯ���?2����6j�z~��v�����Bk`�i��AͨQN`C�3��n5
\��aL@܆N��ʟw��CW��"&!m���$-���i�&K"3�n=�X�~�O�8f�G>C�X��GØ(����%�hg]�Y���R1YT���=�Ma�pm�l²�@�mC����
���c��$� J�=م�M*#���!*ӌp<����/��ß�#�T�j.e���H���pbe	~y�u�uZ0�������^���h���"���d�5<�	i5Otc�C.R<<�|ue��~�6���ε\2����sX�x��"}�~]mb@��
���4U�{��}9q�]6?��S ��D������I_��Q�Ld��KU�R��j$5�=55�o���4]��i:Z�Y)����b�DV~����h%�|�3q.�v�><,�0Xppg�ۓ!.�tb�~RW}��kL��5��߄��:�@��e`�XZ(`\:�5��d��j
����=�AZ)C��a�RF�D�	ܻ����M�t�L�3H\�nl��s���;%�2����m ���ov̵2SD�N��s��4E#��vHd{��{�Yڐ��fb���fOeJ�\j��%҇�j�F�7�y|�.�~�a���r��=�'���q�D�g�FP���O<*�ԅ�t.�	)Ι���ōaB�i�3��E�4��f��K�Ĕ���6h���M����� ^�r�>g�U��\��H�(���l���ī�pes޹v��YE�'t;��1����}�{����BU%�$:��n������I�* A\b��
�5p�5��]��O���GP��"IRj�#2Hv�(FE�-8�,z�I����A�M���)N������P"�Y��v����~YE�;������/�f˷�o�$���@Ą	��*y�g�0=�����]l;2�*�>ZVUi�U8�WE�&��˹�B��!7�s�[�Dec,(�����g�8¼u��K���];wZR:��@��D, 5=���e����f�5��Hz�˾�W�4�`Z"�W{$C
2<�*�.�y��*��B�zG�*����T$U#X *��p,���7^�^�o/]�1F�mX�/�D�*�b�ՂE�AT^�����3n�&���K�����ѓ0��g�2�r�2˃�>D��JoH����O��s�- E�oFp~�\o��Lk%�)8�p\I�ہ�&?�m�������OAkba����4\�t�G ��(vD��Fp���~�Y����밋��$1�Z�e����$rn�p�ro�l�]9%č߃@+(��
!*šV[�6 �*f�$w���F\W�3����׉���ܽ'3��7]r�#��f�i� �Xc��Qs��}�\J�i� ��*x�"��si)����w'L�_�����~7��$��U�ĥ]Ԥ����4�=Pא��	fbJY����Ϭ������\J$��:~�j�QM�TF���R����57_��H�4�|׊�qR�+��Gp7��nʥ}�m۞0X�c��`���R�	�:P�uX��� �<���R4���!��۰�i��]�kU�������2�M	�n��˾��n݀�C�C{�K��!B��M�t� �V�{g����[p�3��+�B��)�EAT��S�M�`#�2������4�Lm�MoDb�{�6όe	�Q0��	MQ���d�a����R`뽈�~��A�����0��X"�I잀��'U?�U�W�[-z�;����g��1 �$u؇�W3����~p���^M��9j�1d�I�	Mƹ�(��(
��h��~������˲��Qi��^���¥�6_%������Ð"��x��f;]��omހ���aqm��d���#M6,Ef'j��qM?bF���c�va`gpn�&\m�d�]Ո�uyVi̢�*D�wp{�o� �{=x®����"�jP"�R�~W}hhƻ;p��(V�? ?<���T0򜡃�ex�_B� 9¸�&n�8g)w�L�fv�D�QT*2��+��L��rU=e�Bb-�a��Dns�ė�mi;���x��$�r�!�O��� (%a0`kj�k8�Mܧ�O��ɦ�R Q0V�!�a���ΈWf�_����R�ƞ�5.'({x�����O��f���q�ET��@�����Rgl���2��	&��SKWࢴ������6E��i�uB���%Cc�Ph��N�0��r�K��Fp��U8�^��n���Y�������w��x�Iާ���'
�z����|;-,"ZR����R��`�8��ș1��wlÎ���au���>�q�m��ez�~�N]%�ߪ&p	��Owp��i�:G�OϿ�Z�V�xm7�TRYq�{1j��7+óCLT�L�:'Jr0���a�±N�7uX���D(4��)����J��3F�A}
�MfLbǬ2i=��G ~\��hk-��;������!���f�λ2`�J�}Bŗ�Es�(�I��"xٔ��o�t�3�	��s�P���R
s��k`����AiJ	�}N����\3�߰X?�����c�q�0=i_�-[�l@M*��3�XۛM��)qS~�D`�?�Y�/$�
�FC"|}ߙ۞������Fu�O>G�WZ�.A�rx"g����"�+����#���p��	� ��ރ�]������i��y;�.`�:������O�/��z�2,����o�ѱ`��=U����߹�����)��뭬Ru���!�b��5L=w�q�#���e�&)�9�u��01'4��!h���LL���ҋ�D}�d�Tmd�8�[ik���+n�Fy@�U%ܴ�����lHt�U��'����G��g³� a�2δ�F�n �q>�դw��;�0���v!˿��}�;����U�Ev�a�q�~��^�������8��^�k�F#*�>�����0_��"�&�=�Ɛ�k�W#���!��A|G�E�F��,s���N�7��>OeϿz�q8�r�j�9,��Wf;	�Ʒ��ހ��-8?X�m\�Knv-���̻1tR������x.��3ۆ��>������-��ɧa:����X�[��&�j������f��s�W��Wv6��ހ�޹��-�x5���Q�;�AY��O��_
�K	^O��[(���6�db ����Q��F��j���ĥT��{ZQ��f���PY8�Y�R�D�pB�]�(���K����y�V%���u��ɉy$ ������&��6�*2�(��d��gD^�;��z����TI�2�ZB?��XWӳ~=�H�Z���9F���M��'�M�c�S�B�@�tJd��ØR���ӭ�'�5L��X�ʵ3-:�������?����߁�O?�U�a�Ӄ�V�`\ST��1R�+�T�8XO���!�/���t~p�"\�6`���1�dh��&���z��fI�.U��BаB���n��r�=���g�ع��@\��6u�U�)W�
%A	޿�^����>v^�v�{���_�I��p�R�SX��жblm���bC4��ڒ\��$-��@$㦑��ˎJl��y%R�rs�����-Hfv�o�h�v�T*I���5���y���D|(�f"P�U��BĚs������)\�x��g:?��)n� ���%��&���i�{\�Ed��/&Tf��J�^�a����F͂�=�p�*���,ٳ.&�D5T �;m}�J)ƨ�0/-+�d�iN��*(m^��Fv�;�I{�i��~��h���w����&|��x��iX.�pl��.-�����(P�����8WhG�,fs�V�=��p�ع��� n�>�(����L<qmAo��U�$�빕����8lG��;sXBcc胝ͨ�ְh�]3�w�n�g���z��0��n�u{~�8֔Ru�"omo���ܾ~���S'�����\��ߺ <W�]�ЛM��7QU�:C���P�ɒ����*岚
+[��	n"�j��F��:��LB�eʈ����R� �]��Y��:������kL�!@Z����$��F��p
Lxz��x�!�OFǝī&������c"�KI��Ɉ�W��� ґPi�:U�mY%�:㉓kC%�BN!�sc��KI��O'җ�}
��!�U:��w�N�K��z���H�朙5�ݪ���Co׸cA݋���_��祐j�hg�?E�H��*����d >����*[�M
kс)ZYC�sH}��ό�����P�P�􄐥�
v�	L;]x�.޻��^�'z���cg����#lXͨ@j+�������k�3�#	p<�w�߂�o��b�����'\�����4�21�����{c8�#`����NYuT��o7�G�ކ�^��ťP����;��y�21�~�Tu`:�6�4���K1�+���S���;����pi���.�h8�\��{"kK*��@5|0��� QG+Hk���L�(��4$��%����ya�e%��&MWt&撧N����c_�mm��	�S�.���N���H�*�����H$3�:�xܡF(�1IK�f�Q���VQR���Q�5B�:�b2I��� =�1F�`#K�F��>aaꈰGϜ		۵�d�,L2�=�{�.�߇�c\]�D�����Wo"/���*�q�ψ�9c��]a�/�Eayn��`aP:O։8#���^[�L0���v��sa�Ȧ��K���=X$82Ԫ���~��v��S](�0L�A��g�+�.��준��$&�!��:m��n�{�'c��i�UD��D{�)�l���x��[T�1�:	 (�"���/·n��m| &Z����܀��t˄a�_0��z�'���g���A
�2nf���"�#j���U���l�؂�� �;p�W���l�&�~�G�|ά��yE%��Ș�l�ܳ@�2Xw��*��j8\(�ѭs��ą�g|�K���ud��TT��釠i�d�@I�R�9J���۬B6T�7\����fu[3�[IgrK�z���[m"rF�-�E�.v)C���*Պ�mxn ( ZEr��2y�2SgHq��ES���,c�@U�zd�qGD1[��d:S	k�k;���6�*u~�8f����9;p��*!���R�9���� ]\��}���䂮�+���F<��T���sQ79X!�D����~X���Y��g��L�==�h;#�-P�_���5��\ނ&�x���za���5cOS����j��A ]@)_��M�^\~���%F���� ��<���_��`w<%����U��t	�j#O��gw���یH���aq�K�X(8��[-x�����6��?ܩ����s�g-? 3��z��
��(E���.�%�.�^���_aByn�P���q\E��H�����Ô�m�"QE)�J�*�Q�K��K%.�.���4"�N�
A���~�D�Q{�|�y�߁���$s��3�(\��Hm��A�=uI��{�a�>+�̩���D�M$�%f�%��g�C6l�����LUi��c�ci2�2 a�ɾ����iV���v,^��Y;e��cm)sL�L�NjΪ}�D����J�g�6K��М��O���)f����Z߳�m�!ג+�K��5�[;�0��m��(K�5%W��9�5�#��ݝ�8��=b�2m����l���V�OK��g�ܔ�ia�d-���?��)�X���_    IEND�B`�PK
     �9s[�īd}d  }d  /   images/ef87c5cc-d843-475d-a868-97060fb00c54.png�PNG

   IHDR   d   l   ��9   gAMA  ���a   	pHYs  %  %IR$�  dIDATx����%Wu&�U��:��yr��h4��Q�H� ��MX������:/����5,�`�0 #PD('4�䜻��sN/Ǫ�wέz����mu�������|'�[A�|a(=��S�җ��o|��于��{���|-`ِk���>g�����%\ؖ����׼���hU�t���z�,���N���_����.�1_�ի�K�4q�5}��|ǥ,��K���+��K�Z� :�M(��~�	�~y�,�԰].1��l��� �2�be�� Gdq��Jyo��W��V�7����c�"����8�ek`&���t8�
?��4�_�u��2��o��l���-�meq�z���cp���㸪lz-�w_mD�lۓ�Q�%���x°��6�0�{�XA�E0�r$�I��!~q	�|�ﹲu��f����1��ʥ�""�	��FP��:y�yXn��{�y8�2��c�1��:Nut*���������b{��/��%�[�"�C`Fê��8�,�/
�}f����-������^o����c��a�hY�h��uu�rъ��G U��QQ%*(%�k�b��p��T����R��A]XG5:	!i��p+�%�9qù$��s��E�f�%~�\Qs+��,_a�Y�Bm�U�D+ep��B���iU*%����:��!�7g�bH&���+K%Bӿ��ʸm�X��F3oa*����ܿ��Q�ϙk�U������.��^O,* 3�=�I����@uR!�2�j�Gm8�Mu]��Хc�ϥp<;���:��"�]�jr�fuEb>�r/�n݈D��rI
��� �3t+iQ�f�D!i-v�he��7�pd�Fc,����nE�k)sYo@2��l!����K�i�V�VC��r��J�(��VW���x#���it�&�`fK��%%B1}m����Q��4�"0'+�p#	�.L�кm��'Q���\�Wem}'F&Q(e����r��*��Fk(�L��l1�������ι�J���Vl����l��;6"����V'���o�pi�cq�%���s��h�����`G�VQ[�jb���6���-��]$.R��x��TrQ�>�;x���B�K!s��[w} k(���Kعv�?~ _z�[��s!�ꃟ��|
��i�.���k���9�����_F4ڀ��A\��J�������~�@�F���s絸o�=��w
:z�1����;ʶ(E=���G>���.
b�����-N-��P�a������i̦p͆����>��.��?LW�{��P-N���[v���G���g���o��k�_�|7�6��r��c�Cu�����b�2H��1�7��xw�N��B�f9c���v�n������,5��:j)%Z�j�`p@�©b�S�{W�P��~�	�!��bh�v׆�]B��ʊ/�nj�5�wcra+:W��C�i��|���[H�֠��a:���V:� *Ŋ���hB�m]ؚˣ���r6�	MZ�X�K��W�ܠ��Ќ�VS��:�X~�um$;A��W���l�-u	l�݊�D6v�������.�G-�WW]��00������ih�Gڷ�N�Q �q�Zb	��&�x^滼�v(�͉N��Z0�P#rԯ8:AuȮ�a��Xdq��xm��%|�ej��bpnۺ6�~F�NH���/?�1tpv {)�K3��q!��ҏ^}�t#�1l�^���IWh�2�������N��ê������	\/�Rx������b����T�r	��B�{�'��ŎU[037�0'W(��9xz��^����믢�Ω�/sqVRYv��[���'��[��Ѓ�������D���/
�>ZCm���=GHg�8�ڜ�R�u���R�U�ǿ��
6�^��vߍDMb55�Ɠ?�����PZ-i����ԝW����|��2=��E�C����PK+��k�?���8<|�N�Xaws;~��O�w��А��G�Ɠ'_#L�	F,�y���������(����T��e��ص�
l�m=�Z��8���}'^;G���sn[V��-�o�:���g~��ϝ �0��L���ť�q~Aqn��q���/����W2��\!M��d�#�,��J���P�Q���MBPQ�C3-b��/=��B���O���cx���	���|��'��]ă�yS��'̵\#�o>�#�R9|������8�w\!�����}�O�&�-����=�׎!$��B�Hj
���;��$v_u�<�sL'�)��"���z����;?�U��?;����H���8��������\:�KS���D�s��:���EѹF�r3�aX�8.R��5�[ą�$V�w��Ũ�_���>L,N���T�'h�"o�ؖq��w,�˝�8}K�J��S�}���O K󟝝E��+��I���F��{?F����7_�tjVWWԗ���m��W��1d�yL�̢��F�!�(q1w�݊���A}þ��x�2�8d�=������ݛ�������M�KH��+������T�L
Q�ë�*�kۻ���}T���G��P*\';��p6���ø����KY�&��1�����1i�����7�#у��V��a����C�����q���d2Jy�ʢ���~ܣ��Zl�p��=#*\vο���oQ�~B�(�v����ߢ\�D�'��Q e�ܲ	/�{���ba�Sc�Γ?F�k�~P���E^��=��;%sF9࠳�U�"���r���ã�x�k�Ggk��D� a�&T��g�`xr��OdnAY��It�6^>�6�P@�aC=�2K8[�bad�k#��޲ʐ%�j�F�f����Q䜤�!dO��2y��d�V�4�:�>��6ln��@Of��f�:�/���c�����
�XQm�.~$ส�?���m����B	K�{y݇�����W<�V�|�
"�q(�'�|��I?���o���YeT>a��D�?�G�!�hD���Xhc$����'�c[�jܴ�&B�?a��)R����^������8�x�u�pa�j����IMc����".O\�o��c��7��P�?�'���tn�lm3��G B�#��)��Ȉ��V]��P��Pr�gώ��s�~DEa��w2�u6�'�+�c��7'�q]�&�LtQ[r�?3���qL�O JS,-$�ʆ]�F���Y�q�����[O�+���"|�n���?�w�t�vu�"ٌhx���E����.�fV�v�];�`�o�p`�=�-�
ܵ�f�}�(�}�mH�7cln�V|.�x�T�1Z��k6bC�Z|�w���/��s�A.�]��+��s5޽���6\�k/^:q���<撋��9<p�=���{���+�y�u蛘����j��}�Gc�6����᷿�x~��C���"��Q��9�����N�3-Ж�����O![Z@�-i�A㐒h�8�<�Rs�,}D?��c�$�+U
�
y���`ɭ�KDӄ��,��N�.ѺS6���;�6���o�L?5�~���W}��s�#l���U�('5??��7�́#d%!���܇������8.�C�����f~y�;8�<c�F<���8s�$�)�P��̠)р����H4�^����ʄȊSB%L+N%1<5����_P��46̹($(2�$�±L�?~�g��¬r@aա/���.cbv
����$;�"s�s}B��D����$�$/%�Y2����.(�` ͸jQ6(	01�'X*z�P]������]���5FĚu<_"oK���9�`�O����q�^8�NU�����C������_xg��0J$4](�\�k�<��C8}i��. �O#,J��0=p�/a2��^;SȢ>'T���gF���_�"k�157�E2���a.��Nl̗2��G�['�`Mw/�i���ӄC�7�2Oa|�'c`bS�)��&:X�Q��A�a��"��j�4@;Ȋ#
��^�Ҁ��,犔����&]����?�������]?�NGZ���S�L�V���	/�n�ƪ*��5xxq�|�G�e�K�J�^9}g��+f)� !b!��Dd�P��]��J�E��PH#}IT���gi	_}�����[��������g�zɔ�'X�QAu�2uy��^|B����~&�1*96I��w氦�%�n�O/!D�P�v��%Z�M!��|J�?�%Fd��ۂZ�VFq���z���d�d��J���z���i�՚u5�|_`~^����1X�G#c�����9&Y�p(l��Z�2,L��
9i�8i��y�<a̯�~ ,0`j��ҹs�onbL��˘!LDȈDXǰ� 4ƿE�!U�n[����hE%�ɎM���M����,�z��|
qKր1���������3J95M#�& �!*�:���z�\�$����nhۀ��� ��!S)��.��043L��P+���eDmǨ�f����^w]+IW�N����UOS'Fg&��y�Р�1���g����~���ш.X6��t���dO;�|
��F�� c^�p)�E,Vm�Մy�L�x| -�4�z�'-L^^�k�D�l����T��@f�Hbsj%B�+DE�D�h	$����ep4��R��y���Mp�Edf��\\���φ�5����O�����CQ[�G���B�O��AEuZD�a��~��G��wo��5-X߻o�:�W��=��{�6�iܴ�F��?�ޗy�k��|
}#cxr�S��3h���ן��>~md/r�o=��fG��4�u௿�E�$bh�5j�0�Z�%
9��JPX6:�@��F%3���m�� !�v�NN�-^�I�!��tp��<�kj01��	���\�����0??�ɉ��JY,�ƶM����З�'�>æ2I�ۼn�[p��%�F	3�3J�Mմ���l�x5F��0<4D�/ҺJ�󾥤B���,�rY_(��ˀ;R=�
�N�Jr�_��a���֍��5�Z\�t�7nC<Z�֦f�
���[��\j���Ok.f��M��-��O����[�}�������B����Ϙ����ks4�=k������ts��c���SL降�6N2�	aaa�v?>��UJȭ��]+V�{�Z�ajag3}(4Q
$ x�����kv�C'�܋o�H�hl$��"����w�V�����o1>>^-��Muq|��۰f���/}�(�u��RR�U�������GN����&����g12'+U�*�v���"�]G�E�ly����nR��һ���`���� ���7[�։��^���&�
��ZZA9����RfIeJ%R˳������'98��q򮦗���\�]�v#��cnn�B܋�Wr�pr���JR���8��GUYZ��d$�N	y�H������c'��tS���&�/+�9d�2�<�3��q����s8���_����ɳS�>K�}��[C�����ɹ~�3i��Q%~�.���IZ�C?�T��=#�(m��)�b�Mh���I���]���L�����j���J-O=�{��F�`?:���j����q2�ؽ�
DBQ\"�Ţ8z����t�D��"Q���6l߸�|<G� ���6K�V�
mSR!��.tut���	ZP��Y;��5~~�۹
]=��kq�lV�����vጦf��ظi;��8���21<@�*S�T��R��^HcdtF����c<#N]�l>��s����l�>"*) ϱ755i~-J�29������E;�9?;���V��/ �Єd���c�$A��okoC��x%bɝI0��^�#G^�
��3�����61\0�}����� :[�a���������'��:���M�z�o�׮C'������ï�7ܻ�f$�t����]������ܔPp��!\}�6��Goݯ��D�z������I�POGǁSG� k!���[/���;��Тb��sx{�!�O=v��{�9�x��8t�.����:�h��ID�#��F��zGg'Ӌʖ��.�43��<]�V����I�?"B�{��o��΅�S�j��X���[�<Z��M�,+��g~](���i��\�e�!~�0W�u���76k5,Ɓ?���r�\�b�����o���[�a�&H��]WߊG~�(�f'q��9�w�=�1��x�_w#N���ű!����Zj]��N�@c]Go�JH܈:����F�P���G��@�����vvoR�|��a6����.�j�����i�7��c��D[C+lYe�R����3�ӚKJ�S�ℎ)��I2 �4Wr�.Ʃ\(K�G4=*���>*���$�q��j�N�.0�>5�.����vӴ�,tLK����&hi�д��;�Ğ];��"�U&߽c��_�2����ş��r���2!/�A�[����?���*�޹S�'@���?\�0����ѱ��s����V޻d��t��У��B�{$�&�l��T�`��-��fI���"��9���s8x� �5bR�V��W]�k���t�8jdQt%ZM��]�w� N��_WW�0	E��	Ӓ� ?��_}C=j�1�t��7$(쒩��ԇ\-�ڵb�^���z$�g�����ç��'�,�H2����Z[˝����m��8@����_!�����ܠ���^]�/��a�E��ױ(�+�6�<�ɮ����S2Eq�����XZt�l��% �RR��j<���Y%�U�  C677�Wm��+�����k�+��c�H�$�*��\�[Q;a:�R�tD�w��S��7�X*R
����܏157nzE���1�$�z��zR�%���-��w��8q�$�صM�?�����}G��-ZR��m��&lM�����/x<D�]C�"��D	�с��*�	+���p}��LJ���B��������y~O�V�Ԇ,�d���T&=��W˗ɉP��>C�����6����՘D�[�v"z�j#��w���3��(�]m�x�s�pg�r�4�;� iu����Y�0���x����wǤ��"b4�cH����5��r;.�E�
d�ͽ��{?����Ǹx�⅐��O��4����CMlm�����e�Q�����R�8f2��R��$0.b�|��|)�-j��y鶘x2mY,X���2��U?Ro��I�M�%�\���=)P�-��⋅��I$./��T�Z5p�B��%G&�Mʻ>K��jUY�4a�2�t�Z �k��{\jK8F��d��or�=�l0U����9<��v�rx�d�LR8ID���O=�4����J&R����B�,b_BQF��	R�N^o�xǗ�	B4�5�k*����UW�¤�j-bo6��$F$)��D�P �qLPa���d`��Y�+�-���i� ���$/�;�b�6�宔	�b$Ky�P��Ö�Ŋ��5��Y�dm)��c��@��Ԕ�	G��M^��n��*�PL��E�� !������9���1:9������h'��w>�o>���N�8M�`a톕�:�f�N町�����,�V���nI"�AT������p���� ��مy�뷮�"�cȁF"1�$��*eL;*IE-W���)*NT�)���Q%%^<d����*TTR�1:�K�R��(�m*�Ƶ�Q��M�m��3g/�,���$Wt��6J��dQWA����q�0�J������	�lV��M-�8ra@�A-�Y�Zס\�y3]�'��	^0�p�]��c,T���(�$�a:?
`Ug7�f:�S�H��.�����K/R�j���-����05=�}�Z�H��&�PR�(#ː���S�c\@+�5�1Ei�d/A}���,��3��4%�181���ndK�������vwtv`th@3���gg�(�N@}VgK&'�11��%�	.ǟɉ�ʨ#fx���I���b�*�H2ֈ���;��#"�m�kPb0�\@F�%W�~ㄧE*��U�z��i���d��ѐ�BE���/T�,c���y�v~�L��LE_D;)�8IF��p��PP��_Fz�`�[����;Ǡ'��h@�A:[ę3}X��S���1��AHw ���U�q�q�\*��Z�#���HW�P��y�K��!�^��{�0�\�3��{o݋{�w���/���˷��E)��}�^4���D햺ȳO���^~����{n܉�?�	%j��ˁCG��S�jzgu[���""��o����=��7�`���=�6A��(���y�e>uZ��[�ۃw�t�Rc�k�p�~���j1�{�����bu��)E�R��?x�A�"i��Nl�r�+����ỏ<����8:�`�����R.�$��3��Z��ճZ�LLN�\J���$�ΨPu�i~.��\Z}�����qcg{�883T��|���AK�i
e6���|E�m9�D����*t�X����I���.�)��s�h��J�N&�x��OhAM�ɕ[6��;oӔG"��eG1<<�M�!jo	��ﻃ~'F%���^ƿ��i�'<�p�u�y��(��I,����9�U=����S�������O=O��Dᷡ.�����&��jGG���>��Q��qܰ�]�y��\�0ЬVÅ8m�8պ�Z���X�`�݈��^@�NN^�y��)�E5���MYL�I��\!�ճfb�z�]t֗02_�\�����ze룵ZȒtICs3�G\��19��L��z�ԺYj^3!e|r������Z��<Q}}�h�|�l�55�kVb���D� 	�6�MA:�Ī�Qaf1���&*g#-d.S¹�}j!�aF��XR�P��Fb3G!��F"y�D��>I^(�q�2��	�JK�221Kf	�d��F�	bx������`9��E��2�q<u�uT�p��@)��S���]W��W_F�6��h̝�,	8�U��yDB�fS��ܵ:��%U�M�1����E���%t��E��Ke3Q.�������� �z�W���?��+ʀd�Ī�e(�-�r��ţ�?�'�}A�M{�9�\��6
[gxt���_� �����,S���9j2\��c�>Fڌl*ڏ�}	Ͽq�K���*L}}��|.�?��Re��&��5T�X�P��~�!��:��tzW]�	C$�(?�{7~�N�@�����~�0S��^L�j�׎���9޶������LY,��pCg �tU6��k�
SS��"(c�_��ij��V)�<�8Ny�ˣՔ�T&ˮ�,��l/����V����DK����l��O�lSK&�j�!��J�ۦfb�<aȱ��с��B�FI���d�%.�S�����2���Br1?���M�������4k�"�N����:X�u�GY�P�h�D�5�E�1���fLg����Y!��ٙYL��1�f�V�TNZ|&�F�4݈%Jdm�#\�-L��@?#Q�]$=&�K��t�E4���I�ߣ��\0��-��@\���M}����.}�&!���E�Ԇn�'i(�$5�~b?Q(_p�5��Z��;�ྣ��>e;���S�R�f��~����ZQk�K{%����KN�Ń��UB1	FmZ��_>���!���KV`q�>�+�?z�9I[��7_e�S�6�Ò�
:����,Q�4,)X��!�2��G���(P�r%Uk-�K�S�i��i���@���f�j^w=��7y�
���^V�2m�~����z����ʋ��ZZ��Tk�:#��(��P����R쒂Tw���Qk�WKw�M�~��5�R�S�.�7��K�hY��i�n��[��=��W��������cۦ�u�U�?}}�#�,���n��Ԃ��M�׊����%A��FM_������]1�
~�S��6�f@&y0���]j�����vj�������
�5�غ��5����S�۫䯺e�e$n,D7�Z�����j,E�U��dVUsͥ�e�x�uyW�m2��l��О;p}��>�e|p��x,�".����2(b�157��ck]=�����F���!�+��{�,j6^���9��A�N3e���=u��R�p���DK:t���Im���_ܵ+��}��7)�D��޴t�{+���t�h�ZP�}1t��A�ÇP��tݢѰ:�p �~H��R�֊&�@z�²͙�x�Ԉ4F��T:�����[�/�(���X��f�A��n�v4�E�|���׿�9�u�%�p�� ��&�yd���l�<v�.��-ل�jYV&&�m��6;"���qѣ(�dJt�i�)~ϹZw.J�SE���HO[��!�p&���|K�B��]�5Y�P��My�Էs����#pea#wH��qE��јM�T�ZÎ
�@�����}�t�6#�EI��~Y��%Y)הk�R������˿���d�����
�U�r�0�8��m�莶bln��E~�G*�m����I���k(ЯH �O$υ�#��0�]Z��ZB�����4R(颥��y)X������Ӎ!l��S�/X���o���_�׵R'[�y-��Gj�&1�ir������˞46C�F�ȟ�S1cj]#�GMƖ���Lj�Iz�jk"j�E��c��)HXb3��?�C	�|T�k��F6�jK���{�͋���{����U�p��$�猳�BKU��ދ�G����I���rrP������&-0�2!�V�!,�H�i��&I$�����Qll~Z���̰�T�\f���T-�cZ�aK+���J�22��a_�sUW�Ŧ�������M���mr5�I��$��D�BJj�$���Pv�}�����������2.Ro}]�yN�I�U�OcŪv�����8��m�KG����
.Mk�^SG�AB��� ����L�kUMI��J��dI������| �:�dt�NEyY'����"a6�#0���e�2�TӪN������$��"It/��^�q�����y=� w�0�(���X�I�\hnK���:�,��� �*�֞T:g�e��$�)k�#ԇTax��W���:���t:v�~�-7�����@S��V���M!S�kKha��0>qA����%Q�ѳ�Qy���E��"�t�N�8�r!i�$ 1�*V$�n�@$�'j�Բ�-Uj�v`����u�P|x�R��*�m:;�$��\H���5�f��7��F�(���b����Y&h�<\YX����E��(9'ΣX� �,j]M��	�hU`�ey��r��B����f~��ͥ�������^³_����ػq)k#�S�� ��C��ؘЪX�p$���B��d�%�S]8ȉt�:�|�QzI���ϭS"D���
�Y�n�g��w�갫lŋ%�@L�w-�P*��5{�sU�<z+�@д�h�M(��"�����	iR��"y�E*��A��㫤"<�KsHC���2+v�+�K�w�@���D�'��Rk�}Y�r�^<��nP_�%tG���_��`Mw�NJr7^UZ����+�J�;Fj��+�,��"��D��-�/'E�dW���թ
\Np��-�4GH��r)��LS��i�Yta
�m��n����j<B`y8��E��TW|�d�i��$�֍<́��R�:�t>F�!U�D����h�X>^=ңdXVA��`����S�%|0�ޟB�B�����4��ʅ��j)�V�Y�3S���O��
W�W=5I=:=��#�,�9eL|��WK8�x�c�/#l9�0�����Z�;��X�G�uq�٬id��J� �Ai���r4 ��G*��N;"Pk�/���9^���Ig��ԹI�ʳJ�����>���D׋�5RU�|���`T�]r�B{sٜ�>7o6#Q ��R������59& ��=���ʥ5�N��`�����ڶ��#9(���z�P"�'�j}1��%Q���HSf�RR[��I_�@��l��c��/�Y���1�@o�K���Ҝ`�	1M���Rт�����ӜsS'+���GūKXz�T8d,H�l�D%���wٖI�d�Q�s̗91����}�?/`���\+��O���bc�^	�'���%A���'~ז�NB�L�0:4��L�8q[φ
 ��#9�S�,�/�4��7![)i���!Y�L!�ԙ��굼$cy)��4	�M������@���N*G�$%���������V'[��N�1�[���=7�P��RqQ�B˴�w������U�wf�; �@��~Q8~�LPIJޒ5t}��i�;/L}����&�Ə��G�++)����hM=7m��2a��n��fZ	�KʹR_�P��B����.��*����|+M��aڶ�Ɇ�J�W|�6��6����fi{������
��<�3K�-�/|�^�T�*0$��*��兎9�F[�̑G^�����쮞�e��P$��e��xIF	T����
���Ľ�b����Zu�B�DiH��jĵ{���sg117I!q0A�P���s<��Q2�W�/�+�R��3�w�؆˯W>Ti�gI���SZ����\Cn*�X�=�����Λ?��VT��OKaZJ���O�-��C�X���i��{�C��V��]�)��.�{F��=p̉��A*zp�~=�}9�"��\�҈�\,kl"�طo�F��b)�/��m���PFٔflݲi�S��R�Y������a����uL�8�vCZ^? �e�T�WH$��M��5�=�bN�s�6G�v��\���z���9!���y[�j#�mT�#�Wf���w��BH�WȀ|�U[V���&75�,�:*�
�����Mv�"��kC1�r�U���i�Ɂi�1P�Y؊��P���~������a���
&�#ΰ�4����q3V��I;l�A֣�>�Z��������Ӕ��gϽ���YԒ��y��hhn���;x���<�Bܴ�{v_I�kNN�e�e�쥷��'sڳ}z����Da���ko��ܼ��^{�X����n?���$��=��oi��ջ���G��]��&q�t��M�x��X�x]��VN���3g�`n.-�:��S��o���xY08�'�y�Ԣ�UKK7�a�PD(ij���B!��N�ZD����ڌ˺�a��H�����H4���~@q����x����Qw�����F��K	6�*��^��-Gg�e�
�q�̈́׬:�hm��x^y{���\o�S�x��O)���7���{]�yԐ]>p��ز}+#n�U�2.;�F�N;�w�#����E1����g���#G�i5�j�o|�~���5����u�Μ���a�5a�绰�ʭ����w�Ͽ�y�S���6�X�@�u�_����KXA��@�f�
�01Kٸѝ��f���Eu�W������tY Av�C\�4����)'���ĴRem���_|��tlV�t�ɒjF�!��p��ID�t��]���0&	Y,,d���^W�j{Ñ�i���U��8|�ѡ����� ����¼��K�x�}&q���6�\�d8��L��}���1uxH��T���Ip��Q$��fMͭT����`6�h�+`:�]��J��p��7dvaSӺp�5{�&gD����9�O��e���誻$d�8*����A�����4� 熱��1��M�i�&�lY���W���������M��Mϧ4�ٶi�R��,^��o��5�A��ШF�m�mڵXF���?����6΅�"I!	�����`����}����T��"Q �U�W!�����y�|�I�i���\����wt��O|��� 	���b���ʢ�H��Q<���úrrzQצ��u�t��Ν5&�אeJ%ShZ�j�nJ�Աpf)ʔgg�vɆz	"e��/pr�1T}��q�'!�}�W��f�8�l�5h���S%
T���YLS!$]!�_㴄�X!�I���R���5)��F��k]0�ɕ�\ӭz�tN��@Dz!�^Z����:�ךNf4��%قZ��hBK������17�A9�D��M}lH���/�wQLI��O�`eW���X�e�`&4?�t���$�3�*�����
%M���t�lA���}y����#!�5�4-.���P55���eE�h�mR�v�G_
6}j���ES�(9h2!.V̢�EsH"ǧ5��c�@��NDM9p|r����y�#dkq�Z���am�Mmt�$�ie76Y���2�t��;���xa1��(ܥ�$�IBV@�5�ؠ��Q��e��;��i��&�J*�-��AL�$�&�J���A�����46�q
J�T漉�kk��؈X���S�!y

�	�XR�x��2�h�f]v�6�	�)��G/m��H��X�n-݈֬7�ս~シ�K1/Y��Gran��\�.��ʦ�����̒ӧ%$��Mmz:�2H��k2({Q�$��Z0�.h��aَ�M'+���5c��Z:y]�m2D�W��*cKw�:�=�� \���K����d��ӗ�`�#K]���0�G�����e��X��4#S���")������s�.��ne>��j@ ������ڢ�?�����ځ�K������m�5���,�?귤F�7���c�r��8�3=�Y��t�l�zµT��+%�vŕX��KǚԠLbۇ`o��f�f��o/���kL%iB�&�4����s�� ���'� ~�POض-o?���75*Ā�L���9����7��CI�H��Oۣ�����g��?Lt�t��"9&\:���8n=<Ew͑M��{�T�.�X
(<zO���}WeZ^�\��B�F2�%�_�=V��+z�G��hj�Q�����R���\"� �5�j>�Pt��F���+,U}��ߖv4[�w�@4Ѻ���b�	P�kXz�L��=�pL:������n�4�|��ud�4�6���1���i�f�F�z�����=��%tMj? ��R�ݸ�E��v������my;W]�.WsW[�]����Zfg��$W�px�mo��R�βGp >;�S���㚖�_<ֲ�M����;��K�xr�x�zt������g�*`B}ǲ��"�l�SoYh&<�8�_B��j�����	00#���b�S�a|l�:;pvq���^��HP��k�ݲ9t�K[��L��%9�7Uߪ /�4���g��Y`�z-BҪ���*F`z쓟�W�R8�~�ԋ��\����&{aڿK�÷({����1;���=�����Xz,�R�]�4{EOu���+jLs �^b�wb��p��q��9-�n]ߍ`yN��ǃ94&���Ӎ��4��������-�plx	'�C���&�Rn6)��,��M����kTUs-/�����2
���߿hYK99q�K5��&@-��ꖴ�b�/
Ĕ�%���~)����gy��}�]#�u���A{٣/��1������z�_ɚv2p�O��u���㟿��&����������kW�$�kAea���E
l!J�Z[���V�+��v�ʘ�$�''võ�3�
�U
��y��O���zf�a�	�2��ݻ��?��;̈�Z��ru���6�])�H�j�_�i�c~ib���4��u}�x�\t�}~��$�wv�8&u��$����v����ޏo}�����]Mu��������מ���ch�EҼ�qK��HJ6�&���VL��Rn?+��Bf{@K[+i-�.q����u���=��!ݶ��b�:^��țǒ�-���v�f�$)�E��SOq*�d���W����TַN��9L;��]h���>�#��L��ã�L��n	��䙀��.q�����=��[��e����3%ۺzV���ٙ�b�Z���8�
�j{:��~ij�7cx$� ����F�>]��!72��
,�M�'o�Ys�Kʿlq|d��ַ���;E-{��9��K�K3�t,���* !
BH��7�z��b��W�֒��-��f�+9p��2���*�������&ym�U8�qvz�/�M�n4F���x��$ΥS��~��۟��2Nz�c&*g��M�㭣���]�ؼ~�9�lZ�^�_(�p~v�傁K{�@\�*�KR��J=�c�ŗ#�ΪZ�i{��
'�P.����(Y^���r�`�\-\�R)��.���)�'��8&0����֘Hj҂*mNNɛ�Q����Lp�>�{���d���s�ʊr���q�b� 2�0��C���C���k}B���߲/��c��(9��B�_���1�Z�v�d���1�d�T�s�#�����1�ڂ��s,�;��V���@x�b�t��ʥ�a�Pomړ�ǹ�
^�k��S7,p�/I�%�㐀.$G3�S49W�3��{���?
),�?�լ�(1���F!�B�A[���\QBy˩����:)m)�>fy��NV6��:LC��0D3+&�u�'�I.YH�q_�I���Q}�߹�s�|-���a�c��ߔU�gm/+��\e�&GKzdk6�FF��M���02g�r��?61�Ԓ��v�=�j-0m>�z��.�-f�0D�Ptt��<0-i#�/��ڨ����>�"@�m��^�%BN��$�.�e�&GG��i5�٤����M;�WbC�L��jD.��cd`b�����F�6�����D��)�8��hu��x�9�ŝ�,,�\��N&��/���ҁ1�Z�ď�P�
}�+���]��]�G���Y����6e����3ǎk��;,�A�B�dr���4�d�Mm;�iDz��Y�h^VG��*Bs���R���-ɨS��>�w]�G��O�,�'�cb}*��9Ɓ�c��v4vaK�U�;u�C���5[p��|f�<��Ggp���������V�cT߁�T���������5ZX
�G�z�Y�4��h$<Kv�qt���`�8|�_S�7\�.�=][����є��s�	�cX���h�����\��;�2D���f�=�HJMr���kE�.v�A���b�X���6\�ۦ#�Z�r\����F�+V�B�q\D��.ɧ9^N��*,My��t������c��̐�F�Оb|���\qn5���0��Z��͞�G1��,Kv/GO��]ƎUkP'O0��ذa:Ww��#�0m4�4ò��ZΜ������a0�&Hܟ��7gz��2rF�c֭_��V�l^O�Oq�>���K�s^�uB?�<�j��Fu\�W}c[����!ˣ�FbX�q�Z�F)�9�ۮN��!���KChڂ���D�_�Mk��V�6Yȥc���Ėh=.��ǆ.F���\��5�0;�A��S��nNL#Zߎ��,����Fkk+V�\���V`�R��.��Ag� ��կ����r�7�sx�p�w�������~��w/�(�!Y�{�͸^��W:]����z��X�����V3
�j����.��ܠlR-U4��7."����jH�s�X�$q��:�5��p~��X������1�c����4/^Dw�������Sغ}�&�����\ߋ]7މ�=�4M�����]������c�z��y��]͟yny�j���YՔ�(�3c�\�f<$P���
鵣Ǵ��f���r@Ot�k��xQ�^�?��lUz�]�Z�q|n�VMxYj���dM�7Kk$��(��}�2%��u�D�'��8����%�e�i����[��E�L����$Jo�\�U�;896����K���@=�1��ԩA���_yN\���k�
�*a\�s��Lb����\�_���"�G�]6N�#�b�4�M��#R-�������/�]]��8&�)��Xq
Ք��K�ӫ+^;�n[�>+=��4�ێ��柞�%��eT�X�[��jP�u�T��=�������"h�x���<��'i����}��5�*S�G����H����a�I�.M��61.AX�(��i�k�����y�{[��*�цM�@��<6�'6�\��ڄ2'9�y��E�r��*���Y�����ػ�@�"�E9�U�/�ONz�](ݖ�E㼇�`�cq�9*{I KN��-�~��ή
���Y�r�,�zh�Q�qm�6[������YJX޶aK�����V�I��*�V�݅���5��P���G�F��-�f����;�P�mu�j��v�9U��+���}�7�}��vS�,>�w����ac=�9�0�C�g)�!,�E�LT�%ז`L��\�����0���-m˚ٖrR�/�X�:/�ޙ��f)�f���ZF�_F����'�Yg(�D4����=�>
T#u�����G6����rƺ�_;�`p�Xƪ������O���	��r�4G�3sYl�hA�.��4n�}3#��:�unSMD&��\ZbS���#�~�Ώ��k�Ɵ~�q���y����gY;�c��S���ǆ�p���L�:˶�fm Of�8t�,���?c������r������ݤ���E7����!w�7D8 }S���C�}-�{V#w9�ӳ	��aW���4� '�ɳ	�8}_��w��-2�;7_��{�'Иh1�]ʣ8�Kr7�6�?��0�Ě�����8�_z�f��{5�[݆B}�I�^��\�eZ���G�Av�n����eܲm;��v#~��eD)�����ܖ���<^:��r�<��s�r���51L�����܀�0us&�pX�+��	xc�,�����ym���b㪭��?��O��lњ#��b���ï"A�H�+���§� ]m+<�`���:^>���"H"2��/���"�q������NE�0�����o�� J�Hq��PQ�j�T|����X׾R������r|F ^Z��B�L�6$�����'qy�V�Μ|-yBj��F17���V���^��D�kWa.^DO[&.Fjx��@ѩ���;q��k�&]z�0ͅ�=��ל�lӾ8t	��܅_��~��Xe�>��$?��Y�v"�+:z��N���0�ɒ-�o_H9�~P,h�������Zŝ���B�#Cصc'���O�Δ啪.�l���p��ݿ~� >y׃j��Ξ���spæ�����ȟ�v#�Y����!��X�x���y�Q�2eE-�j����-MXϨ|n&��G� ��Fa��u��%��8ƬUQ�gQ.P{�I�C..�\���HM5�PwO7yZ=�ܱu��Yʡi�r�C�u�����3������A��#���f=���c%#}��Ǥ��|��hѩ9х���BJ`*d{Y}��1�^����u稐##ػ��W���d����v �mعU�~�K8;pQ᧖$ᙷ_���룿�E�F�eFm��@��/m�u��}��c���9e�F���}�V��6`zn#�؍=���>�O"��j;�r�hY�����EUB}�F\��V|�+�������G�R@�䈷����I\���������	�����:k�l
�\��-�Q=�~�_�{�c���N�]��Or1K��xs@T�&��%G�������Ӫ{4�-�
���L�U`��j���1����%�L�:2t_���{x����TH��7��[=Xǧ���G/(�8�	A}���&�`"W����˙9|cߏ���%����/g�����ڋ�J�/���0ӶQ�����wg�3ذz-*|���q`�"ִwb���z*�Pi�y2���g\��m\��-���u��S�}UK�w_3���o�����AIȮ��NV���;�b��+��ۯ���!�n���?��8p�^8���?$�t,/� �on��={n�v��ꁗ��C�m�u���O|��ƴ����D��6C���5���V?a���W��ދ߼�n_�ۄ�q"EF���'ݷi�����J�W(��ރ���XZU�2L2>կ��R�UHy���x�M�ʬ�B��Q9��2�l�&O�<���T��6�i����y%��PZ�>q�}������ۏ�P3]A��O�������OᑗG)h6�Zd}�ں�~Z~�����.�լAn>��'O�������܁����ёsJ�Ÿ"t�|�}�Э��������W�Y��y�#�������]��%y�	���gP	W�{f�cq���?�=[߅C ����z�{������$��Ɨ��Ǥ|�ҲCt$�N�ԧ��!�Z����hs�A���s�țc���T�X�i�'p�R���ӭc��j9�_�@�A� `�������'�(��}��_��o��~�kh	��g�$y?y�X$�b��yWm�
҂z�	��(���t�/�?����a3�no}�vB#z��׾��]��q�/�o�:.�*)����lZq���7Q��bmK'���R���c��J�ʃ����ړ�qXǹ~��Ua|�+���V�a�	���<3�<�]��z�ů�'|�;��ܔ�Pb!Ao'�<\���p��NA�9l�Lr�� i�M��uupR)��k��#d0�e\�-8���W��.���
�oO(�<�����o��m�GΓȳ��(�}��/�r><}��W��]\�?����M-5�غ33�f���4D�\�j5y�W�z7��nك7O�Ã����ۏ�}�pӦ�hkh�-Ͳ_š#o���#������O�y?��ݯb׆uض~'{��X��Fӆ`�FO��"V��VF�(�U*�G�� ��m����x������I�v�ܶu3V�իc�kѵ���vL�L���_�Ƶ[�G�m��oEi���$�	���u�@�j�pٹN��,���n@c�ZLOM�.��S޷�6<��9�$,ܱ~-��t�u�]ь�.aCov0�	`*WĖ�^L^�C[�Z6�L�)��QM�q���'C�ɢ�~�6[�R������DH��:[;�Y8�6~��wcmc�nڍ�=�nش�Z���QЇ�A�̒��h�m���L��6�݋�ރ��y�'�c��[,�M�O�!�Ok��Rl�Ʀ���֡������ٸ����ů�Oܴ}+��t�]�d�m��5:a��Zݽ��G/��fZ�]�Ş>���̺��j�V����!�x���,/Y&�׶����?}�Yr����ꔃ��?C���-�>�	�&�aMZ��19�(��DKf+(�\F�I�]��-im��x��Y71�lb�:8r�pD-��~-x\[[A�XI*G�pq���@����~
���`}gZk[��A�fm9�UL]��N*����"�H_�~c�s�.N��������ӣ3�h��^.�˲�~���b�׀�|�S�w�4�j��ڋ���hm���ǵ�yf6'tM�_�ͫ6(DI\s��n�'ߠ�.��\<���D�"��x'9(���_G(�����{�T���9$�Z�ܹ-�98�Q��d��`W�p�zW ����WT0� 5erv��1���vpR�[�b��,v�߂�+����3����^.j�T��H$jQC��{��h'5���֧��p��>�ݗ��u�˼w @㝛o��ڃ����3����V�_�n���:H��$��9$g��d�7���u��m]U�{ZlI��/��4ξ8���I�
I;P(SZZZZ��ӴC��2e���3�2a(��!��Y�8m�4ISgu���۱�}�l˖,˖�{����M��{��ܳ~�;��/^"��q+v�_ٰ[6nA>y���I	����9K�I:���E҉�|�R�75#��E&���t@�Sʶ������G��{ �ե�>�zo�݁�@�M}�:���񳍏`��B�Rd�`p�,���I_�����	;&H�Z/�����OqJc'HUѕ�£؜���i��2�a�T����Q>g>�[�)�tæ/ F�ߛ�Ei�$uA�,ny[�dF��7@����>!#c�|ﺵXB��!)^�f������Ңqӝ��ʕ����#�s��0� �������b̢��*-E{{�Ћ��X����Yt�ǅG�l�\ܪo�kNc��rA2�ѕ�"B��|��	T�
a�҃�7:��H-��	��R3�C�:�΋G0/� �ω`|� ^;�_��јg��8���Q;�f�=8'�����d0砮��S�gd#��A#��]�� ���p������lᲕ���u�RD�mn>�si�k�Ԡ��Ӂ� ��<"��͆:,-���6o �Ǚ�G����()���|A�ѩ�9����2K}����lo�����%K���hk�X�����*���u�h�E��,��=��t�IgI�L��q�<��������=������t�Nl!:H�d �ͪ�(��qL�D�B+���!�[m��U|p�!i��xd�>	#Í�:�����&�k�#�-.���M�tw{�[�J@�ɿk�:�#ү!�t������l\kkBin&��ط�F��e|SN�ᫎFE߃d�jji���s��dȑ���}ȅ������� d��Oa����kp[�=��`�1ic����A�����7$����d�����<����p &�ϐ�|��2��c���$t���2�5DB�kM�?8��vR˥2���+��1GÜ=���xf�Sp�2kXԻN�8�-"�C����h����w�ZaC�Dvn D���v�N��N�#�'��"E�!�
~��'�������M=�����.��&��J��d��+Ld�"1r���cd[�p�p��2����x��\k��qm����Hjj|S�ݸ���f����%��э��X�LJVߨ���9����^ũ5�����{�¹H5�Hǧ-��(yx�>� j�l62A4<��l����%ݼc��פOQ c,�bu3Ej��Ps�Y����!S��ɵc�0�ߊb�i�+��p���D�|Sf�����'�@e
g(�ڪ=�B�M���q�r�dÁ���ş�����t"'Q��I[��,n�㊡=>�j
���}�����B�ψ}/|�yT�:�d�~�8.�0*m7�F����@}� ��!��/��1���>�ߍE�d�M�p�3�ە�Y�x��S�e̓x��]��f�e��\�9G6��J��N^��Y�9�<1E�|�\��-W�(� N':�v�����4CQ�3�/�'���;$r���x陙�&Ł�8��4:=����g�ō	EϪ���p$����s�Hҥr"P��{e
��q�������G?zR�9��
��I:����g�㡭�ӧ�8ԉ�,/���a��W�G��'�Nbӆ�b5y�!�zn]�Q��9t�-��ہ�Kg�g^�����T��G�c0�FFEr������^�9v�6�FVv߇?��+d�2P[S��+�!)����)(.Bь��0���1��^RDv��E�����w�~t�)v��ŉvӎJO�\����^�g.���%��9������v	��0�����<CW�i]K����pU+ә�Ț���E8�^7ޯ?��7��G(����+hki&��Ӈ�!�������g`��$�
�Q�����~�>�a�u�k�S��Ұz�z�ͤ�?��l������T/-��=E�m�j������n'y^�X�zz��<�o��;%�>��ީ~���x���������݉@_���٫*�Y.��� �E�9y^k}�ś��t���"�Z;�}{z.Љ�d�?C�����N/^������H3���[8K���j�QL�$�=BQ��M�M�n�� $�����+m� 9�.����ӈw�Z2���å�N���c��P�T���0x�����[���B���_���*�����ϖ�ۨ(���N؅���'+��hӭ�¿u���_�}V������ 9Y� Us��^|�t�W^�0hW�WR�}�!���?a��ش|��#�i��9t�'�
���n�蹅���K�D�F����t�R��z�am�2��|Wv]T4�q��$��o�ތ���6&���K6�?«�����2C��N��VQ�{��L"T&�z]��j��lR���c�p��xf���'�����]��9�MS�I�h�E˥.��H5��c��x�67�\�KA��B�4:�A4�V��������d���t�����2���ن�wje�0�Z��N�e�	�ǉ��t�+�᩹���-���j�I!����-C�bCL:!�iy�ZZ).w�*���/��\2�7xp���W��R&��@lӈ
U�PvE�ƒE��������&��\��J��y��0ݓaRR�c"J����
3�(G_��5B�������JSLp����CF%� ĬN��^�!�J���V�����b�s:���f���2O>�u����a��M���Lp����vu3Y��f�"0��EE���ʛ�g,���h�B���T�t;���D�d�&N�ڻ�����,���54�����+�t5�n�0�B��	���©4����T���fD�ʝ��&)������-B����6�ϗ�åB��df#��J3rɶ� ���C��%Ver�o�F*|��)ך�5LC=v�6J�&��i�/�p����n��iX�k�0V��v��0R�� 4�v�k�@�sɘS$Rp�6`��L}��;h�)*V;��h9v�F5�$�A��;����#!dQa#5�!P��Q�@փk+R��f����N+��@�75��1?��w�R�Q�ۊ ���}�+���GE«�9�?�����z���A-�-���J
�'��i+��%\}'�m��Ҩ�5^�Pn����h�Vئ@е3�Z�VK��ʚI����܂C�t�s�+���+�N��F�[8���I��NQD_�R��p��co�E�g ۝��y���ݢ�e�$E��@5 j�#d���`�,�2��LxTB�mZj���$�������oL���@�x0`Z�oM�ѵ��	yN,��M��cKA+껰V��S�	B�.e0�i�U} �_�z8ug��$�sl ��⥜"��*X�+�q~�nr�2�����8���M�x~�
z�:��!4Dwxﻁ����)[\Ԅ��X�n�Yᦪ�Y��哛���#�}�)�r��BK��\Z��ٚ2����k
��Q�)x`C��M���r[��BN��ba.24r$��X�~Z�l)65U���&8���1Ik���՘�3C1��*NE�Iv�Wc�1
�ʬ�(�g"	��M���Zx��kiqEV�A�й�~4��c&�i�(X��$�=Sy<<ʛ'�	�-�)��9M]sA<����$�p��U^כn�<�q�'�����Yݲ�]�e�&�P�l�%�	)М�6�
�z�d3Mm]�Ko��wI�ֶC�'�!-\W������.ڰ����ڌ�� �P�nڃ�!�By%n�R    IEND�B`�PK
     �9s[��4k� k� /   images/fd3ac6b5-800b-45c8-a4ce-2476671127d4.png�PNG

   IHDR  �  �   ��g�   	pHYs  \F  \F�CA  ��IDATx���`S���w�)KT���T�Tq�OQ��P����7�� Ȕ%C콡�����ۦ�i���M{o���W�����m����;�Y�������*Y�    @��Hiu�7&�SWUA~�����;{�:    X3G'7v��{e~����.�۰i�T    `՜���V�c�͞���>l��-�    `S�&د^>�K~~���J��    `K�"د]�~ha�"v��m�7��    ���>�ϛ7ϱX��c�_�G�]      [$�`������]6n>@     �J��>f��Qi��/X���J̖    �%�`�rɜv�%E��/�H99�    `�d��-��_h�Z�:v����d    �u��111�E�V�;p"��S     2�ʂ\������w     ��U��Y6�����,�H%%%     �d�Z1�YaQ��E�~S���"     �C����z(��������	     *�|�W�T����{�|�]{     T&�`�|���iO�X��     @?I����z��L_�t     �'�`�������嫶�'%�"     0L��>&�Sג��u��8v�"    �q��ʂ�o�]��~��C     U�\��Y6�մ�̧-�DJ��     �j�
����w_Aa�G?.��rr�I�|}}��ݝ��ƍX�� ruu%�JHH��  `���E���(v��mNq�)$E;v�o��V��~�����������	 ��֭͝;����H�bcci�̙�  	�����SOQJJ
����'�`?o�<G�}Z̮?����4IQ�N��P���FR�������ѣ}�����HR6h� �=�= H�=��C'N>���)11�@�$��Ҿ�r�F��� )��H�6���~�m����ӧ}�ᇒ�����5k�= �)���1HW��5�f����yq����3���ݻ#}r	����#�܃M��>�@8�dذa����{  ��:}��Y��]E��y�l���l���z�>��c�����۔�-��9<<�
E��0r���������e�u�������QXXX��1r ���H��h���kT~b��BQQ%''@M�Y�����,�[����n�.'���}��7n�������iڴi��=F��=��4c�!4�:p� ����TPP@R���O�o�Q�q���ܻ�K�۷7�k�����^��{�V�kG�E�'O��{H�ߟ~�)-Z�� j�N������N+���L�����<��#4g��W�<y��_�������὾poj=���7)4H�uҋ~ʠ�;���t�y���t߾}��+�Paa!I���\_�ǄZ�����B_}��0P���?��5��N�y����������A���/_:�𝋴�4髓`߼�����Ծ+cv��<��c­o}������^zI2��uYk�wqVЧoQ�.$uS^�����yP�?#��Н+�g��0a��B��=��]�r��^�m۶B�Qnu�|�r�_å�����%��>|��y˿�ڵk'|�ȑ#��!>ץ�ZO<� �|�z�_�d΀ܜ�ɼUQQ���j8p �M�;ҷ�~a�OJ�����p�줠�ߖG�g�v
z�@J�L�#���Ț��^˓&Mһm۶m�-q~��2�{ �Z�f-[��������7�r��)S(((�>��3�����.t�cyyyB�T��U�VB)N�z��'����Pz��W%W �W��>fٻM�J��%+�(R�2HJx��w�����?~�dG�tYK�wtT���ck��������� z~j��"���3T�ζl�"��K=�k �H_�|:.����cǒ���01_�g������5y��θ���;q�I�s��I2d�p\!���{����X ���`���=�U%�6n��u��U�>�8��}�{�n���\B����=�|�;!��v���`�����S�i�t#�����7o.�;�C��݇_<����:����)55���_h5����߄Q��byܡ�@�������%�qf��/(33�|�P���%��s}zup��� ��ȹ�ˀZ�l)�0U�{���bͲ9O���b�������{g'G�̝_`���5��M����C�������73B�ٷnЭ۵�n�Q�F�`����^\��;;h��ɼ>����ł�=�f����ջm�ƍ��[oY�ի����%˝�� �a��;�I���|>���?�P`` B=T[����s޺�z{ಕ[IJ�A�n�s(���b��za~�8:���@O��r'���G7S3).�]��DW��$���Y�e'�Z����N�JR���/�S��d�:s^|'�r�-�����K�}���������edd�M��\q�J�P����6�[�������(2��$?�J�oFf.��ʢ��T�t5E8�����P�{����G X��\H��'z]�;���f�`�j٬��g��p��Kk�f���6a��#}NNtw�Fԩ]�:x����Ux����5���cW��_�)'�fo+V������?Iɫc|�ޞdMZ4r�O�ѫ�%�%����U�Y�(..N�p�n��2׎jƋ/��HE�=�>�r�J�={v�����#u�>�G����G�^n�[�����kK!���>���������]�/�s9�= ���ӓ~����>�|�}��F�ѴiS����Z�c��)�!�����װ��V���n��,���\Kǥ+5�����(��@rsu"sp��ѥ�wwS�{��=pF}�a�����.xv�T�<ڗF�&kԩ�+�H�|�wb,��G��n��򅜱֬�W��^x�����Ϲft׮]���ǅ�]Rƭ�j���NAw����[���y�/����ZR��Mh������kt�r����P� @Mq���
���ڵ��9O��9\b�s�N�X,�/Z4ݥXi���=�=Or�믿�(�{y�Ҡ�Pd� Q�GG{!`�n^�V�;@)��d.��I5�?7ć�<n��^�w7w��Q҇�Ŀȍ��Z�i���O�
���-�M�6	�Մ�wo��^xRoMB���y�>��/����h�>ؖڶl@�>Hi��_�����R�='���*�w�u�nݺ�{��a^�_��Ϋ�[�K�ł���ӷ�/�wذiي�_=�;y���s=(Л^|�7��� ���H�dX?/z~�ق�}=)%�XX�VLj�v�k�U�V��>}�Ї~h��Ay����]���Y�c��7��L/Z��>�|5�  ����ps~�Z0�X<Pd�$b��s�=����
qY7H�u���,�c��~�Vz���ne�. mڴ��8߆�q���{jX�S�������](v��t�tY�$;�?�%/��+qE���x��j���a��p~��i�2�i㒜~��Uk�k�s[F�&�c�¿��A���s  ]\%�u�V���f^O���_&�2�c�d���I�D�+ˁ��>f��{KJ>]�t#e��%t�҅�|��J�o߾�N�}`���ݢ�^�ܓ�;j�a�/����Τ��/G7p5�k��G�ڵk��/�(����`��`�d�װ����O�G�y�; �4.��U����+t4���V8�q�%�F�`�r�`e	���v���kId8S�P��8I�'�%�H�������8A��''�P��G����9�Up��ꀿ���2�,s��œ��C����pכ-Z#���/Ƈ=������J�q+97��JAA��E����Q8�C�BM�8pp��=���yX� @�g�}�Ya> 7���-�ϛ7�Ѿ85������M�պ�P��B�{U���K.\���8�n҂տ&�ۧ��<��|߉l8����h����3���N�t�^��j�>\� Y�׷�^.�GIz�!��;�L�����Ϸ�522s�/_IY�̧�~X�Q�=�����t���A�|�ݍ^)pל~};
sf  L%�dV��7�=��$$$�G�`���ٵ���׬�wW��V�{;5�r�sO���x`ٲߍ�{߰� �N�۷�;��~nլ���zϐ&ѡԬI�=�zݪ¼���f_�|s�_8|�py��^ƶ���thU�~��%�����kŊ����Z�rS��������z�7�lZ�~c?C�[ԧ��&���j�b�>�x��0�!J�_�t������,�d��ۥ�n-+LZ����ɫ��[�qXu��e�����ӣ��ӱm�������܅D��U����M����G7��v9�{M_���%�5\]]������/��|����-��Bu��q㿹D�>��G?nߦ�\Wo������   ���K�U�J~X�|3�J7�Ǻ��J�-��3�ϩ�q{��-Z��='�G��9��>!�>BG�KW���s��UT9��W)*m�c�wq�~�U��5m3�YP�5�6�ˉ3q���_�i�K��j۲��BQn��w0� L��c"�(]�~����(دX1ǗJ��~ݴ���k$��������n����,,��ϖ-[�\
�:ڵ�0zr%ܸu�/d}����-����<ٻIth3cߋ-�
!^O�/�؈~�?!�S�_�|��{//�j�+ְ��n��F�~=�f�?n�W�����_Ǽ9ap�������6�� `��g��1f��ӧ�9��V?u9������4h@�����0��]��Yc���A0>!��I�&�II�O6�p�Pǜf�Ék�t�V���J�~Z_��zP���5_���v��S�;v,���&O�uss��>6??��]�&���yt�Z��b=WRJ�����PIϓY��   j��`�<����i/Y����]�)4�������.ߺX��[��tP��)��D+cߏ�y����}���JU��C�B�_i��|R�7ܷmۖ>���8q"ݗ�n���jҤI�c�m�)7���gx�����+bwm����ܼ?(`��FQ�zg�
ߏ����N)#��Tg��^��w5Y��'�qxA��0+��,��?7�`
�,[PPD���[�V�~��!�s�gd/W������ �	��8�kz��
��!_��G��:_�P9�K�իW+|���
�}���&�j����S�N�5	2ޞ6-=k���y�v�Z��Iƾ'{ i���J}M������V5����A�Ν;����;��0U����%���(UK��ܪ��d�u��~��^����9�TvߩT�����F�Bm���|Ⱦ<���&�+��W�W�}P6@��XS�o����)Ő��O?	#J�����;���&S�O1���!G�;�֋���wޱ�?��JA�j��ϙ��?O��`���@�6m*���_�~��uG�u?���#� O�4�222�|?~<4���� ��V�����,P�ۺ�/��'/��rs5~K�@UxD��\�bKf���*��\�꺘�r�ܕ���-�)���U�XY�&:й�PR�ˢ(���ڗ~��E�w�(ߦ�����+�\���Qz�ɷr۴iS�צ��/*���ڹY%���Kn�9����R�.M��Q��\�8��*��o�֭�_�~@x�����~�v��M�ׯ��k��
��KgΜ)�Zxn�F˖-�n7�k����/�m�6�AAAԩS�
�EEE	����煁 �&���:0)b��^x�����m=H��裏����V��1b�:zT���J���W*��,���EE�`�����I�+�B�G7�k>���J]zO!www����/��=VVs_q�^�x�������>�F���5Ǐn��R��p�g�����Cre�`�\),*R-߾�"8��[��z���	��6<���9.\�@S�L��5�b᭷���i��׷t��?��s�z�۷o�̙3�$�?���4l�0�]	5w�9�/X���n�J -&���߼��=h���l���>�%�'��CI2O�� ��~�/*�����)��ꕚ�3�/i��=��������K����ݻWy7))I�P��>�����VW�\!�*)6|�89:*��!�~�Q���jrs5|�]P��/ ��Q�E����_e�1��������Էo�j?��5kݺU�s�BBB�7ިr?���#�|�`/=&�U�f=XPX����6PN���«Jn���x���mI�`?fLW'��
��Mkm(gz�gyiΝ�z��ɯ�>iwʑϨ=�	[;w������]n��s�/��|���9�{����;y�� ��믿ґ#�U����6TyGS���_�/^L={�,��d�¿�O�8Au�zx��v�4c����;�<��._�l���݀4��;%`�*�}̒(I�*f�.�����[�F�{���P��I��+vy�؂XU}O�D3i�bm}Y��rUi/r!�+U�{�Z~�|�<� -�x;OWg�gH�`��������u��K111u���2��c�ƚ5��ￅ�����(��FF���E�]Tvʵ����/�n�W)73��h��eP���b?����PcۓRn���3b'�+UF��:�G�Tou���W��{V��y|}<�cl{R��?  `��{W{�o�^K�v��;���Fr:�������3fx�qKVn�^��5��vQ�[��e8���"� �=��T�ʷhde�Q�,�-&���k��U�W��|����ް~@���Yy�a  �0�c��z1#;���J�Ŷ;1Ӑ3�{�0��=z�߳gO�V��#8�'���p�޹7l~B�6M��HDV0p�����k��'xq�\�9�@��m�wߥ�������3s&��td����FjlϜO    1�����O�R�����QF���nW��W���-�j��x��"��={�^���~���Q�F�9!�%P;�x�	�0a�h�k׮�ّ�W{V?< ���[������0�џ"�ۇ�   ��R�_�rV0S��{�/\�')�K�\���.�\�3r���xjռ��}Z4�wϋc[�݂�O��ό�;�m�����F�m�|5�@G�ұ�]xis��^􉉉5>�ڵkI�RR3�¥$jbp�V�����cK�_�q�9���G���e�'��s-.��lso  _�`�k�t��xŚ���k�苧���B�[]���)ux/_�Y��ZG<����g�Snݿz�N��c�upk��u��V5y��='��K���H�(m�#���S��$[�6�2.��Ug?��#rpp=5j��{Ћ���'�QT���n�x�6�'��x��Ԝcc���XzĈ�^~��[Z6�oUs�w�W�  ��
�>9���I�=V�l'�w�9���ҹ���G�4�I�qs�)�v���v]ӷߠA��|��gDG����r)ʳ�o�]��Y0��c���V��FQ��T5�[~��gyA^P�W
��e��O�E��B�2�_��w����y<�2�v�+~ު�����{�z;��8*�io/�*[	?u��\Ca  O��Ϛe���������P{%-r�#n��NA��F�sws�k�&rpI�rpttHZVN�����x�JU��d���� <�/��$Ym9����Ȗ��KZ��v�0_­HK[]rKҚ�s�f���P!�{{��\Ξ=[�b"�n��0��}=�����j߾m�(��;*"zhjv���}���빻9��6�����\�u�   &!د\<��J��q��-���~��QTTB+���<H��NU�oooG������Y3��V�; ��E��
a�*M-���?�P�R*ȎJ�
(��[?�
�(�Kt�F�5���ܜ2˷�-�����?� �{6o޼:[�E�

�h����ܨ���\�M2��mP/ @�!��7�9�w?g^���  ��aŊ9��Jպ߶��~�4nӛ�{P/]����äpPJ��b��i����n�=��W�?�Sp�/-��/������j�:_���~E���#�
��
Y|���o)*���d�֭���_��|�V���F�F��13�梜ˀ   ��`_�\��ћ��6}Mpg��w��!�����"�QXT,���o����4�S٨=OeVڕ��+�����}ݯ/�W�zͤ[��+р���Hs�Υ�m�
��R�o���p1�qg�E+w�ޔ;o����V�/ ��
  ,�Kq�n�r�s� 1)��Y���LQ���'�r��6}Py��l��0�΋uq�/�'aG����y_��������h��BɎt�Eʻ�K]�t>疖���)??��4��S��w���R�pQ��p���� �JǺ   `9B�=F���u�V�m#��m��͹F�+,,�=���?�Qq	V ��#�kF����p��|i�UY���cU(���ׄz�}�l�رԿ����x�JKC����)~\�;�ݾ��ޒ�\kv��(��?N	ݳ�{  ,́@t*�9zYhgש}����Y�cdf���c���_�)�쌪P���M�Jp�>���^�׭��j�������]w�Eǎ#�>����?�ȉ�ԹC#��.�|}ܫu�@�V��}^>�_  ���5������QtdE�� O��v��'���ʹL�V�ҕd�wSPY���*�p�YuV+�<��15
�R�j�*�ӧ�г�M�<���݅��`��������/��mP/@}�z���[��n_�v+�����KW��z|� ��!����q����z���Q(��=K���n�g�������;T����r�?y�$M�0A�Óh�����ӬY�l���O�>-�1��/��Mw��	.��aaa  `���iӦ	��{��!K+(��@��T�o�!k�	���4�\�A�>z�S��B�ㆾVj���G���}�����~�СB_�)S�Pa����̙3�222诿���s���۴iS���O	  ���7oެ��/���^}��Z	���A��`�
�թ(%ź��W���6�U�rc���cR�k�.a���5e9}��>��_PP@�B���N.?z饗j%�׆F���4]���l����  ��ܕ+�[cʦ����Ӆ�{�=�Tx���_|A���:�ܹ��o�s��Z]���_&9���~�tCթ�Pp�S�׶�~z�g���'ooo�=z�w�}'�{���5x��7���֭[Wx��=�Y���?�$9����������˞�IѸq�h���  �t�R��w���`�=��şKTtý���p�[��>44�-Z��6�ƍ��SO	����ڏ�{<�:~�8�5J���Ν;y/��ef�=���,z���{^���k9���
�o```�mW�^���~�RSS	  @æ�=��p�#�
�իWi[RR�
����9D7��ژ���|I-t<�+�#F�k�Y�6m�r����,[�L�k�����/��*m�~��p��+E  �f���Y[�����N���+m���?�<��ő,�9�ڷt��\,r|)���8W@���j�xŘ1c��?�q^~���#GJ"�3k�|�e���B���w�x12k�  �@�/c-����W��ѕ�ݺuK���\��+P�k�'��S�-C�+�&SNn���˵�\�<`� Q��}�v�k	�!!!6}�i�^>�}�c  �ƜAX{-r�<��C��P���.ܾ�x�"I�������Ǟ��X�Ur��� �R/�3׼y�h͚5  ��`�C����ˋ~��jܸq�m<Q�'LJ1�kX{���PoK��|�[ZFEEU�&��9  �.{=��===�P߲e�J�8�p(8u�I���{���%�p��s|�����b�  H���.�'v�ԩ�6��}��$����B�n�a���B�?q�Ʌ��{�������wnp����%���3�#��B����  @�����&����"V���-u��Σ���\n�%�#��-.A34r/�E�4wښ4iRi���ĠP(��Ύ  ��~��T\TLP��͕�����#�����>�΂}��]�vz�]�|�Μ9Cr%�p�P/<r��]�-�0:th����Oo�;w���H�B!��� �Np���P�� �T*����߄	�n����+�P]ٿ?M�<Y�Q�w�q`��J��p#Gr���1q�D��>;v�Ο��u�V��nƌ�F����;�\   0��\��/���޽�^{�5*,,����_�����J�m۶B���>+���r�������G��w�o��Fo��Q]Z�v�p�Ξ=�*�:滄\���/RNN  T�^�&MV��g���4eʔ:<���̝;W(�֢E!����۷I�8�O��B?�
�&�N$U�!�K���=M�>��|�I��ccc��w�z�K��M����D���܎���\�  `���%Ρ`���z�oܸ��~�m*.�ք�?��C����W_���s�m͚5��K�
���͛$G��:S�pG���aԱ���+��np�������z��^�Z��u�R�e��B㣏>�t�����9w����9  �{-
�{�=0`���j"������{~��nnnn��j���������w�ҧS���Iړ�4�@���M��:�w�>��cz衇�n_�`�ЦV��m�FB�-�;o<gf�����+ײ:  �<�2�Bʣe�z�һ]�@��&�~������^a�j����7���$r	��u�;���*�4�OD嶵R�eu�Ǐ�[V׼y��93��  @�=�����d{��w�\B���Ç��=w��A˗/���z�H���5�kߝ�P��%-���;��������"�w޸�nɒ%�.�  ˱�`���h�Ν+m�P��'���ŋIn�9"��sW�
���p��Z��ő�5�k ��///ar��E�xB�̙3��3r�+�r7�Ӡ{������{��y ��a���C�js[H]��ʕ+-��v���@v
SQQ���q��)�=�q���������\�~���s[Y�z����Z���U����/M�:U�sI4������M�V�ơ��6l��s;8ؓ����A�R�/��q7�3�{�-22�����-R�� ����t�牲�B=w���7�G��� �ES�z�M�n;���Rڭl��J��$o�%5��,��s����p�w+���GR!����e�5j#�7h�@�����x���z�sKH)�i�B=��兩�Z��NA���QTկ�OA���Z��=7��RӲJ�߫|���ra�]V���Ya[Æ����z�\�sI��E  �ʦ���%����=�JYS�.NԹcc��.���ܪܷ^���v��M(/���B���̬�}gϞz���;�����KRam�^Ò�>((H�h+�k2�RSS���w��	O>�Q5����NM��]Q���Zž��vg�½�=�('��+=�sj�r�ѣG�nW�u��~  �ͦ��><�_�P�#|��}����ټ���PѥsS�8���`��S5����E�f7&&���ZC��%�=���
�3�<(,�T|W����Б�W]�p/՟}�{�i����.���R��`ޯH�#���f��ƴ���{��?���q�._�  �`����b|��h���Q�pqFP9d���9�jV�V�|�n$���.11����C����!��믩q����'N�F�ssk~���V>��s�^��w���oݺ�䠦篿�������BĹ�ŵ�|�ߪEZ�v?��f�},���   �"�0?zHwa�]l8^�Ů��N��f'stj��AV�54�~�G7i�?�p�/�С����˗�I�b�zƵ�<q|ڴi�J�<)��>�{[���`>���wٌ	
�q��������7  ��EcG�NN���+�N:<��n�==q������l&�kp��y�[��}׮]��<'��o߾Mb�U�5jDÇ�y�v���G�ЈA݄s�R�wÈ�])旃��x  ��������,�5�~���:Qnn����?[�`nܰ����k�����a�X4�kpi����K�W�+�R  @L�5ē�?y�ɷ�
�T�7��s�/�ĩTT��h�������\e���:ӷ��� �p���'��|Q�_ ��q9�y�
�Jx�GG�wW����y�\��'�C�����[k�1  @�}��ٖ����O��.\J�1�D5eŊ-zg�����9|rT��)�A>F�cr{���D�V�&���u,�Uz<ګ�0�*鷳/]I���՜�{�d�ۧG�.��]�FG�����b�x.��Ꮄ�}   ��N�������O�~�P Ј�=]������i����nݢ� �3$:"�Z5�O'�X�dZ1��¾mkX?�ڶ�0����:s}��s�ٳ���:o�C4U}��n�O�ϭ�7x�K�i�4�G�����   � �`ϫ�6o޼��w�K����7��x���?,��lu�;s&)�6~zd��ڷ���X� ���xXZ��@o�1��;���y��#ǯ|�����sܲ�G��{����0vq���{@�  �H>��B9��9}�44�ꊟ�5oft�g�U7�k[�|���vh=�P �6z<�g�-��zsB���1��:�yw��9~�zluC���˷�tvrk�&�yC�����t5�&  Ԕ䃽T�ժ�p7���Ĵ�����y~\�y���Ӭqx��K��{� ����LO�
��4_��Ϫ�1��vm"�n�r-%����y�-��¤�lb�f�m��   
{35onp��\�~󕥫��5䵤�f�ot���Qo�l�8T�å���(�&�W��P����*��J���֣���ϣ�7o��n�iX?�GG{���wɆ����  �������D!�>�'ܸ��t��Ub=߲5����>޴IX[}۝�),ć�o���PT)Ы���zh�����4��q4#�R�xTXX%&&�~숈�F^�����ap�����˷m��V���7,��b��F��{��P`�7���   ��@�7CP���2�Դ��b?g���e�wmm	��`_��F�(�J�q2:�XQ�eo�{**�{)�ݻwS�޽�9(?���5����E;��!Chذa��t���|�����A�缕������`  5�`o_O��ss׈���	���C�~ƿ'k�/�k�J'�k�W�p�W�n���4���R��o���'�{�I��==��3��S��z��Io����qII	M�<��;F��������<�2��3+7�G2�m��  � ؛�W�4�HQtD������n�tww��;��Ŵ�o�Nw�^_�Wjz~��'��Ԑ��TT�Ps�d�J������{��B�/,,�	&��ŋ�v��Z���s��֭[kt\777�����̙3iǎdM�\�����-��W1��\�ީ����A�O�����  `Y�fp0җ��AQQ@�%�7���H��m341���J�H��?7o;S�^�����c��������C!�Q���lz��h���B=�=��#���/���kג��w0|���o�^��z��_�:��}rckU   �
�&f(*.1��ßCIr���b?�����a���b�%��z��^y�c�9�F4��%:jϸ���^�+VP@@�h�]�z5͟?��Q���G�ǌ�d���b>���d���l������_  �{3������ҞD����suq6x� /�����|^68_9���fvU�H-.���iܸq4m�4����N�<I�f�"k��k���/�k�~�K��z�w��Ά���U�;  ��fH��mt����p�;Q'�z8)��iiYd�4���u�Z�^Y��ڇ�s|~�}�U
��3gΔw��Ro?W]�&������K5��   L�`o�����"6�(�>�������~~C�m��"j値U(á;�����*M�/�J2����=X���wc}���������mOJ���  ,���E��t��������̈>�����7|��55��K�J�iuɟ)�G�}*�@
��%;'�n�fPP�������G�5r�����x��Cz�nP/��������n�.   �)��t�l��`�"��۷�7[�l�q�l�����t�8{!��"L֬|�^��V�S{ԾfOB��2��'�|!� p�A�V����ik�z�����u�\  ���L�O]�^��6\����<*���5y����[al��'��-��N9�����]���s%$$X]���ǯR��Z��盞�S�a��<�K�>��a��c�9q�   Ā`o&�}~�t�m���>͚������~3�W�٭v�|v��_�jQ��}�o����Y덌?��\]]k�N�8au��'�������}Z6��}�3���~��'�y��zda�5���	7n  ��k`׾�Բy=r0�b�M���'Mx����׭�wٔ���7�������SU}��{N��o2iWi�����F�����&�B��N�	��k���<y6�ZF��v$�rܑ��

u�ּI������{N  �X�k 5-��:O=�knt�F!a���}}���f��~��4>`@���>��5����VeC�������$�u
EY���0��
���.�/ݿ��ԠA2Ղ���S([���5�kz��M>>>d�n$��_�/�=ݯIth�za~q>��ϸ��֪u{���oȐ���\�W�?����pQ}��'����T  �}��{�ESx�����\�w�n��:X=ܲE����܄⢒�)��<���CB�}L\`(3+�����:�*�/�sUp�/}P!l�铐�deeѩS�Lޟ۳j�Ϝ9Ӥ�iժ�U{�m�q�jdp"�����k�&�q�R�x�&�YY���E�)J�O���C�:ȇ����s�+�v���  �	���JJ��z�za�C���R��:C�}=�o�ԟ63�9��K�����j�L�W��!�y�����p�Edh.���J�4y�|d_Q��R����s�Z�EŴJ}.=?�Aruu�r�y
��j����9���rW��Oy��   &{��ے�{����ȞE���B�M��/-�)M�&�
a\�>/�g��%�Za�Ғ��DoG� \j�({���{�v35����KO�A�Ύ}���Z�O(  ��Hn$ߦ��v��!�����"ϑ_PD�~�O����:z;;^rV����ޮt�*��?�J��T*��P_�MQ���z�%����篧�e����2�?  �%H>����+=���OR�r3��Y����י�5#1qK<.���JSO_�9��W�����\�	��ؽ=�Y�Vq�X�h}Y���+�ϵKsl����;h�=,��ۚ�
mr  ,E���ٙ3gH.��
iy�Ԧe�ӳ-y{���x����?��X>tB~Y�no�	���@�*ߩ�1e	^;��i�ڗ�|E��딝�O�WZGP�ښ4o��߱��}�ͮ  �G��^�xe��g�]���]4���V��o�g�?G/ӡ/RAA�~��T�����l5Z�R�q.T�=:�/�k���V��*,@��(��}t�]stq�>���$L�  ��T\R"���[P�5�
���)P����k�D=~���ʣ�i��&��s��*��/ou���z^�������?Vy)�Bq��F�q��z��������d�i��ԟ�\ނ���qt(5��O����K}�:����Ŕ���>�����W�19  ���'��[ޙ#%5Sx;���
��֍[���e;��}��c�L�--�Q���s���7Z����b̘1�裏�֭[ɚY��M��!������Ѳ{  @��u̚5�����҉'�6�V(

������Qy�K�ҙ��	��h���+��+*>���B�9?%%�-ZD���?��_~�Ν;W+�W[�oxx8}���  `��Z�lM�:�6n�H֠Q�F��w�QX���z�R�9Ze9B/��T�=�o�X��w��������i��ɴk�.�mڴ.��w  �16�.]J�[�&7���k���|@4���Yt��E�sw��[�������[�+}�^��N�U��i�����Ҵp�B�={v��>����K���h���$g�z��?�Po]QQ͛7�   4l:��޽��.�����
۸��Krx�{ʔ)TPP@r��O�;Ｃ�67//O�ܹs'ə&t���k�qS���y�f���F�*l����I�&QTT���{B��Q�F	�/��#''�&N�H���#   ���4l�0�;w�p�[W�>}���u�ii�X1�/J^|�E��D��7o
��'O���7��&��^x.�����o���͛W��������+���۷I������>�����}��E  �f���q��!<���c�U�΁?&&F�R_,�G�y0w@ч���q��ƍdm�ø9�S��og*i寙�HNN�ѣG�G}D<�@���۷�U�V�K/�DW�\!)�2"� |������2|�.�A  �]�e
���]�vM 
��"��KyR�)�ꫯ�C�z����4a�I�2߱?��=�A���j�����RҋӒ��B����ҫ��*��;��v�/Ój�|�СC$Eܹ��<�h�B�v.�����|  ��^O��ɤ<�ǣ޺�4���m��$%���z��[���}�]��9�O�g&ї����Y3��S��t�2���Hx28O�������~������	�k֬!)iܸ���P�*�(�I�J��   A�׃'�q���o__�
۸��G��ی�jv;w�,]|���_����I���)�W�K��p/�PϸΛ�ٳgINbcc�I�򽼼*lspp�iӦQϞ=�	�RѵkW����̙#�  T�ހ#G�А!C�Q4������\��[s��c�g|Q��<x��*����Y]���;Wq��.+��  ��`oDBB�9�>��Sa�^N�nO��S0��p/�Pox������м�╂y���'� �� �W�'�rk9�4�!A�Ƙ�g�w ч���w�i�4��{������>�,͘1�@r�����嶖   ա�����(�F*�~�:W�L��[o�]�I*�;&��KOO'�:vV���ҡ�'vRm��.n))W���[�6���Tp	�k��&��U   �P6��������5I��q/{�:W�5�����p�M��^rv�ӧ����@orr�h�Jr�T�>�Z4t�����^"�s,Z��ڶmK��{�s���-[�L���Ӟ={��   �p:j������5rh���������@|��B>��$w~�D3^>:%N�sEno
�w��Q  �VB�=�=��̜9�~�a���Y���   �W��Y�{ �ؾ}��f����t��ͤ�Y�x15i҄   @*t�A��B��222L���   �R��%�=�x���=��_c   �Ko{�{ q���N��/˷�(   ȃ��)�jki��);WE�cn   ��]y�j�����\�3س��PQ����lZ};   @u9T��=X����>~3���7س�G�R��h�z�{   �� �,��NA�N�{ڹ�-?Ɨr�nk   �ɤ`���^�C��N������?���оj�[��駟���   �dr�g� ��Q��������T��~����   X�j{�pPs
�N    u����!���=   �ͬ`��̇`   b3;�3�{     i�Q�g� էR   ��j��=@��   �&J�g� �C�   ����=�i����}?~<�X��   @�D�L�G�C��/�=@e2��t��1;v,  �<�����s8���=�=ԊLE96>��M�/<�~;W>YUU����*����`O����p��8    .�{6xĔ�6�:4#�׈
�e�\CiI'�`_�Fe]iTz�:o�8+�ݭ4���:؋� �  ��,��=ԵK	��t���h��&k��B��@
;Y�+%�=   �͢��!�C�ѓ�vvԡS�j&-q7)�ǲS�P�c.{   �Ń=C�yQ��Yj!)�z   [�{�pu`�R�yeY��Jq�  @\���=ȁ����^e��\)   ��j5�3�{�M��r�.:��{   [�{�p�V�Ӓ���    ⪓`��A����[pT�    �:��l&�  ���4�3�{��ܖ����    �:��$E�	���   ��D�g�`	��g!�+,7��\   b�L�g� 6���vlYY��J��99٤�S�o�T�G�   �I*�3�{S���M�UB�^Q�?VR��S�--�����7��F�1y   �&�`��A4e�4<ϩގS�Pz�
��eK��J���,Y��\   "�d�g�Pm
})J�=�w��oǣ�����{MW�b �   dB���!�CM)4��v��8�e#�L�RT�_�s=   ��$��=�T�@��8���BU�5�˪TG��G�����   �M���!�C�hFޅ$_Z��_U�����
�{��o��   ��d��=�Eqg�lYk����|_R��8    #�	��޺��׾�C���/�0VQړ��즪�e��Ŕ�Qh��D�vTڊG��   �"�`��W^b6)�k콲o�$i�J� ���.�Q�C}����l=J�}��   @\����Cԅ�z�H]���8���"7j�  @l����K7L�����C{   �	�{�pUQhf�R�қ��
${   ���=C������{�
��&��[2{�`.   �>���^�f}�J�������Q����
��    &���^��n��S��wC�1Y�W�iIt;KI    b��`���)�f1�{'�v��M��   ,ɪ�=C�����b"+.;G�   K��`��AJ�  �6Xe�g� i���   P+�6�3�{�k�l�F�  �Za���!�C]�/��    )V��=    X;���    ���{�p    �ʦ�=C�    kds��!�   ����`��   ���l�g�    `-l:�3�{�����   Pl>�3�{�����i��|��g.   X�}�{�;;͙HӿH������FGGSϞ=����t��I��ӿ:|�0���   H���{�{u��9!�
mٛm��_�>-Z������瞣nݺQAAA��ӣG�3g����ȑ#)55�   @��u �׍'�x��/����������*ڼ�r#�������
���;w�����:օ��z�P�7o=��S���E    M�z �׮���1�D��;4r��>>@����̞=������y�}���TRRb���g��5k�P�f�h�ܹ����SQQ  �� ��p_;���	O���Є��"�~@�	����5f̘A���5:fBBM�8�,X@w�}7}�����믛}�    ��`o½�u��J���}��n����p�<yr��7o�]�v�r���K��;v,��Ջ�N�J3g�$   ��* ܃��?�!W�ҋ���\�裏D=>����׏���h����n�::q�  �t ؛ ��k�SRRD=f~~>:tH���o  H����A.��%ddd   H�}5 �[�	}5���eg��+ذaB�����M��  @��	��r�\�J��d��h|"���������Ua��<G;�myyyU�ӨQ#a�R���������)�  ���`o�{�pu'���g;�Wz�ù�@o,�kF��������)��H}���ڤ0�VC˖-��vvvB�{S��Je�ˇ  X{3!�ˏ�\��Y�VA����0˺��T�O�&M�?�e��eU���	   �����A�uC���/��z�*��d58؛�  @��k�^4�ޔ�xaE��IVǎi�Ν��~�V��?�z{Sxzz   H���Ae�1�*՝���(�(���0ُ9��m�FG�ջ}���F��t�"���/<f@@ �w�}�   H��H�%J3y���Jg�^���������zꩧ��͍���i֬YB���dõ��Ǐ�𘓓͝;��N�o߮tlggg�ꫯ���G�<66��  H������5:s��ҀnbJ��8NO<�,|�\:�$$$�G}D3f�>����iӦє)S���W�}�����^�{PÆ����{�B�wuu�/���ڴi#|�c�z��r   ��^d�W/{���zoK��晐x���(����>#��5;~�L%���ެ<�޵kWz衇�����/L�MIIF�۷oO~~~���Sk֬��^��E������-l��v��Qxx���СC4i�$*))!   �{:j�k��>���z�쨔��"��Bv%���Ttt4EFF
�s0ׇKtƍGǏ���Lz��ׅ�������#�T�����B	Oaa!  �4!؃�P���	�Q�z^uV����٬�,!��X�B��OQQM�8Q�lѢEt��M�9s���׮]�^x����	   ����Y�\!{��e�Y||<�3���n��9�sY���7ұc��'�j�}}}���@������-   iC���C���sH��^p��U�:��℉�    O� :�L_VcOh�   2�`V��\�%8
�<Kq   �6!���Y�
   @�t����Z    �@�    �� :x�^��z   �{�j*���>�w�������p�t   �`V-",�\�W�R�&Ö���,5�ʪJW�e
����G�U#��79���V�m߾=]�~�>���r�
  ��@����	��0O�0�>�W���,�(�(���ή4�+x�L��ԩS�G>�������OEEE   �����2�
r~��:�������CY�W�z��)��c��#�w�޽��4���s�   l�=X�	���7�9�����$�
����   �{ +�p�B�Gc�ΝO   `;����U�����ԱcGa���͛	   l�=��8t��   �	�    �
 �    X{     +�`    `�    � �=ԩ%?gR���hC?�9�JZ�5�    �dCq
���#y�Ɯd�dJ0ق��6;�N](���=�H۶m����ڬcxyy�'�|B�6m����   H�=Թ����OShٌz��d�

ա~V
9�o���ׯM�<�
�7�,X@yyy�>N�.]��Ν;Sff&�ڵ�   @��Av��Ky�*rw��`_T����w�nS��~eߛ{3n�� l(-�-��Mh!�a�e��� F�*��7��a�v�#!���ݶ>�G:ґ,����mY�u�d�9�y�9�]��>�"�·M7ݔƏ/���h}!R�p��駟���ߟn��7n}��'   �`����S�0ҙ*����5��}z��M7�x#��׋�<�w�Y���]z�4x�`�f�mhҤI"�gƌ   �����$u�.�eM���R�\t�E4d��x���t���WY���3�<SD�@�'O��;��͛G    { ��O-���Z]���i��h�=���s
N��{ٲet�嗋}4H���N˗/'    �= e����QV��Z����{��?�Y��s���?�\���9��Yg�6m    8@�>��H�)5�[�b   �`��ፏWS���������#�P��Ü��s�x�xy���?gΜ�엇�   @p�؃�p�_3��_O:�t�|h��貪w��E�.]���;577���/F���   6{P<��
Z�,I��)�,\�I��Z����𓆳�[Xi5k��&͜93�6����/    �؃���SW�M,˹���o=�+�   ��� dt��5�:뮻��xĈ��۫W/   @p��2���s�ѣG[���}Ϟ=	    �b@�8��C饗^��!�E^M��d�M|���   ��� ,Y��z�c�<�H���{=��ӟ�D��	������{,����_�Ýh.\H �?}B   �b@x�'���H����J��}���X���{��/���;w.���i�m��4a��4M��s�g��ٳ	�ba�G�l @! (������N�s�����|�馛��O��ǌCg�}�c��������z�t����������կ�n�=z���t���o�A    { B3��k��ͬ��Z��/f\������s�=Իwojll�L&i�ʕԽ{w����"8j���    �	������ԙ?��Y�����G���,�Gu�y�4h� �7o���������#    �= !c���Էo_�y�=_����NR�L�>�ƎK�\sm��6i�?��"�    �b@�����~�ȋ����E���(7�{,�9��Xc�-�3o�<���/E~=    ����c�/_�<�mX޿��;q   @��      @�     {      B �     � �      @�    @M�3��-��[�n�b  �*$�I1�  �˜9s�L�������z4B�    @m���A�Fד�i�     �0 �      @�     {      B �     � �      @�  ��v؁���  �?�-[F�?�x^�@�  ���w�Y�   ��ﾃ�     E �      � �=      ! b  �����[�r�J  P8�/�{�=  ����k��  ���      @�     {      B �     � �      @�     {      B �     � �      @�(#C��x<Ns��)��F�A����p�B    P�؃����k��;��k��>��>��#��}���׺3f̠�S��ZwԨQ���S]]M�2�n���b��=�\:�#h���4f��駟    @�a�M6��o������k���v����_��WY�k���t�]w�H�t]�	&�}�ݗs���S}}�x��f�Q�l�喤i��у����   ��=(;[o�5�z�Խ{w��t�҅���:M�#х�����F߾}}o�b}��g�mn��&!��xz��%*Y����o��d2i-�W������Σy���_n���_�B?�0M�<�   � �e��h���V�SYX��-[F+V���L�nݨw��ԳgO����Xͯ�v�m%=�m�ݖn���of�ܹ�駟�����q577�卍��q�xn���b��q㨩�����JJ$�c�������o%��w�!*���C��#�[=�����y�AѠA�跿�-�  @`�؃�q�G�9�#}ժUt���ӓO>鈦z����O��O>Yl{�)��ԓ���*�~�s�=ž�U���C�?���"�',x\p����cN-���T�   D�=(9,㧟~:{���W_}%�8*��w���H2�Qe>�`���R�G�3q�ᇋN�\y�5k�8�o������>���m�hCC��"B|ꩧ�N��x>��Â�Vp*γ�>K   @�؃����ZR��+���f�r�,h�͝h�=��C��������W<XY�9%(_�~�m:묳�t�m��F�.p�(��3g�
    �bJG�y�Ѝ7�H����<���E��Yg�u
���_t�E"O��k���������k�ђ%K����    @)�؃�p���d?�v�B.���~1<����V
�ϟo�=w�    �&{x�������R��    PM � �����1���ŋ)��6�z�`�    �&{XxH��.�̱���?�jÝoyt�^�#�����X;���L�=�pK	�j����t�R   ���fe�eN��������&uuut�����k�w�}G�<��ҳ�F��v�m7Gꓛ���_eZ��K ���&l��-i��7���P����jÁ=I>3���x8o�o�ܹ���Si~3��b�0s�5�Іnh-�1��<�̒LPU(C��������O
T���)N<��رc闿���mx��K/�T�� �]�ҟ�L8�@�����t��>%_�<_�}���3U��H󸤼�E�u���n�����ӧ��]G��NɎb�_��o�=�5�F�AÇ�5�\S<V��u�����կh�����7>�5�X�v�Y�r%�p�	��?(;찃�����O�7ޠ��
�z�1�P�޽����/}��G��O ��<d�q�ݩ���ϸN��	J���M{.=��k$�*�> Ȉr���{��Gs� b1�bZL�C�|����]��2��{�9��sKr�{P5x6�q��e]���?��**χz�5)V6N;�4��/��k���x����f�ԩt�=�P�~��s�ؿ��;���?/�}衇��7�|�����6����cb�`��D�	C�-����R�ʕ�� \�p+��E�2��x�jW X���}<7�MѧY�}�݇���O+�p!��jp$���5-�G�s�y2)��/Z��"��#�p���;�Ǐ��Y�f(-|X���;ebƌt���Ӄ>(�et��U���|����@�=�@��
���S�R�2ߑ���b�H&E�����΋{3���WI�Q����>ӑ�r��5�@�^S3D]{̖�8�R�q]�K��s�z�~c[�f��v������)S�:f�=�,no���ȥ紗��[Ot��!.U��ŭR���^zID��X����8�{�С��8��p�I'ї_~I�p8�.'#�<y��q�o��@r��裏�e� Pu�q4b�p!�	C��'M��Q{N�R��*/��t��G-���+Q{�/7ľ.)+�q˾��k�_ϼ�q�O�?��\���c�؃���n����������;ҟ��g!�οg��O*!�駟��W^��m��V�~�_X�x�Y�e�s�˙���F�����7+R_f�L����Zb �-�|��D")n��#��	�z3GH�|2�rdJ��7W$�;�
�o��z�k�\G3Rv4[��5C�㺺3�3m�#�v�B�n�阔��<aB�����? �����뮻������z�%�G̩V��| ��S:� k9����&�d{����577����#G��0Ýb�s��7���Ջ@���_��5m+��@ ����)����Z���ӌ�۷��'e�ތ����j�=����#pJ�3P�y�.So��o���转��k	#�>u]ǒ��#_���o~�უ�g�q]}�մ��{SP����/��V�Z%����Ξ����d�������O>��ϟ��{�0��r����[�G����[���?�׾�:�,Q���縘W�1�k�{d��p㍭����~##��7��uU�M���z�=(:�jv,�-��y,�Y�H��>�0�>&;ך��ܙV7�>lxQG����௺�@����oQ�=zd\�%��9�<�'��\�SN9����k_����M�\
�����ӛo�)� |���0���GH���h=��i ��>}���6I��,G���J��ݙ����0��d��=)#��q�;9b� s�ˤ����ɰ=�Õq���� ���s���\?>���c�M����̩'N�����￟�9��r����:JTTn�����d�>:::��SO�[n�E�=�~��7<�p�/N�����γ����{t�}� �t4�}����v4^F��w��c�˴1�	CY���N�q�����Y�4�UI�h�L��H=w�M$y���kqk��sժ��b�G�9�|ʔ)E���FK)�����D>�m��F�W�.j_~;�r�O��Rβȹ�<�	��{�����ȼ
���������� ��B"n�Ȇ[�y2+�{Ns����(H�_�V��
ڹ�[ՙ�/���;�;�;�ޖz�ػ�b>p&㠿,(Y�?3�ߔzcHV�^��9��s3�c����}]T�"/X�=(9�n�)]z����n+�Ӆ���b���Bָ��3��8O�>��}��֌�~�>��~:]v�e4f��afQ�m�ӟ9f��<~����_���ʺ�+F=z��袋.ʻ	r�-�̹�[�w�e�����HGj�[��w뭷Z7�l�dd��G��(�����~�̙I�L{�s�zsXK����z�1��E�%�$�^�zE�y�z]�� �2)�=���dZz���Y  ���v����O���c�=�;���H0�쳏cy�N����B�7�xc1�գ�>*���%e�s��x&M�$�+���^���ܩ���T�#���p~<G������9r�-,��W'��N		s��Ӕ8����8��}w2^k��D��dE���<����x�wO��'@�>�,���Y��3�/��])�cd��D����c]t��"�ʺ���j �\J�a�I1I�f�ZS���[�u{�'ym��u	bJΧ�~*�Y懳�q���3l����l�]y��bX�yB+7,�2
+�H?����L�Հ#�\r���se���{�8�?�0�qq
W
T8���SO���{�M7��by��Ư�k1�����irJ������~+���o�-�&���=��k�l��t/�ׁ��<�U6x���k���=��#ZPx4nq���E �?Rl�4]���N�)F��� ��b����k�Df�2{�2���*��C�AY�v)�,�G�Yι�'G�8B-�u�sN}���8�����E���	�/dmU�󞣿�Ύ,}��n`8�����E���i��i�s���H�ﾻ#��p� W
�M���%K����}x�[���p�'�xb�}j��s�J� �)S<n���^Kp�I����9��+>|^8e�+Gj�;)���9�ϝ���g�yƱΫ��*^ �57^wߒ��Tx�^ӐmʏڙV��$3�ٙ�j�2V,��C�A��xN{��
�/���^���l�2�
�Q�L����s9�x�Cr
Y��nˑb?��Lkk��'�|�
�#�K�.����o�b��RϢ��
\�#�8B���J��[o-n~�:u�H��[�U�M�&��$�Y��Q�:"�����;�>��C`�(=Y7e��b�؃���矋��W�|.������r�Z���]��K8�>�e��|k���g�N�9���������;�иq�Dk����W_��o�����<<v<���3G����+�^r��_���u  P~�tF��zZ��i@�qw��ø��z�F�(�� �e��{�Ο/������<ZG��|y�&,b\pm��F4{�l!ʹ:<r�5�����/�R����O<q�\��θ,���#��E�|r�;W���lpw~-)��w�)>���Y   �d�(=٩:�b*w|���Z
87��8
��>�j����pE�o���s� ���2��փ!�;�n�c�+O���    ��Mǌ���Qǽq�Ɛav����   y�}9J���3l�2Pw6�a/�џ��/��   ���Bg��D�Q�  5���[����)e�bB�:�,Ñ5�c�>�jt����:@��αw�T�犆؃P����N��o�YLz�����i̘1�s�~	 �U�^�V�u�q-���ˑ��   @ՁÃ0"���H��b   ����N��Aδ ���a�*    ,����YU#�kxo BO>�{   ��jD���g���PR��4�   0�#����4hР���y�|��c�$�zB*�9��  �4�F����o߾%=��������P�h���=  �H����<�+������G<�����mD��/ط�  9�,���	WGZ�?��2~=y�>+��,��  �,��L��u�1 A��R�=  �HP��VK�3�o���a@^���s�  zT!�Qm�	B.y���i��TJ�ϟ/:��%;�[gGi�<h��@L�G�����[z�  j�лwojni)X�}�	����Ƃ�[�r��|��	T�J*J�@�  D��c6�fϞS�����LK�,�>}�.�҃��7{   �%ӏ?G�L,,�Ps�����.\(Cr@X���{   �$�464P�����m
���R��\ JCm~�    �= �b   ��\r� �@�A��ի�9���ٳgO�����[lA����?�D"Aa����F�U���۷�����q����K��� ��2@ރ	�I��ȱ��=(�n�-�p�U=��cǊ[��Ŋ+(ll��Ft��wW���k/q�6��;͙3�  �$��k�
��j����b   2�U�ʕ�������;:&Tʱ.�_�^r/�o�g�b   TD�G�^y�$>�\�xM]��?:�|�xlɽ�|��Q���[@�A�H&��j�*
;�ù�Q��X�,��ݟ�(��됝�!]
}L>�{��X�\�4��烮�^��1�'�1� ��=���=��v�3�믿NQdѢE��;R��ҥ}��'@�@Ծ<�S+DY���X̸��Y��s)���/���y�O7�>�䨡��+���C�  �;Pb2��˴y�ٌcR��
�bC�+/�ħ��麙�c�}��[��kre���6�@�  ���~�XB�DjK}]�OI}�\f�h��!��ZL��G�uq������ד2'��i����C�  ��(E�!��H�ф�ץn�uu���cΨ��|���lXRoF�Eڔ�'�I���ä�	�e$:��t �     >���R�ެ\��.8�L��C�ˇ-��Ui�t��9���n{#z�GS�!�     >�beg�X<&��u�:Z�b9��ґ�4*Tztc�{   ����('TU�S�x�ȭ�R��{��4h����^���p�B�R��}(��J    (!���f��������uu�DR�����Sb��]
έ����>�羻���#E���  PS���Ѹq��/^L ��S��1�c	OT&���4F9D���>L�h���n�³�kbd ƜS�zl>2�5�s�'��u�.N��=$M�՛��h�=����1c��|���:::�f�����fGY�,YBQ�}�;;;	T�$��{�Ȍg��↎��C�E3���cKOx"���v�y7ek\^Q��gщ�����E��ݺvM_7�:���w�y���o?�K�.�L�?��s��9nO�XE��  3*�R�B��c�6-�m)��RR��D{��v�7D_,�Lձ��"�N�q���S�7+ο{�^T��G+Vo �    ��nL{J讜�~}�S}}�H��L��^�g�53�I�k��^�ٗ#���EH~�3���   B&�*-~��SQ�z���1l���Ï�G�wt�O$��v$]���J�Y͎�Q����z�b����y������!�     y ����}y��TWWgE�e�y������֜Z��kim���Vjmk���N+�^b�=ҍ[��J(?Nj��8UAH�S��	M&�@�    �b:����E�e��Ï�x]��%u�))v��ň���w��®��*��P���m��,G�;ĠF4^]��Ƶ?����8IQ9�V�	�=    @4름��p���655��b�"�,���"�<iF��M�cg%��C=��#�Fed��T9"�{L�4�w����׼��ܑ�(����    �B�xn��ɝi&��X���9��!�W7SW�H�-���-��U\y읝I1�oRw�LHԿ������n������DWQb    PFX-9�#؝�VԞ�q���Qb�uo�a�g��}�gg�JL��N�(3Q���ђeK����s{wߚMV�R�|�
N �     e�'��aX�9�<�C@�ܛkP1n߿_Z{�5�q��D���n�L���ͤe˖��$^>V�k1cr+���ѪU+i�m	8��    ���=�RRςo猓=�;��<+�k��k���G)/(�(�_S�#;�x���}��Q��aYU���9�u��K/P{{�x�+�Hb�Bc�F]�kgj�QK,�G5���u�Za��=��JJ$q�A�����C��4�O:#�F�ɹ��:ݺu�79"�����]��t�����]�И�W\��,�K/�������:{���6m���V����=����7Z��n�t5u�������;����~��'N��U�H��e	��As��o�^M�d���šZ���u1���ϧ�Xa�Ck��3�;����S"���[,.^�`�D�M����h���z�@�'��҃.:�?�j�����K�����/�Gv��/XSR��kS�it�m������4��A4rD�%&?���<�,���9�h`�I=�׎=�>�ѥ7/��~� �9�&I��c��h:F���yUWs��<���ռ�����d�ӊ��K}=566���Q�Rϰ��~Š�������۱�M�l�j�S-��.Ɣ��Ƚ�[՚�3��[��#��~���~�]D�.�����>��L�!k�Lu��b��B��q�f�!����j��%��=�W���S��״����?ݺu%��=pP�R/1�u�o���1��}-K�$��9fvݡ����\�$]�ѓ!�1)��Z�����i�F���.;�ڝs�bXu�����Kٯ�s�(�C����ԃ���7��Ǜ6�Q}����Չa<�? ���֥^�W��$|����K��}��1� ش��QkkkZ���jJ},%�����3�&uR����L����d�Κ��뎔���ٕ�R�^ePF�a�׌�iE冋�z��c���![1d��x<Nu,����߯�@� ,R/�%�a>&�܇I�%��>�瘁�\X���ȣt��{Q�=�f��۩=u���)3�)TNP%W��x�֚	��'s��9�Y)8��f�J1>��S@M����vO�I��aObe��9����Ē��T �=��K2�}�����0J����S�$�瘁�\>��qs�)fu:xPJ�����FcL93m���g�Խ\���N�r�'z)�^ϰHw�n�\�X����ߚe���m���}�	��KXh�?�N�ؐ�(��}��z�qc��=�}T�1��V�觟������v�v;+����Fz{%Rʫ%�G�-E��r���H�)�������H=�U���L�*`��@�#Lإ^ҧW�n�b0�|�R:���57�e����Sn������'�����]���s̰�?��J���V eě��Gmmm���%i��tvv��-���Ev�]�=��W:�)��c�7J����(Q�zI��q����5x��(q�nME� X�!�����<�Kcc�x̫q��Xk�FOj9#��~��Όu�]&�V8����HI= ab@�0�u4F�!�C�x��jE<?��[o���_��!��MK`�j�zЬ^	�g����S鄨}~@�#�C�:~� �di�����5޼�����1�����ۭ��5i��i��zR_ {    �"Ft�b"j��bV�X#m��1�%�9|��h�Z}mW[��>�T�{ ���B�Ɏj�  ���ec����H�#��I1��X�\�=�����)�>���/��8:��#G��4�}�@�AE(�{ǽm-	o�ʭ��7��S�*)��i�E �h�MΠ*�ni�I9ּϜ��C�3-���U�}��wA�y1�8��<C��A��r����^�B �A(���@ ���Y�oD�E���e ��=(n�p4+�S��/?�{0��`/�*��5R�b��V[%�Zn �?I6b�T3��}>��S@9�؃��I�U�u���:� �$�Z���zp��K���ˠ�̹*1~p�˽,H������� @�X#���ΰR�SR�'��qd��2 �� ��������kz���rF�ZZ�}��H�^���&����Tf�_S�d�h�̥h����8����Ĉ�k�5 P*t���#�h���=()~��^����H�HF�ގ�#z�DW�3�U��Tn�d�y
5=-z_�2��⮨���UqQ)i�����  ʃ�m�҃2�eE7#n�5���ֹДsT�mѵ�st������ev����VˬVj�侚��*am�l�Q+kծ���%����|���r?Z �/  ��bAʕח)jm?w
��n��Mhʍ�۲3�<��W[�T���d2K�s�^���J��{�=+U撵J(�1���,x�^�u~��b�ll�d  @�@�A��ZS��ʱ|����P�����ˣ 'S��r/�#(R���R�I�W+6s�{*m��D�)�퐽!������V	�m5[vŋ�i�ȔV�Uf���(W��XI  P�@�#H֔�R��[�T��&�p����V�4�h�)���{w��d�X�E�*�cR�ZBO���ߏ$m���^�QU��/�U�qW\��>(��I��Z�<��n�����ˈ�(��Z    �=(3�%CnY�D$[ț92�+|-�72���Xʽnڐ��TS�S4t��ˊLң̖��"�F��^���)�V��QݴJ���&�ʚ�*a�o��|��JpټD��6GZY��Lһ̌�JTP����
  ��bJ���$�|[�D�9���7�=xHL���:i�!	RSz4;���OP$H��,_��w?���k�t	�L��2t��I��i�=����P�+/��Z%T�����]��V������z�j�y���R/+2vK�3��Z�FMTb��'U��y  @	��G�J��X�E�h�'���f۝��>>z{2�1x:�uC� �D������Y�u�_�O�>����[��Qk~b�cV`t�����3T�,ѩ�Mw�W���FIQ���cԵ�]�r$+l2��N�^ie?-Щ3A��[})2\��t@�$5t�QLm}�����
   ��M����J�nK�����]<f�'�QzwtW����~��Q���}ﯱ�Ί��h��[eU�6�c�tD[-�����7��k���s��f�;��z�f�|�
[P�e~��Mh�-v�^��y�~����h�F˽����
   �����(FޥnG�Hg@�4�H���l?�
~Z%���ԍ6�h��]�|9}��&"ݚnG��V	^�J�?�~�z�Uޮ�fR�Ϛ���_R�e   j�}��$����2��*1�s��Zm����F�s��~^K��H�+lK-  P�@�A�)މ4�_Rv?�\vL8F�t�������-��ɛ�)V�no�Uy��(}Q�V��:�y4�H ���k8���m����rI���؞�)��z�O%ڟ�'   �<@�#�^��^1�ՠ�s̚94��-�KKy)�%�^�V�񵐗  @y�؃���et,$gh��B��]e�ր��)�#[�aj��k�3����}>�ۇf�+Hx^�%�g!�   ~��G�J�Ɉ4�� y�b��M��)�ֽ�L�:H�܇��[O(��3-�e��i��gFN6Uо<N��s	   @�AYQ%W�
��\M��'_ѤW�l-j*M��3GF���)]�)���絸�#�\�����J������b^-��   ��=(	j���D�F��[DV�")��);�$ɨn�9�M,�q,f��\.�_i�uTb<Ҭ
#U��ٕ�@S�
��l̨�i���Vf   ��Rɾ���ƨ��xGn�S��B�
Ma;����ẉ2S	2噧�Y�oys���T�J��le.�#*l1�\���b�k���::��˞�yjnn&��A$����K/�I�  �bʂ��A�Ф�M��5uk�W�u��R���4�ޱĊֻ����l���-I��Oj�b~Ԕu��x��+�ZR/_?�ԣ�u�%;����<*0A�ش��C�Wiv���bϡ��������K/u,{뭷 ����A�iӦA�){PrTٕ��H��a��>�9��Ĕrk	P��6�=?�pdm0�sb"�I��2��gE�)]��!�^�㣋�tZ�x>����][d�M����iX�NKp�s�:�ՎX�2�k�u���Y��Fy�װw��.]E[�"��V�����   @�@�#H�b{n��B�{1�)��-�Cʽ�ԫ�y=�&��
2#ښRn���A��҄>��V���RP4s�#��K��\{v֤�|*}_V�Z��Rq��xC%�*���������z}v��JEM�������:+n���  @��e#��Y*��3^i����~ ����
�%�f��n��g*�5���_w���W�^�#�V�D\�'crͼ��U"��׊�[�)���En�R�\eR�.��#~O�g^�!,YE��G�r~�#�^r/��7)�^�����mRS��I�+]�Yn��ܫ��,�W����dk��O��Z\w��
�g��2��A)+ ����;Ĕ��ZF�u;�%ˣ̾@ ���d�{㉴ߴ@n�}Y�*���T$�Un��܏�8 e��*!��i����$�Y+k�s�Yfc{-�2�� �b�i�5R���ӧ9֔i}�6zV���C-��p ��,xɽ%F���]u� �^�"g��,��G��"j������H/˧��I�2P.���;"Һ�$;b��:�dҺq?�li6�k�L���"����+��'g�od;Hd+�����|�W�L���V	+_'}{q�V�Ld�ЈYZb<��� @��y�՚��;�+�L�'	�fʽ���o5{PV�t�#�����r�˥>��*�����5F�y�Uf��kQyZ���@��U~xM�,Ch���Y,�dʽ����N�LtR�#���H<(�=��h}���a-wTZ%$^���9l�v��X�yX\#�O,��_koo�ztttPGg�������V�}TPS�@�@�#H��'���[���*��(� P ,�)A�ҥ�u�����j�H�[{G;���
�g�oO�D�ތ�g����(�b�� ���V	-1�D)2_,.Ʋ!Ƶ����	H&"�����-������-љ0��k��u�_�~.��.a�� J�ח��aMknd=pn}�:INW��o]��46t��F�K��mFn}�έף%a4-�u�C��bA�9�D�g���h>D�:Џ��uW���(���7�r�*Z��,r�Y�F���9R/��d
�Fk�<��Q�=  �P�W�y����b��ߤ�B�YHCA�����_��V	K����h�j�6jo7r�y4�3m�*�Y��H�)�}��? �?�Q%bB�j�.ԣ��V�\�ab���������ya��ƞY�� �i�dw��(���5���1	��
+�x]��>���  9.XX�R/�ӧ�����d��+�jNZ�+��u\䪜Ɋ�kr��ې-Υ��������et�U���  @�hmi-J���.&�������X��|y�Γn�GoN%����NRIi�.;���3����4k.k��<v�gx\(��C#w�#W�=F9X���G�` @�ɖְj�*q���\�}��Ґ!C|�뗷�~��M�������
�' |!ǋW��r�J��z�H��3�]\�Z8� �Q~3�^�p�<�߸o�����B�{   @!W�3K�iu�B��}�R��k�t��+�u���o�}�C���~���׻�me�hJ����py�=-a���ޞ������}"Ʉ�  %�=��n�P�b_ʙ?�D�����x%�{���s�׊f^;|K�t��$V�sJ��t��Z_�ה�d?��H��"��5������"��3q��^ �� ��\ @4�#���\g)�^�b�3�兮�GS��\��N�P׍q��cq��jb�Tz1HN��3֒�ڢY��Yr�v4�-��?y�;�,�J����k1���fc���9�FN'＝���5�c��@�b   ��jPF��b�)�M�qo���a����;�,}]<)d�%7�ԕu3����DJ�9���Q�K
��TN���=�Nf�*��ԹӘ���7n�hOI}GG����W?K��餄1޿�#�gbE� d�3��|��ɵ����޶�c��6�4��꾊�������b�)�Is`��w\�h!��?м6��%݈�;/ig��W�s_��<rߪ��p��D'}?sf�ϚU�I&i��b���#��b   ��3�O��z�g����Rҽ{w_�A�k��y�X��.TϝB�a/��|�f��ET��Z��T���-*1F*Qg2A��	����\M���]t�]��g�EY.o�ٓ�<�\�:�5�oߥKZ�hM������  �����i�=KI)%"S��j������9s���dDύ���/��O��F�x)hf� �ŷw�S[K�ͦ���J7�$���T�[c���F�E�7����S׮�Գ�=�ܳ��[n�8��
>�>��r�s/�
?��w��Q�ܻ�ϔ_��.��7('��-:�1���Sb�G���K֞j3oۙ{ݘ�-i�񲄖0�#�ʦV�V�c؞'@��D�ez�����߾{�.��NQ�C�AE����jɬI
-3��w���7�>�����-��C�ˋ��ԞtVwXyss3}���h�7��򂘒��:O5w��o ���ԣT�E�qT=�H��Ug"&'����Br�������װ��+CZ��V����}y�744��ux:E��!��"[{�E��S�\�@�(T�U�RN/���X�Hf:��w+�)>���{_�߷���a9SI���)�^��h��������b����Ǔ�Hp4����3d��u�Ҥ�Dro�׬�"����J=��"�ڽ~�
�T���/��^����r3Ş�Z�X������t��u���D�Ant3Z/o^ttv�SO?AQe뭶��/�BD�9R/;���z�B�9'��z�C����Bu"��uN<��� ����I}�O]Zv��]��߳r�Y�3(�.�wf��J��w���(�x��\��׭�p��� �n/���=!�]E޽�4&��/�����ֽ֙�ݡVM�Q�������Ip��������Ϭf6�y�n�%7c���޸�l�+#��}W�ܙ.�|/� WZܔ��^�Au��dq����.%K�.�}��ȑml���Ff�/���:#W>�GJ�α�5��"N�D_Vj�fM�+��}��H�����	E�=(9�(������9��X��3.���{I}�J�3�o�)D��?����Y��.U����w�Ž���J�ʫ��4�Z�*k 7RH�v�J#F�(i��믿���ISVu�f�G.dʌ���~�a@�:��Th�.�)m�P]��p����zF ���d�zUnu���9'�p����
�q�R�%iR����23�+��� V� ��&W��c���\��UB=��Ŗ9H�5�?��Rl���s#�Dޒ�,[�����a}�i�*?^#LeX�^�U���]��ӌ�R��B��+r+{ѫ��Cҕ@��4ۙ˭H�)�A�]��z����擴r+��I�+)���J��(����{=����л��kA�kHx�����!T�YV���	8������.�nݺ�>,�;��>c^��|�O�ñLt��я{P2�Sk��r��m�Mi������NэI˕�O�U���
��Ie&J/w,f7U�����*�E�V	�H��������٫*�e�)v�+P��s.T����nk� �䍩���7߰žĴ�������G��	�%�;�k|!�gP<N:e�O[!d>�ݤ)�^Q�jD:sUf��'����-ʩ�sA���X,]�U�D�m� r��(���W��W���ΚV�g�ŽWy�=���"��D7?�B�y(�DBo	����ի+�~r�[���C�#H%.����S��DiRd���%M�ٓUȘ�W;�>[�E�uS�~��3�����M��*s��� (D�Z%4�5ƫ���n2I�u-���l��)�q�*4 7�zTjǰ��[BORgg�@�q��V5�=(	VD3�����E�8������i�?����mꠑ�;m�5m(h��j'a)}�Vi4}V��4hN����e�n���Z�R�e��=�VXU�
�o�m����|Z%�|r�3��V����B��dR/�̢��ۧ��V�B� P�XR��]i�G��!U�T�q���!E=�H��L�'���^���"�%�1
9S>�ޗ~�����o�Ak��b#�C&)���~��\�y���1�L�ӧ��������ޚ�"��ь赮����*A�JۼE:����\!��R�q�Ƙ����Խ[LH�Xϣ����,���I�ڤQXG��'Y�!b�P���'��9*�b��V�  ��G��7ti���o7�>�RO��BIR�ſ�ca���[�ݒ��U ���׼�ד����/�}��5!P��[���V
���?�{�Ϋ��Fd?�*��9*4:yK_����ǔz0��h�-��U�WӼ����v��
[��R���tz���i�-w󽟟�ͣ���iԚfz�����i:^�0h� ����y䑊�_�D]������ٜR)a�N�#�ֽ����-��5Ro�E�'rm��c?�I*�#=�i8�ޟ�Y;�]P����d;���l�J����~�/_N�,"�
[�Ӭ��.�sۧoS^��ҕ:~6�wX�=Ӭr-�*]tuttГO>Y��z����wJ��QjX�L�BH�(�\{)�|o���~R��f�&B�s�� ���#C�B^�Tr���n�)�����Ӫ��*�yN�����鈼Ӭ�c��)�מ�bT�>�fEM�Ye����DX���:���e��|�嗋s��SO���+9�G�H��d�M�,X@�/&P�~�૽��W>����yH�7{P1
�c���Ubt��(�}P���EԎ�Q�L�Nrlyr�Ø��Jj�R�j�[o�U�a}��'[�X�ǏO����裏RTa��<yr�Գ�w�q�l�2�#��5�,��K>�Ƭ�o��Z�!�؃�BG(�Zd��Vy�Uy�����z�9)��B�gެ����#��\0�&M�������K.��(�R�7�tS�r��c�9�f̘A�x�g���N�\�_LK3��bA�U�-��L�R(�m���,������d�y���D�ro��,~~K���#����{P��
��騅��bQ3'���є�b�@؀�C꫁�w�Y�w��=(֬;��-�r_r?A�ۢˬ)"�E��PL��Z4Nkň��C꫇���|��h>��>���(<���9�xKy�w�1g�Z�\�׫��aH�&���\q*N�cf���7Y��pU@`Sض�񝃆�y����G�3��g�)X��z:餓�ea��=z@�D�<{ 2�)3�S����؃� ��,�"Ups�o�	\�^V>�N�)`v%&��Z�j�ӘEQO;�ŵ�d����5	�K9ObV+�]i�
^k��'��(�=K=i	���ԃ����� bE��=$��b4+Őܘ�B��$2�����Ȗ�*Q�@�W�B>;�)ɍ���z��F�8�X,s���/�k��}h����NX�s[�DA�!�  / ��$dK�Qs͛��ҫ/L4�?w��9(
/�\bG;]���~U���AvԾ�{'���������e&r��y�\C�h��.���_W�D��$g'p�e*g��m�kY�-
9./��X)V�pX�y\�N8�Z��/��N?�t�u�t�B]�vu,�ɧX���{ D�=(V��K��L=�a�U)9�H��)g�%r���9f4W�_LMK���	ZtSMC�`d�F�����H���i^�c�f��]���J��+�j���������AÚ:�
���b�GP�p�)H\�y?͢W_�����X�t%m5����wTڼ�;���[n�X��{��^�zQؐ�OA��6�R�@5�);WJ��53'1i�(eW�؇3��� �|O��j�8cF��L��L��E˰?w�cJ���*�W��p��}nji�4ʙԽsOet�y��&#�T�r�x�T�u<n��)a�m�Ϥ]Q3�g�r���N++�2�4��xE����裏��  ��td�\U�U�O�<#�^�7�\�[+�(�]��*��NS˞^����ڦ�Q{y>�UBkjy\��88�5!�5�5F
��b0Ω����iV���4ˬY�VK��3�9S����}X�H����  �����{)�d�l�+&d���S.P7(���B�;�^,��Η^e6��(���W+��zo��bUW˄�N��#���u\Ǻ���e�YST��h=��|p���w���ab֬Y4o�<  bA*�l/��x�[�j�����sRV ����[��})8�n��������U�����*a�4P��n�1mt1����c9��>_��9��x�2m�4 �0�%G�9)�2�I~��e=� �A�le6���.��2W�l��ʚRIӳ�W��CD���d*��(��)�j�  �6{P�DW�������H���I�2��!����j�}���*!�!�<u��sY�O��k�}�e   
bA*5S�*��e��m�OT;H�*s���؏��"-ߞQS��}iZ%����J�9��   @. ���#���B�tJ]�b�-%9ӎ�,#���G�9.�*WKL��   � ��C^{	�߆�Z��q��P�rgL�2��2QKr���.7^�^KƱ  �@�A��,�� l�u�ez����L���V��   �R � M6���]-Qhy�� �h���6h���1���^u�8�% bA�lʉ�� @Ahֿ~>VZ���;P%,���pg��*�{C�   ��G�J=�u_�A��CO�7Ѭ�۽�-�!�    �>Y�|���3=C�A��H(��y�4.�ce��"��G|  ~���������䌝o/Std�^+y>'�>�@��$Qs>� <��c?�R�%������[Roɽ�Z(�}a  ���������8�c1͜�N �:R��h|�A�:�z,Ӭ�$�9���!��%��V�!�����ܒ�k�\L׏z7�(
<��r�ku���2O���ya%M�j0���y��%��++	��FSF�є<d��\̮3l��|����{�d���}5Zo]�J�"��Pn�w	����v�Aa�#�g\��>���f��I�]1��5�;4�K��O.��?j�[.D]��]^�7Vѵ���Ӯ�O�]��<遥���+��GɴEǊtJ�R:��
��kGͯ��.+�j�}�� ����+o[L}z�i�_t���ѡӹ�R�|5��κz>�|�`���?�eB�.���u��x,����{�t���V��W߶���O�hՇ�R����'� a@SoRz�н�4��2���� �F��c�^^��:%�л	�� ?tv�;�����
\��',�w��8��E+]~�B���Y��XM~x�cٛ��u����'��0��OZ��Pg¹���[銔�_~Z�P�燞O?� �<�΅1�bIMt�Mj1�DRK��� ��ڤ��|��?�λ;��):b�'�xه�GNS9���4��!���z
��N�޲��~����Ko��H��}��+Eε�{ޯw��?�7�	������::�_��U����ǅ�<?��J�)�9�f� >���'������S5t�xyt2z��d%@��גʇ���K/���\9MUJ��u��53s����Cmi��Z�2I�|>����4��_����%�rJ޳�"<h@�qL/�u^x}M�kq�u8}�+3��Nӟ}c�U�wd�I�_+i��z:|��.7�!������5�>&"�<��N�G1cF3��/x!��A��;�`�T�s�} �� 2]7��S��{!����1���S׳����!���c�YP�/�S��o�&�Z�?܁��H!���T�����5Q��w�i��_��4ݿo��o��T�|5�]\�-m��o��ꕪ��Kmv��> �	K�c|M=%�:���3��dJ=9s�x���%��.4�k�+_�n}���.�^H|,�&��k�������;��+�Qc���8�<�/��O�~;�����F��]t�B�z��-��o���{��ެ�j��?��i��!L������S�T%�[��y�>��qg�zb4%�i�*p~�H_����.�G3�^~&�{]��e���;&�ՠ� �9��kGS���c�!�u��+Qz�fʽf��#���/�m�',���@u����������)����ҭ��-6��}��V:���N���#�9~0�?����v����+�,4���������Fgqq�',�+V�M̐]���u8oF3Ed>��$Ӣ��6���@��W�����o�	�R�q+Z�׶!�u�����!�1e�� �i��Q3��u]vڀ��T���
����G
ik7ƺ�|�`Zw����_�9f�4����ܯ�g���!�Ɛ��4={^'�x�ϴdY�R/������Ӕ�Ө5�}����\} �eZ����K�c��'4Jh	!>IM���H�1BNRF䕏��.��/�- Q���ӟ�����[I�a��)r_gF�딈=�Nf�U�?nmm-��!���M]M���)����Ó�p�x��Z�LI�:��=�y[�Nw�s����L,[����/��y>� 3oA'�t�ϴhi�R/��|�Y?Q��`���5�H==�-2SRBRg&�T�ńܧ$>��%ust�Խ9b��%��^>��+��:8�
�ؿ�o�C�cf��{���:GĞ�}wZXsK3%:���d�'����@O�HM����D��;ST�=���:g�����9�pI�R/ᖎ�U�� �0>�d��_7;��9��Ha`�O��덨��'�q��"=C�XUϰ���f�xe*9�,��1G�e�^�RrϹ��s��/~�����c��9�:���t���O:�  *�������DC������
!J&)���q�>��z�;��fB��t	���@]V���<�"o_��ѝbV����9��:���8���kE3�    U㞻/��!1i��jO�x���SG�$�'�	�xC�����t�W�"��]p���s��(��_s�˖/��{OQ��   @�x�����Hn��������4:��t��BO���@G�M�)դd����Yh����Ya�6
?�V�	�__T�Yb   ��r¸c豧������	�љVw���G&�R�x)�c#� !/��q�Vso#�l����(�c���z�!z�>l�=    �ʊ����1�ӝw�Mn���5͕Oo�:x�([gG�1���uMe�t�G�y]]��w�#���D'M�8��|gIb   ���rȁ�>��w,:�(���R㾦�ez�4-c-����蠏>�����*�a�̒#�    �᱇��ÆѦ�oA��.]�rH��PL��\c+V,���Υi~Hm��yb   �����7 � � � �F��M7ݔ�zꩂG}�i��(�HЛo�I    �} � T��ݻ��g�M={�̺���7�Ls��ɺ�u�]G믿>m���t�W�}<��?]u�Ub\�wܑ/�g�=묳h�6�{��<�=��   �� ���t�ڕ&N�H[m������b:�c��̸N}}��;v,}��"r�=z��<q���j�#Rl��֔/\>΋    �b@a��<y2m��f��2d�{�t��Gg�{ɹ�K������j�+��R�!r   T�= e���IH=��3��H�ɖ��{�<x��{��Ϛ5+��\|��t�)�P�9�s�~ȹ��_v�e"�/����#    T�= e�e{ʔ)��&���|�	�t�I�z���}��W���_9f�����iܸq4cƌ��q���{�I��׿��|��w��7��\��{ɒ%t뭷�4!��g����	    �b@`1�Rϑ�O<����}m��/�O?�D��r��ߟn��v�u�]snw��{�'����[�����n��F�g��J
W    P~ � ��>}�X�y��R/��A$$��/�̸^gg'���޽{���/Fߩ���:���۴��;���    T�= e��q��͛G�rH�uX������_.:��t�j�aw   �*@��a����O��ѣ���.��R�6m-_��     � � N���oKÇ��t��.��     � ����V��뮻D*̘1c��_�:    �{ B�����O�gX�����Cl    @��^{-m��v4h� :t(�q�4~�x   @���P%v�m7�x�s����F�&M�ϕ+W��5��cǎ��_~���}   @���Pxv�	&P<Ϲ.���{�7ޠ�^z�v�}w�o����ۏZZZ    �b@�������>e�?G��j+1Qְa��SN	    ��= U����L�X��{ٲe"���k�����?���xF[    ��= !��y�;Ｓ��������墳��    > � �ί��/I={���#G�	'�@��z+    |@�1,��n�I�i�{���k�    ������c�ў{�I��կ���������    �b@��u�.��Bz�g�k׮Էo_�i��    �b@��a����k����Z�u_*�ΝK'N���>��I�~�h���   ����̰L��P�>����9e�%�G�)%���%g��6�r�c��}��4d�   @��P�O�N[n��x̳�r��u�]W����=��ҥ�;��<�LG������W�cJ&�t���O<Q�� �[x�K�����	    �b@�ꪫh���t�'R<�=�P1����U�VQ"��^�z��MMM�c���?O�]vYɎ�S�&O�,f��äI����3�:\!8p�cٌ3�3΀��'�y��i�Ɲݹ�[�n�5�����M<���<�^��  @��pt���n��?�X��*ŗg�>|x��9u�ꫯ�'�|���v�]w�.���+~���y����  p²>b�1��gL޸b��ؘ��88�b�
0��4��͛G��=͜9ST   �b@y���i̘1"z����L��l�N�J�_=�������O����y�<{�I'	���Y�t)��Y�fф	0N> 
�9�h���m�6�5�X���p�"��[���z륽>�|�R����W_}E�~���� �	��2�l�2��KĭTp�<紳�O\�iA�����1�C ����_��V[���<�l54h��m��v�9޿�����č+� �� ��F)T�%��P8��7����bԩR�hUJ8��+|�;N�y�7���_}c  ��   �N��(�{�!$Yv�/�A���p'�R�O{�!����ٳ��_��^z��,YB ��b   ���Z��o?���~G�{�.x?ܩ�����q��+w�厰<��2��q� ��pK�s~��;t�PZs�5�q�w�=���裏���{��~�i�6m j�=   ����_�<�@��o�wԼ������k���/�o���p��B��=���[&�w�Nk����P�w7�xc0`�����=<c��5�'��T�\C� ��   � �d��_�򗾷a���g�s*��ŏyX�J��;\���6���ܩ�o[l��5>~6�Yg:���E��|P��@�.{   �ŨQ���o���g���f�#*C[�adK	�<��s��}�o w��~��E�?\)�a{9����W^yE� , �   �	竳��瞾F����^xAt8]�h�
<*���%��~����7�<k�����Kp M�8QTf  �b   ����Gyd��5O$�i6O<��\Z�k�|ni��;O�ǒ�������7�,��Y�k�R@���  �4�G~�Yg���`~�������N<���w�I<��h������3�ϩ<<o�-\� T�=  �H£�q�"o�g�;�r��n1��������C^r���C�~��y�ˑ}ο�e�]�k����� �  9�N\p�=:�z�vʔ)b��(­O=����s�����8�Ϻ{�]w��W_}�  �b   R���t�i�Qccc�uf̘A�&M��>�� �ɲz�!�r1n�8�7��d��{�0�7�t����ٺk׮���-;|�1jp��  �,$'������l�+Y�Hb;�B !d���W(�@��J��e�_ii�
eZZhٳl(6!���'�����s�+_]]IW�����Oؾ�eY������\t����O<�6e�c���*����>�%��N��;�#Ԛ�[n�E�K�;6LF��.8���� ���m8���ذ�2.�6m��7]8�K{""�x�?��jép���{��_���Rd˖-S�$����j��>(w�q�|��B�����ԩS�[���aЌKQQ��]���,X�~��6����u�DD��v�yg�ӟ��B��6>��㜥��7���ꫯ�7�����5Ci�m�ݦ6�z��'���Sؘ젃Ra�M=\�=�X�=	�����[�裏�~�{""�X�����~v�'�Dn��vY�f�P׬X�B.��B���T�L3��!g�u����Omj��S�d�������'a����.'�t�꤄���[o��͛�������2꼱K�UM0|��'r�]w��7P_�2��K����999!�����Zfb ��~�Y(�A����1cl~6�y��}�v�3��/X4�~�0hƙ��cA:�=��<��Ng���0�8����SO�E��6��}��]�`ODD�c�����ʲs��#�<�������0{;q�D��c��/��Bͼw�;�#�W�V��f�<�@U���(X�L�p��N9���$,�F�;:@��3����ڈ�c�ŨQ�T?.h�ZXXhy[���z\P��NL~��x<!{쉈(�`f���/W!�3��19q]m���3�O?��� �w�ʕ+UY���G;vl��(��FV7�t����
�f�O8��� ʞ"���9s�����{�kZab���+����X\���{�M��uV�`��o���>[�w�}�gzl`�'"�����p�3�X����X�� �fRsssUY��=o��p���=`V�EY��F@l��Qn�p�M���l9�Z�� J'����c�=&���TWWw�{����_���r��7ˌ3B���-X�yϰ�}x�Q���i0�����O�g�;�˳�>���̙3�����!�<x�:�v��'�.K���
�����2�K&�B=��z�v����Ԍu"����
��zv���@c���j�W�c��կT�{�W�ە�pv%7x�Q�m��,�e;��k����
5P
�g^x�Un���g8c��8&1@����L���������<R({""J{(���UM=f'���:�%�A5����賡�}�����FB� ���ѣG>g�ѵ��0V��ŢZ��w�q!������|�p�CW�g��l���s��fė/_.� �3�~�����{$��!�C�δi��٧�^{�lM쉈(���f~�:o ��4~�g�z�v�HP�����ΆZ�E��\rI �����S���?�|��R!@�B�����w�E(�E�^(��F��0�=�Ͻ=�4�}�?�,�~��G�z��o��F]�������]�3L�^z���~j�
nvՉ������~��U�z��c�>���]AVl���P��hݺ�:u�*��:��E9���]QRR����ֵk�Z����7�Pl�<���u�>0��a��2�X�)`=챎�裏���3�T�X��}���U��4�������Z2Z_b�^�xݙc.JxP��3Q�`ODDi
GQ*b��e��暄����f��8��1fQ��C��;U�Q�2&��	&�{ｧ�%� b�p�=��Pz�!�]�Ǉ�׆��9��3�'�xb�u���j����ٳg�����^K����J��N��4������f�ƍr�"���o����w�!��Z�z�駫Ё^�f,�m��T���)��/��6�BhB�!Ύ`�"B>:��R�Ѕ���)S�]�����E]�7zo��ڃ�E�٪U�Ծ ��r�(����^��n���t��(���ћ�H`�'"���.+ư�Cp���[�~�dC/xԖc�������^$�u�V�Xpfe�u5�v�E�瞫7��Q��a��
�5��̒�<B:�!������녋";vdEY��y�-�kQO��p�8%�0[\}���.qi�;���v�d9��r�#�!>�W|�>񹵋�'�&�x��S����]׮����ŋ���SevtP�uX�}�}�����)_Kg�DD�VrP�mm�Ri�~X������#�[o���ǀ��YN}-�8J7����Q
�7�y���L*s��=�Q�ol�	S�NU���Eco�V�L�K͚��T��S񂐞]�+9��$�,O���h�|^���)SvIp�&b�5�Ҷ�Eڶ�H{Uk\�>֣`p��$�(�,O��x؃�[UTTHo�`ODDi�81�E�f�����JP�� ��H�Ah[8x�>r�����|�}������Y�&�m��MR�qc`�m$��׃}ii��p�G,�Ca �r�Y������_�B?v��GP��3,�6�8K���T8�����A�3��������#y#$wH�������w���.�Q���}U�o��,-U��y��E0h�N�X��1}c7��g�p�g��;қ0�Q�@����Gk?��T����o��ٰ#dҔ)2q�d�e���z����TWU���_�x�,��{Y�lYH`�&E|���X���s�e��\�����<�L`a.j�q������,2�̿����Wo���}���k����Iw[;f��`׾�;��8s:�6����?�G�}8�S�z��rHް|u�4��e�6P]]/�֮�]�4���5��%��bm��%k}20�QZ@9˩��r!��v�&�=��Î<R��1CJ-��tf�q�4u���T�����#-h��g�N)��Į�z�t��Y����CKE�qt�A:t�u�Q��h0P@��I�&�|0�CyUo1l�0�Z6�zl��윝	'�([
w������
�� ��A�5;���v����h���I��~Ҵ�A�Vԩ��X�~�
���M�PƄ5
(��-���R��b�1������D�XoI�%8�V3�h#�z�jIU%��r��Ǫ@?D�=d��w_uA`G�O�K-R�Sa7R���?���[�N4��ۇ�p��/�Ÿ��{�1@��ͥ'�!���>R�_2B(�0ۋ�G`��Xʦ���]R�g���B���7���u�/�dW��^:����!?h6o��b�΅�gT�4�m��e��m�}į��ju��xVkr0XB;�Llj�`O�"�YNu갼|sh�#E������
ˍ�(��>|�ر!��ϟ��lS�@����SN����@=z�a���3�eْ%���ϫ�,.�7Ϛ<y���GA,X���	q���X�+t�y��U��#$��%;�b����0xB(���	N��](����C��Rj�Ο5�'�|�Fz98�7p�1��j��#�B���c���9���ߥH��(���5Ҵ�swd��(��nP�o��=����{��曻�\�{�����C��-[�c�P��]�ѢԆh􍞌Pr�� �VW߿�Xξ�5Cߕ���2~��E��V��?�y��x����[������983b�f�uؔ�;�	��.��O�q�pf!�݄���9ǂO#�c@痮Qt��;�D\E�3���y��}_g����p�a��wS������E�>�
���n�8�hJ��ȗ�o�b.�ihhP�������j�:1e����zĐ!C�L@���L߸$/7W,ӂ�v�{��:z��3��16�h :�${*#��z�rᥗJQ7f�{ڮ��.o�����{o�wBw���ҏ���?j�3RG�ģ-%���g���{,��}�?��c�2�i�����a18��t�te-���xP�>Co�x��Yo�����r�&����Yz��;�{��3x&?�}�|�#�r�I�ქ��*i���sPYY�ں"�K�0p]�h�|�����3ܯ�k�M\��`��L�r�e�rG�Px���C���n���n�X�i���W_}URŨ�w�kn�Q�X���Q�G˚-[d�֭2հ,ʆp�%6�x���R���p~��>�z��SO=%[���.L��P�o���ź��6�`�^��4B�8f�c�`ɑ�T��yC�g����?�{��x��s��ƙ���o��olN���Tpi�\wܗ�_����ǣ6��z:2��}�~�L~�B^}����{�� �.k���U�څA?��0@�_��Z������N9�D)���@�YUU͙{z�O�N(�=��5�8�aO��kԯ_z�U���S��Y|��we�q�dԨQ��Pߎ�\ ��(�[\�P2�I�x�@y�w[�`�)b�X+��l:������s�����%���v���7�x�Ǧ@�z��C}V�K��lq�qZaF����i� ���$�Y�mn�Mn��s�3�S����q�_��{C�=�,Dv����B|m��/_�v8ƢZւ��&>3�|���(���,g�x��z����6~�xUk�Yd�NO6�˯�F���~��8��	A�����B�S@��lUo��1x�Y�r����kr�	'|���PW��>/��13�M��0�M�0�	0+o^,��㏫�@����T���Y������z ��PC&��9����唸т�3ץ.�7WrOs�x����v����:�s˙{������Ϸ��vamւa�=�bZl����[2�}/�3��Hu���l5Q�d.Q �^�EL6����;dwm���mmRW[�zl#�����w�3�}������Y�E�k�Сҿ�D.��r)����Ps_�3C��fb�mOl ���0x3.΅��>Z����/��1c��!��{�E΀\�7�L�C������{�}vq��s%�(֕���wC�x��T�NǕ�Y|�l���7��� ���Z��O��p�}���>�{b�T�m^S�}/��fx��<�iӦ	�.�}s�ԩ!��}�ݸ�rw�X�v�]2b��.}>&Wj���B���d�;&3|>C}�>6�{�@�Z�/\ gJ�ʤL���ځ������ܣ-��+6�B�u@���eɒ%=>I��1p0�Y
�x@�ʟ���{�E,�ivq���^�%9	�����Yv��<Jo���٥}�U��@g��rD
��]�.��V�[��4'B��wI񁃤ꓭ�m����8�{�m��C=��Ǡ?�SM��Z��`ODD)'���%N�aZ����{��k,�֭�U�k{�BD���5V���p�6`ئ}��~��N��1vF�c���kU z��7T�2.��x�b5�m�a���ƺ�4U`a��kFb�5��&��g齡���d�H���8������kZ���@��h�O��(՟V���^�_�f�ڧ��3��XC��N������R
B�r����Kj	���+�P���i�F�R^2#��z�i�F��=����U�q�E�u�L?�up{<��g�?�`?r�(���m�����+���E>О�dy��'C�=f��;�8y�g$�`A0v�5���F�r�i�v�A��u��z��|��F����Ajal���Y8��ijO]�:�`'ܻ�fK�����Β�(01p�a�-��կ~%s��͘V��DD�RN8ᄐ�k�_~Y����y�4lxcJn֮^�gA���;4�W̎cA���^��'�Z#��Xt(���W����}o��I~X�T�ጃ�uK���^�f����kI�ڣ�;!أ]-0N#���`�37�,�L{���.8�]�ۍ���x��@��Bվ2�aЁ:|Ou�z�v½�W�<{���|���w�8�>�h���#�H&`��^��{���Vl���G$/7/hC��̲��s#Q�C�9sf�q�Q߰a�$B�� ��.���D6�[��n�\n��q�Y�os��$[{��{\ol`�\3c=��_;�?Hhӂ�[� �TUV������#���=�M��"�_y��^�J���_�[��`�z����O-�M�hϻy�JC���(أ�
����ު�+�����`�U������0�ʜ.�_�G�5-�=���Za�(���i^�h�k|�R�A�qS��?^mʖ	`2�S��Y8,2�c[�6[=o���}�R_I���Ƕ��!�_{�5I��/�@��sO۷���+���s�L}a,B{���FoY�0������i8c�0܇Q ��i�����}��*ط��u|���+e���K��,���]$����S<}��g��\��^���Ѫ��3Ă��{�����#c�v���,c��՜2��W)éz���ݣ��RY�_vf5��;�D�k��x����XD�A�~f�q쓀үt�`ODD)a�����{I�}�?�'�j�#i��Wu��$�����9�𞓛��W��1{��h��>�a�_�{��G�{�_�o���s���ذ�5�(ͱc�a�,�?�AtCB�q#��c�;��:,b>蠃�����K��h��N�wi�����E��	.�q�ϕ��ػ"����*��XT��Q�0��k1�1��`0�o�R5gk�s:k�ե�� J �31���=��h�.fo��vR��(+�kn��vM:��W._�@ָ0V�X��5�X0�@��aW��׍�x�xfm1��������~�@��h_]e�����#m}�r�,�?_���%������n2�]���!�cJ����������cx��,G�3��ު�^�ԧs�7� %�1�����%9XL�gL�4���-	gK�i��s���X���t�`ODD)!�j���ٳ��x~u�j#*;P�n���z�УG�
��[������f�1���|���c��-�?���?m���6�k�ڵ���Ѷ���.�H���+�L�,����U�����;�������|����+��b��)�4WՑ���HP��;�]�Y~Zb�,G��pJ`wZ���q��uS�xl��ǚ�y|���cؔ���(ۈ����R�Й-\�Pmޓh{�L�h�i�7˗-
�z8׃�
�}�j���=p�^��ݳ�E��:�������0�P��B����rUnM~A��{�r���$�6gΜ�`���P{��;��uml_�͒^}�U[��.8�W,Jp�3��mnY�wNY���+�U-�޾c`�쒃�?EK�f�v[w���(��gJKKUC�o��F��=%�p��c�������M;���������O�����g��{�-B��s���X]���֫��ה��e8C���3�3����C�<R��]U��H�d���v�����nPNs���>����Zy#�U��9[/�%8��ˢO}ajl<��R�����\�c�;��:��^}�?�(˴A��ߞ#��7�=Q7`&�X�˟~�i��q'�hkQ)�1:̘w����f�f�1S�矵Wa�����e6]h��ru|=U��FЅ�*�oW3�vZa�{�Er��'t�ʆ������o���v�Iƌt�ni~n�c��g��=�ko�K��37K2�?_��nu�}������}��+{���y����:�%�T<0�QҡÉ�����W��??�$[��n���6|�(���7vz���{�Pֿ�����ܣ�nз��"P�zN��VN�@cw��Z��ƌ+{k?�ys�J"a�Ps�ǂk<�v;�$�O~򓠏Q2�M����/�������Y�a�,~���k�_�����y:��@��i�>�]�#��mQ�g/���� ��"ܣS:b�'"��B�4�NC2N��<�h[��Q������j����F@�,�Koe�
����ew�}�Ytc��3f��� �--���B�Rͬ3�Hx��zM�y�4iRʕO�96���ݳ�uV����ݠ������I3^�Nm��mh���ֵ���k_��&�"oα�q-��0�u��#,7��7o^B��ɳfٺ��ի�,�,��s�����P�{c���ii�����xx�x<�`� s$��/'O�EH�lݺUu39rd��=��3���;��������>�ˢ}��l��(����3�wE9|��fwǂ���ڣ|�����|��zJճ@���W��	&�C}�+�8�<8��P�^�_���z�}�
��֖z��+J<�l�YGz����Я�ڱC�ku�1	��NI�`o�J��S�}�q�Fٴi����3����j��短�&d��7���OC[���VXH�7<_�V�G��o��6ha6�"��x�a�'"���
e?Xt��i�yd�� L���U�z��ꍡ;�5�:��^=~<>�c��]i����:�H�?� y�����5��{lбq�Ʃ�ܸ�9�Pd��� H�a��N8���?[���gNf/�Ǒ�%�fG�	��]��{���ߜ�'�M�2�����(V�En�t�҄>t��ӷ���J�!��B���^�z�s盠�C%�,'��8v���k�m7Qo�҂=��d���=������#��d��ǁҗ�+WJ*������{[��38O9�]f��g�����z�%9���8��hhQ�䮋>�����v�N�DD�4�Ç9�ٳD������6,���+��Y�aUO��2cliid�z�\��x�
���O��Z�C?<��u�555!�2R)؏;V
��E	�����������oy�����j��T�|�;b9�ʳ��:��ǻ��644H:�ݯ
""J*��v�B��Y�&��c�EW3��KN�P��_ �����<n�>j����=a���&������8Q���DY�v�*�0=z��
��_�^���m}n�@�L���o�
{G{ˈ�z�v��cql�ߣ��<iZ��	(����F���	��������f(ٱ#z��x�h
�V�o�ho	���߳>P��>����2;�6��V��>��8���������t��=~��D�C��~�]v�T1´��d�u�t���;S�%9ǰ-u��{�<�'\�}΀\�nA�� �30�`����`O�FP�[YYi�؍��݊�
Y�pQ̏���E�z�aÆ��ll"��x��]_��[a�X
�Ne�;��3�N��7�w�M��1ܛ7�
G��˿;m��c�f��c�g�ɓ�׭[r�굔,�=h�i���7�Oc���.�8\�sѬ�3[�_�u���r�ϖ���g��s2�t�`O�Z��m?��
�
-k��2ِ!CB����a�i���[Ԝ��o�Z4믭w���e8� ��;�:��W����5z������͛C���������d3B����=����J��Yy�n�]�����楞]�k+؛N�Z:ૃ���f�E��m۶%�1�5*�m�kk��}�]�2��	ǿ�4�>E�},�u�u����Q;�$���fx��l�"Ʉ=�Sٝ@�*�e�u��Yy,�1B���y*��K�`���m�DD�49��`6�Ƭ\�C*�Km��e8jWY\aQl��8���c0`l����%E���0oެ�㉾sgQ߾ҷ_?�3�z�;7��P��=f��;�?�3V�lPt��N���#��NV���k���)�v�e�'"��)..9�腳�m{�����S���ްH6����};�>��6�~|�nC�N$X��,A�����Jt��6�H6�k�g;g9���OVh�=�&�� Kj��D\@ku&Ċy ���}Ity`w0�QR`A�y�У<Q���,������b��i�ݎT~c숓������|��U���g�u��`?t�pYf�yTO�Y�T�}��	���0(��V�D{G��:ўt��kiPzfl�۷o_{""�h���,��^z�+9f\-��E-.�I��{��b<���z���(�j-�$�1X1{�Nő����n��6����tF��3m�_��_G�0X��=%E�`__}3�x�3�0+z�5֢�f��;���Mm��HV@�n��RPP���{;%6�u&xZ:W[��;���cc5Č��Ύԩ����:���e��1q��9}&�����}��ײ�bW�:c�=�q���BCf���K魬�p ��#�K��0j5��s�x��'C��og��`�j��hm9���8N�����}i�(���Eny�P�o���gX���Je��ԩSd��]�~�۷�`��3a��}���v��/���m�Aa�p����}�D� �;ci����AZz0���u6�}~�g�����d�r)g����b��	��T,�"��DD�+Y��D�փ���$�ȑ�>*�_,�e<X�VR!�����}Ecc�D�a��5��I�뺻쉈()��&������p�݃>U���얜ċU�[*��σ�3>w�׾���1�[��D|~�k$=��]�DD�Ve7��gm�f���2S�����f�]�e�<X�����n#�{3�u�e6�:[ϯ��R��k*�DD��P#m'���B����0������Ot��z�X-�M4s��cc�<�etQ�黩v>�>��M��YO��]�p¿R��؛ϰ$�KW<0�QR����H���	��h�ٹyy�b
lƚ{��La���6�ıl"��}WKq�m��y�n9���~]�z����Ot,����k>Ò�}5������"\};j\5K�D��M����o�g�!��8��lڰA�\�����������M@�;��{$��{^���6��O{N;ą�ip������?��'""��j�P@J�S�h�!���:�
z���{�(E��;/H���%����r,�k*�***�>����Y?O���W�i����?ԛ�$��G���L<�W;��1�*n߾]�	_������0��Woٔ�Y"JM:���nGڞ�i�ƨ�)��Di�A�8�c�ۦ�,�vh᧵�Uɸ;�.�&�l٢�q!����e���Q?�S���UՌ4ڪ��۪��$��g��MP��a~����:ی�I�6Xe�K�U�˵_�����ܱM�����Њ���8���c�����_@BN�Jp|"Qgo,/;���<��f�:I��	u�b�f5jT���`�npK.�	���x�Oڣ�����F�L�vf��7���{""J�;v��!C�$�1,Z���́�naQ���g��E�^��h�a6߸`VT���N�_���ݙ�gu�j��e0ɂ]�����i��<�h�:�v���Lm��V��P�b1���h��w6�������n�*�M��J�c@X_�n]�:�ee�`��lt`iokS�����d�8{o,��[gZ��t7�w�~̏�?�{r�[}F�(��~������zJ�@h����h�8��Y_��j|�nq�2�I{�2O�[-��c�ȑA3�� ��f�������G��Ⱥ5k�쾺h����z��jA8++˲$�%���8c��v��F�d�A}��#M��3=&L��x�����Ź%9�8�}�ξ�]��� 'z�O����Cs�߰!���UADDIc5�jwv3����+��I'E�;�}�*�������B;;�8\�OF�7�N�������.��^#V��dY�pa��%%%*4�_�>��mo�������G-��x�Ӭ���wL��V���������M�<9��SW�Z%������f͚5!ǆ�v���',^�@�WTH���o7d�0��J{-��ǥ��v�}�tŪf?Ҍm�����
�����z�	d����gϖDmqve]��D�m�65h5�M�2�V�o-o�����?z�v�6�#qc�^{����j(�	�+��ߺ�޿#�F�-J��bՋ_DD�lV�ar��v�~�!a�A��?��g͊x;�"�9�i�:t��6- ���Ņ���V���\c�P��?kuv*ԣ��_f�g�8�g/0(J4�`o�ZJ�����O��������z��k�nU]\��������@��.N�xZ{o��u��G�)���-�k�w6	/�Ix]�C/}EQ*��B���RZZt|�]wMh��<G�0b�(���Q�#�?G��K��c�SG�Z{0����U�?�����؝�����	/���ʼ��Z�G04{<�v����R�G��r���`/����.�>ѻeo���k�_����7���s}��	^/�DD�T�c5{,6|��7�86�['�ϗ�S�F��,<X�mݪ�q;f�`ߞ�+Y�BZgd�p!>��>\���h��Oaa��D����3�q�ƅ:��LB/�H���3�1�M��&)߿3�:o��8(�o��^��&��E����`��m����<0�w�W�^-������j�ҥ2mڴ�c�����F�0|�H���T�݃��.�����ŦXH+�Zw�����̽��ܦ�;A���"ݗ�u�@�Jp���=[�-	�%��sϐchK��?�g�V�X!��[�ؑGi+أEc��&��o1k����w{���.Y�'����;g�#��4��W5�v��b4w�ܴ�qV�`ODDI�dɒ�cXt8`� ��U"a�~��x�GX ��3FV._��ꊓ�%������A���{c�7�z���z��	Ww�:�x:f?q���ΆT��_z�yI�`o�J�k�c�?������0�ay]G��f�;��w}�8�\���-r<>�AW�D}��v����B�]�q�hv���=%�r-����Zq���w�}7��g��[�3���Jr0�ݦ�{��6]����[�Y��t�	'���ǿX��o�Yh�>�3Gʓ�yO^^��ٜŋK*�����/����������~���MZ�5K�>�����:Kr�c������G2���M��T��k�ks��̙3�>�dB�.�{""J���VU�3iҤ����_R���_-_���7cF��b!mSc���׫0ݦ�z�}�;�#���>\Y�~]O2���m-�P�E�vJp���䱇�d�:u���Tb(��od��t�QG�
���C]G�cI���������OS�d�gnIJp|��%8��o\Ug�>�z7���g��e8�`ODDI�����~���R%,z�H"��d�"1�	���q�T�NkK����CA�d�/��Vj�%:=��V���6@�h���ٌ
�}�I��2��g��c�_���
�8�`��	�u����^�*-%oDg���&fN�-�grv��{P���$��$Ӡ����W�utͱ�ft?�t�`ODDI7o�<������,�����ۄ?�
-(���srƹ�F�-��nZ��a�R�z����:��Ӽ�6]q�^�hk����'?_����A�7_}U��"���aP�ʾ��K������������/)��v��ϯ_\#9���Ю����m���P�||�iWI�8���yI��gS�FQ�Jp<ni\io�^�9���ڵk%�1�Q�a����ٳC9$)��8t�i�d����6G����C�k� �*��P�|}���͝q����!3�������\[����㎤�ƉE�XPm�&����/�,�~��>����O4�}n��V�&w���-�rv}Ύf9��n�l-�c���}?���.8G�P�����1}�t3fLб��|�c�'"��C���O�SN	:�S���_;ZH&읷�*>����������U˗��{ii�(��ܫ۠LG�G�b[s��x����>��,=~~A�������W��d9��B�UUU���Y�7�xCN=�T)**R�g>k�,�뮻l}>��Q �b���8s/3��CgG�o��b����>|��֖Q�lhT���eڌ%]_}���;{���c�����,,�̶���KN��?�D��*�#����_$�1�$�;�[��G[a��k�~�M���\��-��3!3�Z���v�]s�B���S�L����b�b����s�g���K�`��Ar��?N����������q��cGq�<��3�y�樟��[��)=l�8r�ڦ�{Gg�=���,����O;���k�z;%8u���	�����=�쳒΋fu�ԫa6;�,]��wDS\\,�w�c��_�ڵ�D=	m/�nݪz���g?KZ��o��J���ee� `1B

eݚ5�l��?+��o�҂*�*µ��=���#o����o�t}�.��f��u�5��R,����W��w�-Ʉ����r��t��+��I'��*�W^y��p��>�V�~W)���uWs��M�T�H�}:��cӭ����-ԋ��k���;p�%���
��L�`ODD)a���ޓ��:+�8:���>��O�~�1����N��9�s?a�$��]d���{�l���(�Qi�V��q���`�N9��y�s}����ӻ
�^$�C���j�-=��c�	9�0��SY���S%9��vZ�^�p�|����uK�j�X���4�b�^��pL���fq�M�R��E�jۡ^S��Z���gG�t��'�LJ�����?e""�5�y�U�`,{������G%���ߤ��D8�`۟��>j�e����<���I�{�[�v=�=f��~`��-��q�^zC_z=�#ܣ���/+���%��ħ��V~{��RUY)Ʉ6y���o��V����7�C=4h��e�]&�}����h�aI�d�$ϼ+���Kuc�!��:Za�ڼZ��G
V��m�[|nKK�AFy���k�y]�����	�C��
�{
k��&K��1"���f"D�\��%6�2:��T�
��'`���?�I�����b�|��vS��[7o���UڇP���`6#Ԩ�w�BZ}�9��a^���Ko0�Y��.z@�G�ߔ��e�N>�����t�7���?��O��[�j�>fy�{w�����U���9�,���s�g�}mnqWy�U���Rh����阥��l���6,���kaeܛ����?�����O�RNAQ���'�VPX$DD�\�챈;v�������&�B�%W^)?��B��e�]Ռ}uU��TW��
f�s��=B���7�ԋ�9z���P�0����.��mݲEn��:��7ٰfɼ3(|��gR��3	]�u�o|�c���,v;�`1m��;������o�Y��zi�a�^���u-Lg!໒W{�k����c1w,��к�I��W����>��}^}�U[��{""J)=�ׯ�Q�FGm,�/��G]��������i��ޥq�ݔ�.�5�~KS��i����gg�	�(�Qe<Z���|n^��c#Y�|��r��{K�V-9_z�%Ig�����k������7߬6i���{۽R�Y���^&9L��,f��=[�GX�ZӪ:�8�h?;q�\}��������,=��7IͼJ���a��v�+��"�Z�>��S�i쉈(�`��\s�5A��-�'?��
�Ɇǈ��V���n�!П�+������ż(�=�{b��9�/�s���_����8��"�-R;�����r�A�q�岲2�馛��ni�
��o����\c�=�g��9��ٞ�֎uyNq�z��=zҷy��ڹ�#��5����R��:��U(����~����}�ݧJ�2�=��O�}��RZZt���OW�s��a���_|!�_p�ܨ;;��.��D��N�h���9s$����P{����?��L��c	2cƌ�1�W�FV/����;�rr�J)l�H�h��U�׻Ψ|Am�x��;jr��{�訷���:��襏Ű�v��ZQv!�#�c�pӪ��
Z�b���l�ۓ쉈(�`�7,����˃�c������0�
lbuï-'kA�풓�>��͛;W��_U[�T��%�9�a����c��w�}���_����w�y�a����/�ߗ�'�����M�N.т�Eb6|�y��������y���_���腯8�����:ڬ�<�����y�c�����.;���Eb�}�6�g{���K�b�'"�����^"��y�jF?U��g�{�I�3{�\|���i���W�	-P~�=�Tt�EY����`�����.��sO`'`�E��u�]g{1��b��m�o���m}#=T��g�}˳յ(���{�G�o���&4��ka^׶�E�����c�����/�8�ֲ�v�m)sƯ'0�QJ��g�yF������(�s�Qm�R:�����T���@v7NR	��k/�$o��r��қ��r��^�7�V��k0`9����0�A ���-�֭������R��V)�O���#\ͼ����s[���0�d:�� ���^i��V��K�q{ｷ\��A�a`@��?�Y�n��쉈(eaêO<1�FV�+VH*�f�\u�C�'͚%�M����SSS#o�������^0��>�^b^K�P���C2���?���u��۷�
�x>b�u�0�I��M(�	�w��i��^ߝ0�������Ե�W�ﾻ��P{B����u�F��_�������-�����ZA�5�_��㘉C�N�'��e$K/V��������#�>Zv�I8�1��o��?�ϴ�-�:�4�e�]B�Ϟ=;�;�D���@����l:���7ܠ��c�ipK���7�@
v�+���b[�w�m�lUN����&M���t`�e#,FN�u9=����Z�q��%�����BBc�=z�����g%�mX�N��.�?��L�{oU�3i��㩮�V-X ���|��'R_W'�b���j��YSS�<�裒�?��'�N�8���<����7���K�v�[66J˦F��G
v�+�Ź�*�W֩�����X�`^����ʽ�=��|P&O���AZ��㏒޾��u���G�#ô`;|�H2t��ͦ� v�j�X/\(�׮U_#�`��7�h�`��������,���{�c�x�e9蠃��vb��(s��9y#$oX�8�<5�����MҼ�Aګ�&��c�Um-�5��Jw�uWF-�������Rj�����K/:�:�����S%9�PjbV]U%����r�� �r,�f��1�Ʒ47K�v��|�.~�
��[����_]ztn��l��e�=��FK蠃A����n}���-2s���>#
${@n��|��۷�H�Fi�֢Ztv~W����N���?�;�#�K�z�=���^{M;�0g�4����\rIJv��
�+���V��`�ĉ��_�2�8f���"�@tW]]�\{�r�-��4C�T�ɹꪫT���c�>�W����s�Kr$�,O�|W�q�8��<�nq׶������i���yqq�*O2�-�0�ڜ���a��^#������mq��ή����+=rs�rCv�$�N���,�#�<R�s�qǩ�]�JK����o)� ��Y�v��V8#��A��c�	�����w�Yn��ָ��a�M��9Y�U�%��lq�f�#ǩf��δ.�jKٱìW��[o�G<���nhW�{ʔ)ST�/))	�e�oDo�`O���L��م�B!��6oެ�֡T�h͚5�j�*�ԇ2
�Hw]ա���/�(����{�jW��_�"hr	��1+�]Tq6gz����<��mSʑ�>�l9��C&�0���vh�ۛ1�QZy��e�}���:(�8Ϊaq!�rRiWZ�v�嗫23����Lo,����tZ�l�j{���:���z?ꨣT��jלt��7x��h�588{��-Q�b�'"���N�F�R�!C��s��o͠ť���Q>e��|ܾ}�P0��^p��<����Zb��#�ha�?S�w�޸�����?W����쉈(��9v������v��馛�g}S6`���-�{��'��α���ꫯV�`082�M@iʑG)�����+�<���k�	�sa�
��k�]�0�y�7�:1�QZZ�n�����oRo�2�ڣ>�7��Nu����V�e�	Y:l6�l����P4@�vs�(��s�9�$�͟�y����t�R�Ї����߫3�ׯ
�`ODDi���=�ܐ��I�z��Mɇ>�8˂�̰��u��Y�r�*Q�����|AAA��8�u�'�O�S��}�ݔ]X���[�z�ja���x衇�O>��`ODDi�g�����P`v�	'�n?�0g�5᨝7�M>boQl0z��W� ��a���t���.8�5{�lU��
���9R�q���bu�FiJ��:�������:k�?m  �IDAT�����;�"#P����p��^r�m���i��EX�N�"����J��{�9��*�6s�����?_��?�*kY�|y���4Cḯ	ԦR(�;vl��c�[o��Z�rA�=�DD���m<Z]"�X�Dy�Ǫp����l G]���HȪ����Q�o�,2��K�<��2k�,�9s��s��?y�du̂#�/\�Pm
�q�Fٺuk����C��#F��ѣզR(ǲz<fX�E�/��RFu�I{""����BZ���c�=B���~��c ���B�Δ`v�j渥�E�ߠN����s�=���O��G�^�Æ{{z�M����*�#\c ���A .����H�����RXX�6C�Gy\�Z�p�����W;H�}e�0�Q�@��,0bN�4)�z�棛f��l�".�K.��R9���-�G D�_�x�PϪ��Pu鸠�3��~����/��bf�;��$����*̯����`ODD��7�x�������\���v�w�y�|��B����&V�P�YX�l�Ch���.XH������[Y�U�)(�������_�d	׾��=e,�C�D�D�<3�D�ꩧTW��C�<�(Ű��7X(˚��B�6�7C�{��B��y��n�������B'*�5@I,P��(Ţ��`ODD	���o�6�Yg�r=f)�>�l5�����tꨱ��@��5k֨P��&����N>��3uѡVu�6Agcp5�Ɵ3�X߂G�/��.ӦM�-C|b1�Q�!�Q�{�WXv�@�����9s��C�C`�sʝ0pb�KX\�r�L��^�㎳�9MUh�ED�]o�����㏪#��F8��q��7��r�e#f���y�gٟ0����#����Y�D� �����Յ���Y�b������Nm_o��D�}��Џ�a�!��3fL�۠$���:n"J{""�5�C��W_�z���	��Z�]�?���ꫯ�D-����TOt���v˖-Sk��%�=�*(y�Tw��2d����jÿ��;y��zm�1MbS����䄽�n<������7D��`��`�ٳgK�8�sT�]"�x����矯f�O8ᄰ����k/u�;w��ɳ�|tB9餓�s�]E#�s��N���������A��^{M���~�3{"�1ة�����s�ת>��L�6M]�c*f��3qfg*о򨣎�8Cx�0K�ꫯ
g鉒�����z=�8_x�r��G�N/(?	1႞�~��Zd��]t�t�}�Q]�<���;���� �M�6v"J�D�Q�Y
f�����z�1}m<VJ�G�z�-X���Z��ו���i���f���壏>Rm% ���jg^\"f��.]*=�����D)����2ʳ�>�|�(�j|����_�3�<SfΜqp��O��.؁s޼y�La?�vZ��͕I�&������_N�B)'�n���k!���`ODDd%&w�}�<��srꩧ��mЈ��q��k�ʂ�,7j���yv���<z���(ց�%KԚ�/��R��"���`ODDAyy��{ｪ�%Z>bot���qqAgرc�
��W��u����͛U�w���|<x�j�9j�(�k7.#F��]Jf����?�\��`�Q�`�'""����F�H�r�3f�1�#S�N�����<ႅ�F(�A����U�@�`:�455�۠��4�
��}�JQQ��������w�yG�{�n6�(�쉈�b���.�|�4H-<=�Cd�ر]�O��:T]���Z-��_��܆(}1�u��-.ÆS����L�0!bG�d[�~�Z܋��X��D������(P���t\�S�)S�bU�|��'3�oڴ)�����c�y��`ODDg�� ]dp��`m\��u��vR;�������xA}��cF~͚5�j�*UnCD��������aq,�˘;�`�lp�Q�`!,.�f��Ѳ�nw`4x,��"[,��BWt���D�{1�S�v���zX;p*����v2�l`̏��-^$D�{`!�ƍՅ����W�L��6q^�W͘E��w]i=��\"""��b�'""""� �DDDDD�������(0�e {""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD������(	&N�(���Bɳl�2����L�`Oa�\.qee��~��n�x<BDDԛ�x�2i�$��9��d�ܹ�)�)���U���5����'����%DDDD?�DDDDD������(���JKK�P�)++��)����z��ʖ-[l�6??_�l�9(�T.���6����n""���^y�嗅zΧ�~*������Wۺu����¢B>|�u�=Q`�'""""� �DDDDD�����z����#)��+DDDD_�ֲ��J��"����;!"""��b�'""""� �DDDD��l��v�mQo��w����d���d���os�%���`�������(�de�dȐ!QoWZZ"O���فM��<F��=Q`�'Ja�55RW['���IQQ����1�����:������W��BDD��1�����z���V�"+A��x���Y���z3{���� ����yPV&�+*���E���z+{����$;vT2���W���R�m�Q슋��W^��3�y晲nݺ����O��g����믗-[���O?-�x�D)���HE�v�>�R�0s߬���(6���r�g������n��&]tQ�P�R�C9D
��f@K�K{�������""�]yy�lذA$�W��z�.�@��fJ�DDDDd�o��9묳�����)�������l�Y�;�C�9�9�sd�ܹ�����j�����_�~A��Y���v���`ODDDDQ���ʃ>({�̚5K-Z�n�]v���{O-�E�=f�}�Y��o~#Գ쉈��(",��׿�%#G��SN9%���~r����p����M���������R��1�QXEEE��SO�p�I'�v�V*++eǎ�t:e޼yr���P��˲e˄z�=�>}�,^�X��D�z��v�i*�G3p�@y����/�K����������&N�(��~�*���;j�/��B[�0(ظq���5k�%�=`c*̴#�������n�M.���ۢ��q�0ӏc���������,�}�ᇥ��F}���&3gΔ���ۛ7�B+LlZ�%�=�է�H�9E���!""�ԃ�f���TTT%�=��˸�$oȮ�߱�/�{_��=Q`�'""""� �DDDDD�������(0�e {"""�������9��ZZZ��pH2�k�y�{"""��m�69�Y�n[RR"�p�=�
��=��~�:��͋��n�T.DDDD_��_���Qz`�'""""� �DDDDD�������(0�����"<x�P�q:���쉈��R���^�.D]�`ODDDD�쉈���2 �=Q`�'"""J�s�=W\.F�djnn�L�WQ���Q<1�e {""""��`ODDDD�쉈���2 �=Q�����'�un�[|^�e
{�4TZZ*uuu�a0����ү_?!""��Dij���q�&�2������B��ۅ��(�0���aÆʦM��cY�-x��o�.����p8���(�0��1��)#0s�a�0�G�P�C�����2�=Q��̳^�C��P�i[�1��2&L�3�<S�Ő!C������!����Z(Ԏ�J�z""�x��̴i�ԅ2�}~~�P(���BDD��쉈���2 �=Q`��e���eÆ�.Ə�M�����l`��e�y����$]<��\@DDDd�=�M`�Y����������K;�b��v7wN%""�N�D6M�>]JKK�� -]���}�>nw)).���̙3G6o�,DDDD:{""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD�������(0�e {""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD�������(0�ٴa�����z;��+.��_��wHMuM̏���Q������lz�W$U:T���+DDDD:{""""��`ODDDD�쉈���2 �=Q`�'""""� �DDDDD������.2h�������ec�V!J&��!Ç��}b����<[�mjjR{؅=��녈�({
�ϓ!#w���~��l���	Q2!�_|��q�Ϫ�*Y�n��ێ�u�پ�ٳg˧�~*DDD�0�e {""""��`ODDI7d��kz��z�ҥKcZ3Փ쉈(�n��V)++��-DD�"??_N<�Diii�T�`ODDIWXX(+V���۷Q��1c��?^�ϟ/�������*''Gub�'�tSWW'�w�=�}����ODii��ղ�>����L�:{{
���V<-u��F�'�}������g�x�b!"J7���j��뮻N���?'��0�Sxk�/C
�����6	{�����R�����(-Z�H8� �7o�̙3'��������$~�a��Ζo��V���U[[�,Y�D���j�q2�=�=%�̙3��.���*Y�p��;�y���UW]%S�L�{�')���������������C監�:J���d���RQQ!DD��_��L�6M^z�%Uj�駟&�10�Q�\~����x�%��'[�l���r!"�Dب
�~���r�5�ȯ~�+y��7U�O�|�DD�m�j���(DD$�i�&u2d��p�	�_�B�m�&_}�����S�=�������� ��.`Æ��?\�?�xq8�M&�`nܸQ�&�_�^��Ÿ����X1�� �� ��0`�Z�4y�d�7�?:�a�+�[\�z�)y�l}{""""�۱c��D2u�T��b�'""""� �DDDDD�������(0�e {""""��`ODDDD�쉈���2 �=Q`�'""""� �D6͚5K����v�Gj�jm�gaA��F:V.��j!"""�1��4x�`)--�z����Q�C��_�_J�Kb~,+W�d�'"�A�C(�|>�P�1�Q���z���5$T:�Π��a�|��	w;�)�3�ǆ���*.*��!���2!""J���v���U�>??_���%˙%�G]���_ !�4�nw�}�q�e�f���}��ʲ��4��?�c	w���Jzz��?��8���`��`Oa5VrJ���~G�""�djll�ښZqe�����YNq:��pj!��o���3�iq4�k�z�}^�jG�q�9�O���?V!R��>	��_� �۩��g|L��D\^��x����`.d��^���=�a5�п��:���%�(������q�j�g�'""�^���Y���T�mhhPA�T�ػ���*����V�a�aZ��D�����*H�Ɂ���q�&���D�9B>6��Àϑ��Vg �o�lDH��?n���:��Z���������}8��G��yPb|VgI��k��P���\���i��г��쉈���@�����ֶV�.g �a?ۥ�u�T�CE�7���y�+,����#��A_�j"�u �Z�W�>���Qn� ����>ogP|�3a��(�Τk?��Ƴ���y��Q����-����B @1@�v�+ED�"^l*͊�� ��U�+^A�"Mi
��A:*A��JH%�'����g�ϻ�ξ����ٳ���o>�ݝ�}gvϞ=����}^G��T:����'�V�^'�iqG0�k���Rss3����w���C�   P5���
�ejG�Y�e���a�g���N��22�W1�YX]�W]m�����˥n�#↚$�0H�K4������d�o���o��z@}�R�S3���}�#3���������0a�!���|"�{    T}��l��z#d^I�	C"z/So,���@ �c�i�Rp<B���@�9�٢���)�"R���H�Q�I=f>Q�Bq�j�p�C??��h�j�XD��$��Mvfv��!�iii��.5{    TRPy�FD��4,�"�FF�q����r������F!������V��z�Lw\'�W;R�Ћ��_�i-'�O|����.���Z	�#���c���=�oq'��s���J��ollL6Ub���   �*`Yc1���9@L�؈�Χ���F�V|!���5�օB������ܫ
-�Uq�U,�w��tn��R���8�S_+�?��gBVO�c��x:RWW�H��ϕ��=    ���"�b�ٖ"���Ȉ�zQ:шwԒ�j���H_>"\H��\s�L%��L�޶���;2O�J/�LJ��ׯN�+8c�+7��#?�BG�Y�y0vGGGN�R�b\y������ힷ��+� P9��������?v\ZpժU��  ㍌���Ԋ�8&�D��*��z-�D��\Sb��p�|�_=�l�����u;I���K�^�N�幊R�<9��b�zQ	(0&��{YƓ��y�������=p��"  �ħ?����K�_����O��[��[o�E �7\�p���}b������ѱ��fY�x��W��H�U�3�$����f�C��9�����8�6�6m�g}�����g,���+���(	��FĠ���	~}]]ɣ�{   �G�n��fz����o��Ҋ+�񤩩I�:[_��!!�r�%9�N��U ��E��mVT��cU�Ѫ�):n)/r�z�-Md��1��}�}�̫�r>V��k��g@oC�=�Ā���5�5־�b  `\ٵk}�s���ﾛ��cZ�~=0^�����GGF���c�$L�H�@+����	�i9��닜�5��WI��|]��"���|$;]��?��x���Λ5`���C��r1�R�  0�p��/��~�_��Y~���qX�X��Em{9�̝�p"�5aQ`,^
S�g/k���=7��n���	T&�R�)>N).����C���I�IR��������Y3`���������>�ԝ�= Y���RCCC���@��./��r^���� ��ڵk���'��>��k� �	���j�>�Q�Mq�4G�GFG��<>D�]��D^bE��U5�VMG���yN�wu�Ufd�}�Y�S��ZI������{!��r�cf{�n�QE_��TE_8����R� K^~�e�ӧO��������Nw�u�,�.�x�����e
��Ɂ��g��WEI���Z�2�Z�Lk�Eߖ�!'�JLp�F�-���wJ��Sz�+��ؿ@4�&�4(VO����:�+nc��٦C9�?�3��)�z�M�  �:���u�hΜ9�& ��E���J�u�YfY踬!K>߲���s�����gُ���"��[����D�|�<��[�b�j��ӟ���S���yn}�$��jC�}��3���j�}}����\s��˟��r�Z� �   Jʣ�>Jg�q0�8U�QYϓ����q'@K���˨��~.�908`��Ev ԫ <��\(WD'#!��s �>�.�����+~���T�<=گn�����vl��k�}�~>��\�
�o5�Lϱ:��W��  ()�<��{�@)��X��j:�^��mB"^'s��N:d�_ʾ|�^��|nV �r��3��W ���r�y�筞���̨+� ����H�S���q�����:m�l�>��[�����_r�  PR8�Y���4�.t��TYe����evʹ�eVv �I�lK}��:���d
��
 e��] ş�
��`(9�n������GF���3�Z�(�J@�ye�c��q��ŭ#��|"������~b  ��p����f���" J������Xy�9�k����)*z^x:Q�{���F6W�vٱP������8�P�tԚ�2eH��u�� ]��s�"�Շ�)�+'^�ϸk��O�C�  ���_��8�~�3a�#���m=r��M3ɑM��نz+���:'�X� )�|@�VүH��J�|�����4��YPS���QS|��!��f����v���sQ$ �   JWQ�XP*���1=%t�T��6iw{��?_�X�r�M[ʺ�9��������F���u,�}y@��)@��9V��=���)���J�D۩C�G �   J���	7)�7�Ct�65]�R%�N���g[�àQ�:��Ls
P���U YT
��Ȁ�s�����%AE�Č����<5�F�z���P+�����$ܭ�_�={    �4x���Q��|s�+
ٞ�R�=J��K�w:o������NW<�����`N�SS�d��
Sm]-575SCc����9� n[�pT쉢�6��    `(f�&�F�E�3R��w��8\)Х^J�:����.�����@��l�?�}M�0!.��Q#j��S��g{5��u�^�/��    g
�|��B�F���S��"�ߤ�����t��2���������nھc;�޽��M�f�,�#+�T{    �2$���ٴ��@T��Ƚ�|��w�j#%]���qyٶm�߰�f͜%��T u�m.��6�����[e� �    (c�J�a��
�V�'�Fl�AR�����N�J�v��n�=��A���"5��q��     ��
���L)�I�}f�L�1�u���8<`6�~�ĉ�ώ�;(\���tzm�C�S�^�S$ߏ@�    ��B�թ�~�{�����,��-nW)u9i�$Z�v-M�0њ)W�ܪPr)�YJ �     �s��F�m[n|e�ι�����xE3J3�����;�*��c����ޛʅ}�ݗ    P�x�W�^���ί���!3/�ɷ�a޻r��t@쫌Y�f�    �\p��71i�\x�Z9�{�I��y *�=     (�轜����&��������s�b     ��j;�ƽ�'�m5H=��py�z뭷�Rx��	    Ս-r�X���c��z�O��5+"���p�}�Y�     Tz}|�3g��r�!� ��$��m���i�<!J]]]V��X�����Y  �)��^�Q��L�� � �����׬YC   �Y!'�n�y�����     e���U2XVb     *
���4�JH��@�    @šNd%#�z$_�J��C�    @E��>kVA={�=     �xt��Dɇ�    ��AI�gy7��H�     �S^}���@�Ȓ#�8�3��_�pv�Z��H^#�l�B�#�   T;Fb1�	��Z����7n@�Ȓ%K�P{{{�����h��+�js����&�|.O=�m޲�   �j�)�n��6']��rb     ����m�ܧң��     ��ԛd�@  �q�6]�^Ͻ� �     ��b���266F�`ȖO_-���=     (�(���S\�#��B!�A+b�>�Q%�Ҫ�@�    @Y�J���z�x``����(LH} U�+�=     �5zT�ŝ���6!����4{�l����jb     |�S
��o$�ސK�qOO��ajjl{!��]�MT�     ��8ɼӭ\�	��A�;w�9s�PMM�|5b�&�f�B�     �eϧۭ�F�J��r�y�fjkk�֖V+�^�:I�� �Jb     �"]�]��K{R���2X��s�~�ƍ"J?k�x5�`�&���    �
ѥ��(;Ɉ���cj�yu�bmN�@�-[���	i֬YB��i�l�Ԝ��1��K�    ���&�=���x5}&�\��v�u,��O����{̥��V[�\'��f?n/�:��'�=�    �L(V�[��D���}@��5�s�}Y�GFF�����'����z�������ԛPPLF���{�[.���B�    ƙ��^(�(��B��)4��R�
:��[�>o������Ԅk��7�7�ׄ����jkk��`@��T��#=ƭ�xڑ�$b    PD
��;>_X*sгi�)�ީ��I�����S���r�v^Xڥ��%[�񁯢c�Hoڜ���m2�>�ԛlp{���o�{�= Y�f�ھ}{����/fÖ�[h��m9�K__  ?
�ty카�4Q�[:M.��f�'��tU��(;â�r.�Ǉ�T[SK��V�;��H�	"��ٗ�)S��Ɋ���r��̯�c���@�Ȓ|�����ө���   /�7���DƳmOʤ^)Fo'� U�
㶨�nE�c��b�����`=��)�(�"�V�q[8B/f�5(�=����~&^�ثB�G��(�{     �L�Y�iKOu�#ιT�1��Qw�cgd��Ŝ�ZX�y@*G�嬭R�9®^�vz_�&�J����鲯�%�s�\V��ePo1f��m����{T�    �!�`�E��q�+NR�����Ք]���H�	�X�1���"���ɛdjK� �$�#�j����HQ��;���kr�z5
�֡ϥCU����}#qy=�    @�$��s�o.�J1Ts�������+��\uta��d�y���c>W��ޒy-%(�vt����T�/uʋ��4�J�    U��Ȫ�uQV%W�a���S#�I�c�.#�R�mr�E���g��mB����y�V*�ID�C٣����W��}I����qj'ݱ��Z��+	�L�AU     �$����-]��3rЩ*�Rإ�˔y���Y�nyjn����îW�qJ-Q[��?�&���<�wjo<#�z�D��8�����!�    �N���<�)߲���c��(c�M�N�	�X�Qw9(U�
#��tlF�D�Ψ4����>�kR�qw��s��ug#�~HkQ�+���q�gA,�1�saFK�*{    T%e���R�3���Oc�^WW'"�,�|�N�$��9�]�8�)M�M���2�&Q�]��&�z���^.i0N�m�K�v����\7����U^%��M���fF]_K���   �����.1 U��X��ZW[g�ͨ�2B�% ��OS"�J�[�^Oyѷ;��S4ܵ��8��o��M���2/�^���V���O�QӖJ�3��   ���ݻw�2o	{0`E��."�ʀV���LR.�%5%�A��䥻�KN��<�+��0d�!�"mH?��O�*��܏ERRsFFG��]~ b@����G===R���#  `X溺�Dn���pr�Ә$�u�Y�e�߲��uR�꼫�I�8��ӽ��{��`KA��M&�ש_��Km�6єIVꍌާD�G#"ukhx�FGFE����L�81��+&{ * zH�;\�b�)�}�6 T7}}}B����uV�=`����"�^���%]�E�y����g��S���4�+�����)P)�5Ȫf�y�r���H���1�d��z���P�QHG�+ � �9�}��յ�@zx0ܤI�h�Ν �^8�:K�ۮ���$�٦}d��L�x��,����S�Ո7#��I���9�[����~<X�p�2P6:&��2b�2ϑz�|QQ)��ɓ&ۣ�ȱ �C?�ܵ�@v446R{�w�3 �!g�#�1��(=����BA{�r�T��N@�Yu�VkΫ�\3�T�P���,K4�s����\"������L�|���1��yN��3 ۢ���b{d4��k���MD��+ �b@�280H;v��ݬw~���I|��9 @u�R�B&ēR�}�
�3R+�Xbo���4Lk5J�����8ɹ�߭���!�+�#�ЫeJ���>�i��Kt�����,�C��ف9z?��#F����Ԋ�}��vjnn���?/�= e��uvuA�󤹥%����� ��"��A6e=rq����Q+�oe>��c/��K�I�g�J�C��+j�?_
��KKNӄ�4d4���P���|(�o�ӹj)W)Q�Ĭ���*߈�B�g��+x^�Yhz�t_E�%{ ���
�'�1}0�	 0~H��������Ǆ��N������uR�ժ8������X��GM[
�:�m��N6�<We\��SSV�����HA����ի-No�i=�kd�7�X2/>\�]��R�PdJ�O � �!Q)  ��K�([����RHE��H���`(H�� FS'��MJ�T]I=�������M�0ʒ��y!O������ٰ^���[��l�e� �>������+�Jm�&����K�u?j�ҳdǎ#��g�y�FM���3{    T������)�)�q��x5�c��6F!�r�*N���\�6c*�&�� S����r�ت�©,J���)�5�	96�dj�^쓸���.�꫶c�W��@�!{�՗�����`b"1"k��d)�O.>�'#�ߪ�Y�5�-Ԫ��n�{    Ty�(,OB���+,���s�Qc�81m��	�z_��\��e>7#��4��6�o'���X�:D*QBZm�j��I�~JD�iЯL[��k�[�@�@o�mN�z��`e3�2%r�����a,m�N�~b   ��b�ĉ�}�vjnj���>�Ds��@$!�FrSYIE�0[��T߶��\�>"۷Uj1�����$����Rf�4M+]$�_:�VZ�huW���K:L��n�W/Ȧڌx�y�>��y�n�{    T,��'O)9B�x��(mh$��Ydc�e�{!�A��g�"�)�/�p�*��E���l���t�)$R��b�\�1��YI��Zk���=S��է�t���ǺD��.��   @���˳Qs���O�l�.�,��<��-�D�w�<|5�EY�1���<�[�~}&Y��_�tFf�˼
�  @�a!��0�p�}}}��/SZ��;WZI��L���1�4�
-~��\��S�@�  ���QS J�>C�LCQ���ڧ�TIE�7�4Ą̗{   %�'& J����.cVQ~7(={   %�k���� ~@��Be2��=  ��"'��{�y ���{   %e��Őz  � �=  ��r�q��g   P{   %eɒ%�b�
  P{   %��SO����	  @a@�  ��P(D��~:���[  �p �   J�c��;w  ��  w.��"�k�����'   � �  0nL�0AD�'O�L/���ȯ  �{   q�%��̙33���� �~ǎ�t�RH=  x�  @Ar�!�m۶��Lq�z(� �� �  P0[�l���~  P: �      T {      * �=       �     �
 b     @ �     ���     P@�     �  �      T {      * �=       �     �
 b     @ �     ���     P@�     �  �      T {      * �=       �     �
 b     @ �  P0s�̡��Ѵ�����;�C�H�   x�  @A���4s�̌������N�w秊+WB� �c �   
�'?�I��644ЕW^I�z(���K400@   �b  `�`��袋�_�"�t�I�t�R!   ��  0��v�m4y�dz���'Ry   �  @I��{f̘A�6m"   ��  P2���:��w��  ��  (���?hpp��M�F[�l!   ��  PR�y�:�# �  P {   %塇��;�   �  @I���@ @   
b  ��p-���f���% J�a��Aq1M3�c�{   %����!���H��[�����q:���g�  @��P�@iЅ^]����.^�ϔ�g����;�  PrX�gJ�[�exx���h�L��KU���|_�����K׆*��`0�����+������ĭZ?G}�߀�  (9�R< �K��]�hll�F@,��Մk(��bK hfK�yc$�4֦վ���u���ĭ�O>���}Ƣc�4�mD"�9�y�����$���P;j'BoO�/�c����XR�ն�6����W�\M�K�Cb   ����xǎB����B�Á��������a�`\�����
�4����;*	w����t	���QT��1��P���Vd�ꔨW7�-�ޔ��<[��JiCtn���z~*n��LWF��rd��">����T^��_b   ���#�����2ǋ�pH,2b�b/"���域c	�aX2�M>��=۫T�
�[[������#��,�ra�6��աI�ܿ��Ԕ� N�%/_p��Q�i�΋lO<?�������i������ZZZ���N|��}\@���   �jB680��������h}�&.���%��WSr�"��䞅נ�R���:�s�mkB�Z�
�����������Oy(_�ڑ����SWg�FF��������@M��{    T,�2ם}�#��1��0|k�z��R6D��0l)R�3�k�H��_$���mɽ"�"�m&�>l�-�uz-��*Ÿ�B�J������>_������:!����b�:uj���K���B�   P5p��ёѤ�J�������,�$��y7�wJ��D&	N'͙�eJ�ѥ�JWQ�Ѧ{����Qa����ʆ��	xPu0`�-�-i[|�St�}�]�>}���t�=    ��5��E�l��`O!~�sJJ�)��/ɥ��7���|�*E �͟y�F~.8]����5��u�V�1s�չ���M1��   �*�M�.)lb`�r+#�R�eN������U�3��d{>�"����tU�%ls�Z��� E�d�qe&�>;��G�T���H|�F������Zr�g �    �
dE$��{���2���~4/�hD��2�Z�[�tk]������[]ݖ�|;٤��\��/d�t��"���r��E�%�g�?C�o�i9===B�)�NV���߰��Z��A����ϭ��F�L�����K�����?>�C   JK�+�"#Jm���	�b��}$^�Rԧ�΀��5W��ʭ^S]�8����~�5����l�f�_hdYp+�܉��&�n8�6,��keQ#�9�aSTLb���cTZ ��7,YPO��r�3=��x��C{  �MMM���i	���s��h�N�%���沖��bN�h�>�VNb����i �ڱH'�j�_�xd#����Q�B�t5C/Yj�6��$?��V[Wk�}���=    ����Z��������=�|2l'w4���hM�t���m�Y���Du���3��Rc�D={]�3��Ѩ�8���SI�u�!�މlR�2]9���W�^��9uK)yYJ �    �*&L�@;w�ƆF�7b�Q���Y�y�鄂���+r/��'��[)��i�r��S��u��;��l[�G.�m�����D��6�����S�9� T U�]  e�WGG��d������쪼p�{9��J
	N|�Kq�Є.n�VG 
Z3֪�[9���c�ꀞ߯�~�J9��ZeӤ������v�R}��Gp�i/݀_����r�ܙ�)U�=��?N@�("S&��W����-ZD�V���NL�<Y�aˇ5kֈ(  �3\ɤ��Y�F�9�r�Q������L�s!�	��y��Wኈ}B�j
����̥VG��4��?w*�m�0X���]�d*P��#��c�H�Q���}Q�;E����g���+�z�%�f���?S3^)Iv�,��Χ�@�("Z���SZ��������t뭷����O�6m��?^̐������?Q[[[^�8��hŊ  ��rKKKJd�c��	�Xb���߫|˲�F��"�FG�<����`H��'���'G���ʙp�"��׊t�@�64��}�mu /�mp'H�VrjC_'ѣ��.)E�ґl�?�)@�(2�>�������-���K��k�Rϸ��?B� �jǩl����ɇ�Ɉ��v"�Oʾ.��Xv �>##�"�G�z掀lOD�U�5���,�����\r��R��4ly,3y�8 +
Mڠ�ĺL�
��YPR���zj�S@m�m o&\;7Z��/�4���a����8�wǥ�L���1zj�@Q�u�y�ёG)�s��s�9G\^�ٽ{7=��Ct��'  T;��ˀk�Ny�PDl�"��Y�Ul �{���Jv �����J �����4��UzBA0�S�PSjgEޗ{X��* ��c �&�rJY�S{�Ы篿N��:�}WS|+e ��*Ӥ@ٱל:��T�c_r?�Vu�l�WV'7������>�z�ӟ��֯_����N'�t���v����?��G?�Q���  *�
��URM�(��~���U �i�+�� j��[3�ڪ�$D_D�#�ȿ3���p��s��5a����P�r&���O�<����ɩ�9':
�����@r��^H��v%@��U����̗J���@�Aə==L�
���{V�B�	���L��\��V�!/�	W���j�K�^���/�s֮]+�;����Z��ͣ?��Ϯ�c�, �P�^}�X��|�"�6�]!��nXҎv���oY�m�@�dG���6�� ��d�}Y��I��&jod����x U����צ�N��L⨿^MȺ2�G���K����g��J(�	�%eִ�����ޖ���hl�u�M���}m����O?��M�&��4K~6�u�]��sZ΍7�(�� ��ѥ>E�lWD�)��u�L�W�Qoe:O m�5�m)@#��}5J.nɰj��J@< v_���Ubb�-:!\(�����Z�{m�D�e����n��/���Y\��9��f�*C��ګ	�=()'�L�C�%�z?��&��ݞ��$?����g�s�=G[�n��S�����詧�"   q�f_ͷ-�ԞldT=����K�E�ՈxL��55�� F\���i����jl��y2/����� ��	����0	��ui��d����2�k"����c���EIt�h��A(��= F.b�_�<��t˜r�){  p�+�s�|��ip�L���lO�q����·*����e8b]��Zx�|}YH�1�~�4�� �U )�r�s���b� >?_L
�NN������= W���g��/������۷  ���U�v�-׈�+z^��U ����t�^�*�}Iiw��$�ȫOL�œ��(��E� ���/&�
�'�b����P�#"g�u*Q��>TH���
#�A��7o�W_}�8� ����8��?  (>�J���P��f0�=ΦDe���q �$V2����-����vxd����������phX�=w�uVGBͷw�WM깚H� �	}��l��_�*Ğ�4i  (�D49ud�����I�O�*��U�	�����<OKWW���Sccc<-g,>����0����+'~b@��O��۶m���$  �� ���`+J���Ċ�mQ�j�>VC���� 8�/�r&r��BcV>�א� f�����rA����1   P9��v�_�<��$&�J��'*�� �9s戔���AjlHD�r�1�LdUn@��0��s���'�   � ]� �+ b0�2@�Ysƌ�a���å.���:p�-�F_��DV~b@�q�1�г�>��s;�0�>L   �����VZ����˔)SD䞯Z�"'��}>�L9�\3ߏe2!� T���'iݺut�-�d�?װ?�裭��    �@:qfigX�D*���5�5Y�8r�+��[U!I:��mA�(��I���F�a��-��?��$ejk��H�g�m�����=���ė�m�������_/'���ر�    ��N#s�9uh0^�ٚ��t���T ��b`�k<&f�������J�=��R��w�o㋜V����1����س����t�GX���oӱ�K/��"uww[_�,����b2�������C=D��?�C   �_Q_���i{zz�|Ӿ�q��J�~�=�x^~������~�]����~�/��cאi���\����ϧK/��N?�tk�Œ	�b����n�r4  ��P�krN=Wő�z!���LmT{P�f &��T�}ǻ��/�Q��_fW_}5�^������]�̗��s��ӟ�����\FƄ�  (!)���c�WMF���Z��؃���$����=���K���~�ZZZ�����I��z��$��Gy��Ν+.u���   �)�)�{�˾�쳕�Tn���כ��k��������=m�'����   ���;S<[h[e�T.��Qʃ2K�   ������+�g�	�=�x
��6a�   @E�i2�rb*��SqL��=    *k6�
�{�=�xL$�>�`��W��I[O>�$�}��   �!�F�.�\b@����~��_�T�3��/�  @Y���WB�b@�3g�1��WR�<��c   ��JK����
����n��f�8q���{��/�Pp����   ���c5�Ưi�{P�T��t�hjj�_���4c����k�E�  @�c�w��"�jν�=]t_-�i��{P�Bz���SMMؾ����Vt��Qփkjjj�n����O<���H��~;   ���b���:h6��;���]v�<�؃���Ɍ>c�h&��4�g��~A�m ~+b���}͊`0H�\s-Y�D<����NW]u   ���3͢m[�H}�m��=H�w��}ԤYQ��i�
��]Q�*`����6�����}Y���{��s�1���իE^}$!   �R�E�))�L����[5Z�$���rb�1,�#=���g��z#�����1���FSa��K�g��/��Aeg�_����SN�w��M_��W����   �J���η	i�	}��/����u�L���>�t��{����B�����.���'?��o�w��y���?mM@5<<L�{.m܈�%  ��B͝����&��Y상`b}��	��G�ԇ��_��t�H����f�#o}$6�h=)�z����������~���cN�Y�l   ��*�R���3K}(�G�FE����� ��& ��S�ϨQy5R/��0ʧT&��ɨ�Ν;	   �$�"����������("!ש�,%f�ľ@ �>�%�n�ث�[iy��'�)'�g������>�1��/�K�o�t�R   �}��L�QoY�9���AD�Y�e:N5�/ H�����9����1����> �`���LɣW��H����7��}N��SS����?L�gϦ��?_<nhh�_��Wt饗bR*   e�[�5Z�z����m���4}�t+b/;NQ�Jb�'�z�1��hp�`��6���zW��?T��c?؂Ω!�+��@��|}}=�y��1OR�����Z[[��   �A!�����z	G�GFFhB���Q_����H}ya8��8�ۄ�L���k��8�]q����D��z+   ^��|���$�*�Vn��}���4m�4
�C"'��W*��ԗ�dӆ�^y\�B�r��׋��_|�����o�E�=   �Rh�Z�q�6���c�^x5J/o�}Q0"�'~֬Y"G�gV��A�s R_�X�fn"�1����������N��(*0�s�Ƚ��k���  @�L����%E\��C�y�CoPj:�J=���e����fb��[#������,����_�O��Bu��W�l����1����g�ݵk����z���<-X�@�/�|��y�  P�;��(�w����4ٶ�v�TK�)^�~˖-448D�-���&!���YŒ��H}�x��!��U��˧P}	�c��pX�/�z������]��szδi�ĺ%K��.w �  0�xewKy1\��Cqu0���G���H9m=�<��Z�\��s�8K=�Ȕ�#��ү+�y��ק��!�����o�`�v�$*���~ɝ�R���Kz�Ûo�I��v����'R��*  ��(t`���B���~�vd�He[��o��N�v��~.�cy���Q��̏�������������߇���S�5�9���Iͱ�����=�@�� �?X�9=�}T��J�%�z�e0eԾPv��A   2�V�݋6�D:[���\��J��i_y��z:�~N,�r��η,��N����c�jjk������9OTzS߃t�,s����Q3*n�^���ػ ����D���zA��^�_���.�G��,(
Xj{��q���e<10U{�t�t����\�i����>����΂�H�\�#��3����ۘ�775��b�I|M�F�̫��5]�����=���K��x&��{b� �x�� ����?��lq+��϶-!����|v���\�Kc)�rG�U��e�`���)�r���yMS�-�.��;n�3�:u:��N��٢w�� ۮ��,�b��^22jB���  JM���Txɶ-� &nU��'O�jW{�� Q=�iQ�]F�9�^Ә�pMX����d��9�N�C�~N皩�.=&�Ύ��c�(h�y#`�.Z�@� ��k�Q|� �700@ �]����L�B�V���ɔ�v\=��$�z��o�=���������+����¡��w���y�N��������X�ڒ�y+-GI���Y�� ������. (�d���"�������)}�-b�N�ݢ��:�躚ù�c���\��ƺx�=�D���į*p�P ��TM'��V����n)8���v�1��Ye�uJL��%�z  ({� J�.�R���z�=]���I읤^nS��n�0a�J1VzL춮��&�*�D�ӭ˕l�/�}��+��TB3�sRSq��4�?����z�jI��z��� @i9���ń3 �
U�墊�S�7���y###�z�z�]氇B!+��b�%ET=�r�y�S$]��W��G}n&a�$�ْ�S�_���j��>����8�+B5��B��/EĞ���z  (=�~8�_�� o��^�z��Dʞ.�jv����΂�b��IԔ���8�Տ��J��~��Hw�v�>��7��V�s����?wqL�����V�!�  Pz�>�h!;���
=��v�u�g�SbD
Lc�-®�ĨQ�l�<�W
2�.�=��m��1�+ר�ɖb��g�|��tyl�~Ñ�H2R/;pb���^F���k_�b� ��Ñ�s�9�֮]K �7R>���C��(��Qt���z+=FT�ID�e��U۔�K�$���i�m�ҵ�UU�b��}օ^{����ԏi��"�ruJ�>T��C� �\u�U��-[��?{�v��&��^H��w^��
����}^� T��������)b��oZ�S�]`����X������i�lȥ�|��U���k=:o-�yK�m�d?2�/��`esN�EU�=��7~�� ���o|���Z�t)0ް�q������2{���.n)��/��N�1��Eϗl��=G?�t�_�:!�c�΁S��J$d��_IX�����z���"oFmm�>oS�W�>R�9:�y������5<2L��DjV"UGΦ[j����ԃR�sz�6���_� (����L�B���?�J ƛ��N!r}�}"�F��V�2���d�w�\v�H���9��E�3	�-��A��0��<�(��)Pnǔ�82b/Rp"I��|u�/���b�s�����?Pb����T~u�T:�{P�pJ͌32����'�H)G��V�T,ai���b�Q��1�����٪Ȓg���w���r�� ]ĝ��Qp9ϙB�Hʧ��_��>�U�ƌ�Ȫ���ؖ��1X�9}��=o*^�!��C(X�i+���@�AE�)5۶m����-[F ����~1��-�=j:��.}"��TJQ�᳭P�&�N������d�kG
1G����B�[���&~2�JM�4>o3~��#��5<��Ɗ�8�2N��H�����q�������R_>46hɢZ��a�D �����,L ��6!S�dTYF�Ձ����ɔ�Vk>ƀi�l�E���v�|JJga�<��x�z�S�^V�����F=�����7��������X����-��� u,�|/�-�D��Y�쿶�L	�X��ԗ,��_1�ښ�-���g���?�h@� ����$-Af�z��Z5�Y���y�r�l�I"��T�2���nz�]=H�e�)?�t
\�(�"�7��"'n�`*'����&S�u�M�)�਽mfY}�E�!��9�<n�/R�T��C��)�����n������� ���&�U�^`$S2d������a�<n���n�^�t���j�L��"g[\%����>�����Ӛ�5�9bY���k���R6S�x�t�#	���ȷmmmV�Od���R_^|�S�q�/"�"�����K�Y������w  ��#�2Z���"�B��T�Ϫ]$#��oD����7#���
���ш���UWde���o�������ێa���E?2���@��	L���v������X�yP�I���gI���*J�!��GM8P�cĿ؜?�����&�'_¡�(  ~��3��Y����1G`)q�؊�#B�E�?�O0���J��S5w^KM�I�E�<`Ӄ?B�H���T�6�c$��l�ɫ
�.%���N��Y��S_�A�Ι-��tu���Qccc��g�Q1b�n�t�~y���z   ��S(X�m/q�}쟸���H`$�����-�>C$]s}Q�L-i����e
���ɫS$<�R�|�x+��Uu��8$�ܪt�Ll�jd&KX�}�ف�����i1�2�B�W*B�!� -	��?⊪zy1!�R�!�  Pyp%���3��ur�5��Cn�N.�ێ����6_���7/*�1�8K��n�IR+�0R��q�H�ܦ�So���m��3z�L�%C�2̲{H=�D�%b����ddFF��|�  ��@����Eu�u44<d�.#���E������Hp"�D�n�(�<G��0jU ]�����D�3Eĝ��u�;�\�J���R�!���r�E�����擉�  T �/�r�{�njnn������O�6`T�u�9W��6�N��X9ކ"ݦR��t�J�YgՊ<�,��-�Yb�r
I6bn�s^���)B���\�U�G�l�R_yBT?�)���>�CJ>�Dx�^Y2�jcX)7��y��3��S4h�   ��k�9����T[W+��ZF�fg�`Z��c"",'��G��b�:�i��\���+&����<��Hw�P�b��P�Tߒ�ˡ�s]��s�ޒw�bS<$��"�'v�~J}��4ʽ��  �?X�'M�$ĝg�f���Q!{4>����"�E~v)�B_����C�A��#��5�ΐ�F͸�Gq��X	�-T�  P�p�JCC�m�S��I��D>�: �AY�=���ؘI)3j������X�crϱ�{3a���  Չ[�|��xQ6b��ۮh�ԃ4�����+S���c��q��r/Rp�N   �H:(�B�ԇj�K���z���炫��b/ʇ%r�9G>7ȗU�DG �z    ���T��Ճ���3��m��	G�@Y�Y<�>�X�\�=g:�    (|-��z�o�o�����̲��Csg�D�=    �ߊ=�xO�1}�tjll��9o�&    �rb����    � ߉=�     ����C�AQ@�<    � ߈=�f   �2#
�Y�sz� H=(&F ��P�&    @1hnn���Q࣮��jkk��3�ã���iӦ��+��C�A����d�    �[&O�,���&!�,�7o��+W��իi������o��~I�R<��č<��z    x��3hڴiB�{{{�Ŀ����s���Ȉ��*��C�׸�8�(�W{��   �3�N3�|�f�2����<@�=.� H=O�<k��ĳ�p��L��I[۶m���p���F����O�֭��� �Jd�����3gҚ5k��+��6�۱�]�!�`�	�1x�#��rt�UWщ'��I{O=�}�ߤ��1 g�u���_�>餓�����aq9�E  *�<�������=�\ڸq㸟ø�=��ԙ��Qz��;(N_2J}�@�6�/�R�_|�gR�y����~Wt HGWWW����'?�u��կ~�>����b��. @93a�z�{�K=��t�M%;�q{H=(6n
~�~�t����s�6���F�M��>�l���?�y���v�H�)��<8%����'���������-  ����Z�h��W��Gy���2.b��$�a��G���K�/���O>�����������-[VP����_�R��s{�v��￟ ��_�.����OJ���H� �%<ƈ��z��b��E0`PM��4�����G>��*ö��^��}����'GA/��R��_�Zp���\@�]w��������M�?�8�%o��=���t�A��/�L  PNL�8Q����/~A~��b��I(&��#�n���|F���Y�fѵ�^k�P����}�Q��������_.��87��7�D��n�A\��{� @�0{�lz��'�/M�!� ���v1�4�]�s�=���{北�>�=�Pq,>&�x��А(ɑ��;w  ���K/�_(��C�_˲m $�_������* ����o��6���R   W���/  ���T�!�      ���R     @��D�!�      ����R     @�)H�!�      ����R@���~�     �$/����ؾ3B��o����y���v�߻�����i����%�&�w:&    �E�b�^����MS:Bt�q�T��n��ݞ��b�
z����c������[�3��uvvz�~kk+�x㍢m�駟��+W    �INb�^���޼K�?�cmTɰ�_��.���:/��b���iɒ%4{�l�կ~Eg�y&�v]]�hk޼y��k��F^x!E"�w�   (�{H=(R���[GG�D���R/��}�kt�w����E���~�;ڰaCA�Ι3���w_qժUt�9����   ��d%��zPl�#����W��K�%===t�Ygѝw�i	���Bٲe�w�y�    �7�R@���=VT��p^��g�Mw�u���{���ݻ��_���{    ���b��0�����7
�?��<i��G�u��    �W���P~���b   @��(��zP
�Z?L���nۺ���Ҟ�k��X�n�V��O@�q&�   ���"��zP*^\9(��� ��LjmP9��t�owҳ/Vn     Wlb�OOMM]}�մh�"�+�=���G?���]C}�~q����z&2�?.젋��A�'��/����u�]GӦM#��eJ��   �/��C���R��ґGI~���O���Z����O�h�ʕpؠk.�{�R�����:�?�N�\>HŢ���n���1c���{/�v�mTnL�8�n��V�{���\z�d�|    ��C��â|����a�F���'�,f%�ꪫ��gt�7'����\��1��ߝL_�j��zq&v�	�>�`/Z[[�����[n�ŚA�ϰ�_r�%�w�{   �z������K�/�ԧRWW'���r���ԧ(�]�>�6t�9����ܩ�5�?�3��z�6Z�����X�����f���CSS�M �ƤI��7��MYH����{   ��7�-_��'No����~��_Ӓ%K�)����>?�>qL3U
M���S��m�7�z[!��_���ޟg����(�Z��n��ƌ��tWRnL�>]��̚5��D�  �K(��#�u['�^�#�7�t-^�8e���(]~����+��_��G>B��ַR�s�)�?��V��'Z��hr?�ξl+����v��{,�~--����1��~��{���n�{�i�&��{.}������{r   [BRhnn�����v�~322B]t=���'8� ��s�)����?�D�}fU*\���WM����~æQŁe���I=�̻|�r��]v�i��f[��   ����%G�ݤ��.���~��G)'��Ər���7�e緋��Jfb[�n����w�Җ�޲�{���)S��l��줳�:K� ������@�w�{N�a �   2�W��_�pa�6N���K�M�߷�����
RU0eR(&�����vt���=��ST��<yr�6N;:��3i����W �   � b� ]�롡!:����^�r�����SZ(\e��Y�Bt�Q�t�}�	W�a��Җ:;w��z?K�r  �P�L��iooy�Ne��_�j�H���2���\釥�g��ٲe��Կ��;T.@�  BՋ=׺v�������Σ_|��Ƚ������Ġq���6o�,�~�ƍTn@�  �KU�=W�`��={vʶ��^��W�B˖-�rr�OJ!�۷o�˟�W_}��Ã�ݤ��3��UI�\��  ȇ��SN9�Q�w��-���̞� �=���^����;76l�j �R���R�=W��z�S�N�5k�P9ÿ�N�7�ׯ9�[�n�r����?�!���:ֹ���{   *U-�N���K_�7�x�hǨ	����A��葑Q������M^�c'��t
��K}��2^�������^�����R�cǎ���&L�-���D#�c��3@C���O�W�x2<F�{   @b��0����6L��I{͝B�gN���F���br��NZ�n+�xs#��yz,�<Y��U�J�M���j]��y^�=r���?�yQ������;��܃�cR��_o� mܴ�V�������<ꨳ����{   ���k��R'Ml�#ݗ޻p��(���XG�Ο.�����|{=������N���,U�x�F�MJ�>�rU����{���ɓZ��-��̢`0�q��zZ��L������6���-�
/kZ��   
�,Şs��ϟ���/��a�\mm����B:d�^d'�y��!�e+ߡG�|�zz	����:U�3z����¨~!	��/���.�%�wg�;�!X��,ze�:z��ר`�   �bR�b�ᇋK�:?��Ϭ\�R1c�D��'��	M����=�i�^��O�H+�|�@v�Boɼ���Dz�X/�NJ�&���=�ޟ̜�N��~'�5�����Esi������������  �/e)�~e��3�d�v�+������<��u�R1��&�fr�i{^�Gg�T�����	�7�m��B��@��wp��I'�?���\il��ϝ�z豗��^����   J��#����?���	��G���� =���	$q�z'�g�7����V��|k$�� %�ox'��?�޹����_ԟ#7|��%
i���"   �k �0w�d:�ă�*�*G}p�o��u��R�tYu��XG���$���D�zPgL��o�	����5�S.���z�����p��������'>�d�~&<0�+�p�   �K ��?��CD.�v��n�������k���z#jAs�����'�.��RKO������[;i��nI�Qy+dO]��t�Ǿ�SO<����2@�%sr�(=?0��s��D�#����T�tZip��S?~Hփ�c��#[��~yphtYdll�A��X�~^]]x��I-����ej��}���j9�:{	   �
�}��p쁢�]&�n�ݳ�������nL��>s��ӧ�ݼ��i���<�O��~���'(��Rx�+���^��DN����q���92�^?^N�^&b_�pjW��Ħ͝]����������;��cN�9}��f�w�ۏ'�����[�|�d��  �<|+�'�p-^��q�ܹs�u�Q4c��m۶m��o����'��A�ɞxr�e+߹�׷<�oٴy�]��o�f��>���-�sYL \�+�,Y<�^|y5��h}���m��h=7���Gc�2	����J;{�զ�16��Vn��M��i����/vs�W����-��p��J^��N��3�^[��    /��v�a��<��p�bqb��՞����_��,��ʚKn��krm�7�}�{�9�C�\r�^j��u���a��K���ql����� ~;l�QC�}4&�AY!G��\{T�)=:bA��#�zeٺs3]es�o{�g���/�������_ ��T   ���b�w�Nn�t��lݭ�H����~�����K��z����1���׫s ^�Yf��7��i&+��R�f�� t�pz^��{���;�3gΤ���7ߤe˖Q%0{�$q���Y��l���z��w���3C����{]�6��g��{ϩ�j�   
b�'����v������>����:746~������A�}��v����&�?eI�h̾3!�B��W'���(�1o�<�馛��8W��W������ݾz��7o�ݟ/(�8�����45������ÿ�{   ^ �ϓt����uK��:��������676�9�^s�Q(�H�8j�>U��L���T�>��8^����b���q�J�K\���і�]���X�v�<uάIk�k��]����  �0 �y�%.;�[\�oܴs���>��Wǻ�ާ�M����}fⴝ�~��vZ���fL�H����l�P%7[y����,\�y@�9�C�gϦl�2e�؟�N���m�A�w�}�����Hm����7lܹ�?<�^����n�䎕��=}������2��;   �o���[n�|�q�GAg�qF��?����c�9>�'��
�#���vu��/yLw��-��Cܶs�n���W�y3a�f��7I�ʱ�Ē,�R�/_N_�җ2>�����.]J�����o::�����1�������m;��B�  �o�~͚5bq­��;３��G��1<y��c��l�m4:�f�����x��x{Z�EqJF�������{}̡H�vJ#���	   (ߊ���K�i���1������{�XsS�cy���̓���O�1Q��¨��n�3�zjVz}LN�;쀽��Z�y)jk�U  �p��$�w��t��	�v�#���i��gFFFr�_͸�NϷ�r�\g`��2#r�4jtt�|��G��q��H4&���	�  @��I�F�\���L�'vw���m��qˏ���S5��������������"2�fbFٸR�;3�}HT)1(>x6 ��|AI�ɻ붚�����3��;���1���5�=��Q   
b���z�1�}�؟z�3���g���"� �A#Rh���9ӻ):f�ҕ\R0^U0^^�txj@��F����)䞋�#��td������t �ڷ�z��Cܯ���"  �*b�;w����������m^�����t�wu�Q5b�8��a�}���� =[{B�A#1���G/�7��(�:���p�8oPvv���m���rA��}}}�7�mߕ�   �l������b�`�9�}��C�>f����m߼���='��#�f\��7M�*_�5��� ��r/��r�B��sgx2+���Ɩm]�ΜƔ��#�>f�Ė��۾�.  x@Y�����7:��S֯]�v\��3S���N�;g����I-�g~�#?��w�~ǋ�}N�3��u�޾Aڱ������'����]��,=(��p��6���#�>�s�.䥘y6W�~�m���+頃�n�����������S'8n�:����~������ϼ8��>}�f͜�ᶝ� t�x7�  ��,Şg�䥔�|�]W�g�ϛ������=�<����|��Ť��@�J<+�|�1�Z��qJD�)�3���	��o���F�I)3��h=9H��/��KO��K�ÿ3nb���c�U'�x�M>�|A92��ߺ��N��t?o>   ��R������G�\�ZfrB[S��)S^��
�s�1�̓E��>5k��t���l=�8��'�ݒ{� +�L�O&�F����,�ȓ/_^[�����{�m·ɓZ���3�������L|�� �m�����   ��<��8//[G�?p��>{�1y��'�8��K~���������=��f�n�5�Ѧ-ȯׅ�-�L����n�|��yV{Zꍡow���	(!���i�����3޴��q�'^ڼsա<A\.�sy��-'>������U�h�N��  ��}<���iqLj��9�i�56�njkj�ԝ����l��짎Y8c����uf�ۏ�����N�)�M���ےےcfS#�y�%Pj���JZ��,�A�̂}f��T������w���ٴ{��:h�g��tLM�_4�'�]N   �W@���=�������oƴ�mS'��e򤦕;vv�t�}���Sz�>}��-��Ο7�p�('�����Zzw3��nXUr�F��'��=Qk��O�AO����9?���7{ƤI3�N�ۄ�O��kW��~��'�v��s�}҄	Mϟ7��pؽf���W���   xľ@���U���i4o�)i���>{MOl���o�-߽��kd8�m��XMm����~��p�����~�Uv�0��ט��m�l3����8��y��7���i�����DZ�]����������ݱ���pxBkkÄ֖��ޝ�EU�a �eSVEA�}�J3�4�3KTDDMm_-Ss-�4�J��TD����45-�ܗ�}c�E@����=8��02w`fx��H�w@��s��:�{��x��   9{=q9L�փ4ilr����8:�Y*^���U�9�]_�w(77�@7e��~\9���U���ؤ����uq����89�[*^*|�r{Z�~��+��  @-{	�B�u��ф�^:�����Υ�Q����3���������H���ˣ��l������Y������n���+��n߹G   RC����^��ƌx��x��9�����?̪.w�_��c+{��`k
�9�T����i���,>|8��ݛ6l�@��|��|�[]�9RogR�"��T   ��`/!���j�.طun�'i <�&m�v��g�9�vGM��Jd0��¾��r��Y
�?�E��wt��]����\����w�mIz��gc��G)''�   �^����^�u�?*~��3��'ﺵ�:w�ر���w�/.����3�-;�^���`�p����ax�~�'����zKЁ?۹y����t���T;�����]�E$�u[[[  (���q���ѣG����z�'&.��\����yѣ�Pc?O��,����n$�ѓ��s1TX�G��O�Nu��!c����u�xɭR�}eA�7���{�.^�(����m�7�R�&��S{_j��q�ZU�s�����B|���*�,�/&  ��T�`��_��ό�X��^~�e��=�:~������ɧ�y�;��S�/lk1k���/:e��fPl\*]��H���.T�2e
�=�$����3r��bd�Ku����E�h�a�z���N����i͚54~�xI�=�q�S�/��6���I�]��͙��ׯ��0sy���J��Ч�UE��E�R�P�l�2�֭[�c�r� ����~�ڵԥK�ܹs��s���/���_�}��I�\��F*!!!j�-]��n޼I���?�yo�G���+��G����L͚5#oo�R��p�n�:q��ʕ+�=��={>V�TkkkZ�d	��ѣ�1�|�  ��j��ǋ/�(B�j��_��~����*���+4i�$��>��3Z�z5�]����{Ӵ�=B���`��;�Uý���x���2YZZRhh(��ի̱���6m�ٳ�   J�����s�饗�צ�ʕ+髯�"c�� �����7������=���>I6��7��\�=���������S���۷  ��j�9�{.��u�p��#0v��>7�}<Ճ�M�'���[����\��z^ ���?  �:&�˜�}pp0���;j����ѢE��T�q�>��Q-T�{k㟹W�� �Ws	������W깳�|@۶m#   M�K0�pϻ����j�������8���ɴ�=�����:�~Ĉe�q��7om޼�   �A�Wa��~ذa4{�lT}�����:}!�b�ɯ�5���|:vV�6��;S��=&F�Y���?�����	  �<�j�b�:t(͝;Wm�߲e�8��F9Uű�}>�˨C=�oM_��W�$QzFA�3�p��oj�c�7����$   ] �k��[E�Z��ڶm[��{��.�&V��\��U�3���/f��m�c
�,�YԲ���f�6�b�'�<'Q�M����)�����������o��l+}���[4a���x-/t  ������◮��{ClbU�����Յ�;vЬY�L6Ի8Y��<���i�z�G�~�\/zi6�}U�pϋ����j����B=�1�P  ��<s�e,<�meU���g�n���t�ΝJ��x6��_��b��p��y�����Ǎ}���F������ˊp�Jp������?/s�g�����U���k׮��8s挸S  ���Q�n]��]]x�m�y�[U�z��� :i�������������޽{dJ\]�~���Y7e"�+���f>�7nܘ����ĉ^KaccC���t��y2�Z�w��IMM�)S�T�ݬ������Tպuk1�0g����  U�^��z\���5����ě���Y��F5�w�ؑ���Kz�L&�{�Y)°'5�cڡ^�ICZ5ߋ^��D�ws��gϞ�l�2q�[�Y��B��0���/�@�2.Sƥs< �Y�f�c< ~�������T��/_.�]�>U=�����wS��  ��^???�����ӳ̱������ɓdxӚ��\ѣ��@I:tuƓ&M��;��r�]e����ǲQ}�V��E���'����|ă?^��`��RՃ֊z�'D�:��Q��9�p666���	ݿ_,�U5d�qe�ԩ���O   �1�%��͛�P_�V�2����E�?}�4��;wRNN����0PR˖-��ó���#/wK��/��i�?����{qV"�ܖ&�;;;� koo/�޳g�^.���K� �ˋKϞ=K��W�^�dɒ2� �.8'N���D2&|W�g�����wx�ś�q�  �6晢����\��G��r�K�.�1��<����e���gv�D�?c����a%Bo]���q�6�-3������K�ũ��cJJ
͜9S�{��1c����������ƍd
('�w���˗���֭[d�x@��}�=T݋�;_�݇7�xCܙ  ����N�:�ʕ+����-|�r����_��wUK�5k&z{s�7��Ӡ��(S�p5�����W�qR}�ʙ�[i������O�>�o�)l|ׇg�y��ڵk�;=�G�&c�JÇ]�Ե}�<So�w�����ğ\W��u���C�y��p  � �?н{w�����\.K���#S�7����nԨQ��1^;�5�\g���LU��I����y~���^�R�|�z�4q��~�Z�s��	J���(Œʵk�D�E���������ȑ#ŝu��رc��K/�=)L�{�s�n���F�`^��0   U�TT��=�����\��OJJ"Sr��Q�<y�(�P�ѨQ#�y澪�--*^:Ru�^S���~� _� @WV���D9`���Jm˖-"�3ueiƂ��-<e�����8Քl޼Y������Ҳ�1�σ.n�ij_  ^���R���;wN�T޾}�L�������W_}E��5lؐ���)$$����ɜ����o�I���L��cK�y�½�D������\�Ã��|�j�L<������ӛo�i�e+��g�C��M\2�״)�� ��Q��}߾}飏>R{����/Nc��-���;<������y��̾{�.�M�^�Kה�e�}Lq����|[]�
��|�bj^\��鳳��}<w`�au�M���P�{;pi��w���_ğ��=���R���`  P�����Z������e6���W�{ղ
�������P_&���>�_-��K��?L&/����$6�l�K7���>其��tc�|���w߉���eS'�<@Y�hQ�RA��  PR���p].� C.N���!�dgkM�����G�Yt7C��V���nذ�̂ZsT&��K���FN�ºL��_���)O"+5s/3�j�b�+{�0ȥ ��k�9����S5kؒ�S�U\�\����~��ާ�{��	��]�v�u��  �6�*8�K�k(�|������wo��!6>��\O�3��ҝti�\�pA�ds�rsSj^M�/���%:T�eF�Ɋ�pJ|1�/{pn#	��6bR��I�&������|nc���d���	�5�����ȓx�*�_[����Υ�8��#�@�;  ��ހ<ݝ�ɮͩeso�R�n�� r��~����I���z�q�7&��d�/,���*V~̃�.¼�(�[XȊ�s�p�<U�֫.�V�7�R>�K�x�Ey�W܍��ё���^��G��Լi=�%{���l�i�:����m��围��sb�  P��Km��lM���U����e��/�/ޤm;�ѝt��S�Lm=�K�������D�/I�\0++
��x@��5�%?���������um���K��wlx݅6<��B��p�M�>�]�������g��vҠ�v   �^b��h�3��\�4kZ�����mG���X��/��R�^�`�^�9��v��)��kx���BM�7�֗��w���b5��J0`@���cǎT�6����=���IvNQ��ȋ���o1�  `(�j�����߶X��vԳ]鏃���=��+9[/ޖ�K�z���.T^�������5�E3�������r�����k�9�3ދ��~S������EkĒƌCG���{��=���7͛7O��_sDDU<C?̿�Ne7���tW\�'��C  ��%Ү�=;�Q��/t��h��۾4+5[O����`/+��/^fˡ�̾+�Ǉ,G
������/�C�
���N7nnn��ٳg�Y���������C����x�b��СC��yyy��իETƏۺu+��.�hp�N������7��   RC�� w�xfP�J�I��DK���M��_��Nm���g.נ���{��R��%>���.5Өc�po!*(�m��½ʷ�2�rx7d�_~�����E�_���{�]�8��=�T�s�I�\��%<��7n�K�.�����'�?�ڵkŋ��:���;V���_�����~O�s�   ��`�''G{
�{�M������G�����\V��|+����u;ww��^�.΢���������t3�6A���*a=�=���u��ϣ�»da)+Ȫ��^.��0�O�F�i܍5&&F<�g��cx ��?$$D����{1[o�j�Ԥa�u��@rJ���[�gg�+((����(����������������Cy���CvT\�i����p  `<L"؇��QӦM˼�Krss�*�?�Qt�(OL|JJḼW£vGi{ܘQ�����޷�G#m��?J+��ir	�\��M�[�+k蕳��R����&�tO��ƛqoze��:�w�ĉ)--M�p�����5�g�g�Q�c荞��Ё�E���܈MI���:iæ]?i{\��~}�븬i���[�τ��=�߅V���  P9L"�s�=��!r	N�G�i}LAA!�r_�j�/u9g����oHP�)m[�,�ao�1xy8S�����1��B�b�?gF6[�ă��ӧS\\�h{�NTT�8�t��U1b��a��G�9VVVt��=:~�8͚5�������bw�����+��w���o�r��;w)��?>���Z7�ikk���~=Wj�ʇN��N   R0�`o�zuo��x~~=~�����x�s�۰�#�:Ѧ��N����|x��'��H��_M=a��V˖-{����Ƞ�Ru���ߜ�<��cWƆG����_����cF�9ޡ���54�{=тN���`!7  �~�+��W-jX�]�q�'���yEB�RX�o�C����ܾ�:++�ٞ��lV_��Fqw����h�0�C��(��:�.��]��n̯H�W
��������4�T��ڎ�ԯ.��O   �B�����j=~�z�կ�mM��Y�qWXM{��6�|���n��`/!�2��3�Pofڕs�^����ڍ;f��<߄��ËCG�x��1M��r{  ��}5���x��b�neK�\i�����Ntt��Tw��Ǔ��,E�Ou&{���(���0^�<^����y��_��E���MPS�:��������z�[I�#��w���$�������8  �/�
����\�4��O���~@��۴i_��.�Z6��M�q.��x�n$SuU��U�鑑D����E�����(&ɵ��hS�Il|�刈��H�|[����r>ݼ�w[uǹ+O�Z��F   �@�� O7g��S��jm�W��d~������nN�2ؗ
�*��l��X�cQb���E�91so�ݝ�OI��V��L�s�k��j:���`  z�R���:^���Mm��ɣ�R?gLB�����u��ծ�@PD����+Kˢ�e��[���ԗ��q���xAAA��ϙ�%�`����]p� ���ls,��i�;��nm��?p��|v�lh#˵8-�s�۷/����N��j���l���+Z�*+ڨJ��z*�-d%f�eŵ���L�����\�~?/�_��s��]ɝ��i�ko��&Y   ���Ԍ��y���pl|�ӵ�	�YZhNs<Sl[+)�ϛ�_�����x��RW�Sj��a��`�^9C/f�e�R���>�����M!!!b�;w��bA7�Z��������d;����BE���  #���̺� ����.�$KO�$�,7Os�x�wݛ+^�|־����i��\��)T���>�wi�����>�r�غ9��o�^�_�/9[_��px��M�6Q�ڵ�ۃ�)S�����	ʗ��Z������ذa��Vz��aU��������G   �*�'0f�����e!A�\��wTP��L5�w?[�q��N$q������Fc�̼��s2w����֗-gQK���|�hWYy�c���+�,�N�����~��݋C��СC�ut�~���<�����=��kڤ��s���/  H�T���wλ�_A��?�c��	�KI��zܱ���k�|���S�OM��9U'���<�k�|?�O^��¸\%��2[�\�@_���߅�P͠��
�t�Rε��\s"I��nV�����  ��Ri�W����G����XLlR�c'.��t+]l��.����c�g��ܹ$�mwW��ڎ�'ܦ�䬽j�grR������f�e�ߧ.�WE��믿(--�Ԭ��m�t��x[,��аV��ݹ�������_��hu	  �+3�8#)2�����b��h�u�&�w���K%߆j���:�;9p!�/Zg�u<��s>�ݽ5O�{�RR�h	������<ůk����Y�;w���ѣ��Y��w烈~�|�����'��w]�m~�<\�?=}��_C�x�	���_��M��䔻t7#�   ������1��^���q�?_�4����$¤�9�1�3ű���I��_�y���[�4l�J�%E�=G����^*��ڷ�-�Xc肣*&&��͛GP1�����Ycϙ�������Y�[a��k4��T��˿�c	  @
s��/���?��?��ݳ:��\,|�=Y��^G�\��zg��ѣG}�A_�����zuk�������V2З|[�>]6��������T�Vde����n��f��=��SR״��a/OͻO��gn  �������y�MK�6}{w�s�a��de�ґW�k������+������S6o�-�a��5��7�m٬~m��x%�������}E��K_N)u�v�Ӹ�g��������y۶c���|���k��4��R����� �T��q��foZ���A�?��z�b��<G�6Һ�kc_O_���q���l���.��l�Gs3<�o���K��x�o��!�Nu��"�g��R��>ﺱG��m��`�b�2j���;t9�QO�hP���n���_P@{���   �Rn��Q�]�^?TH����FX���"M���lڵ�4��Q���V����VO�ZWn��]��vm��U�i���
rws~��_����Dy��e���n8a���S���ԯW���W������vw��i�>;{1u��c�J�(5|8Y�Z�q���z��^�5���t����   ��S����"ׇ�>�֒ϣD�G(�ẉ_j֤���qk���u�/K�g5Zܥ]��쬼t�\^`ooS�������^�}���ݧ *��C��|zj}o.լI�f�WW�k��|P�G2�����= {;g'{G�������i�w�Y  ��λڜ��3�Ec�N�#�\�Q�;ҒY�n�����]h��ri�w?�M�����:}L{Y��N�W�*�����b��'.g��z�&��C��u���5�,/�~�=���R   )���Ν[�q゠.��|%��C�W�m�=�y!�M�h����Z���:�w?��"�S�m�ة�Z\>ujM�ε8�Z�ZZZҫ��J�jբ�?��RRR*t��M�����8G^^U|M��;!��8�4�s��0�sq�  ��C�C?z�����x������j܈ѫE�Y�_ث�vSP@wj��F���3£��3ꢱxu9;XP��T�$����{�j�g̘A#F��T���̙3�C����IӦM3�;b����{��o]�Zd��zŠ�k�  ᡂ=�q:r}����o�x�Fʼ���g��7�Rߞ��k�G4nY_���A?�8F99�5�ZP(�ٟ�����zt�A��ݙ���vs��g���g����
�k�ڵԺuk1k���F�1U'E��ߨ�v�h��$�h�5��?u���<����  硃=<}cdxh�q�_\��Q�
E


Ţ�Sgch�S���#19���v��\K"s��/�i�ܢ��q�';�o��e�=�pe
I5ޱcGz��7��^�x1;v���۳g����裏(88�RSSi���T���� ~��4�o{���'�)�ߓt=�  Z��=K���z�&����>����\<��s�{�n�|��^�IH�-f�}�Q�~���Z�e�ă�KW��ɫt�R�d��P�z������E�h���D'��{ݧ>�.�;88�u+��K�СC�a�����YZ�jEAAA��o�p�u�V2'N�S�N��Y_ܵ�Ks�zR��~Լi=�ߵnMo���p9����L���_�haaA���:  ����~���y�k�W��q�uN��D�nݺ�q�F�2e
���z��Fl�x��������N�NT˥�X[�r���|J��%j�o�ݢ1)��-��J<�;~�x2f���8�>��I];ؓ�8x"�f,N&)�����T�N�znn./nW �����?N~~~4g��s��ݻ��]�6m(**�^|�E�tI���\O/66V�Pq�6�v%w7'rv�)���:|��͸O�R3(6.��ݸ�x�4%svvv�p�B�ӧ  ������{71r���A#��MLJ�NH��v�2���%[[��9�gCW�X!fD9�K�kk����KjlmmEiE�~��� $��T��.L��3<�Sk���ʦ)���%���f����nWh(,]���/_.����KF�=J�z�*Sσ��|����=_�"�_�� ^*����X�9x�   ��W�g#�f�Z:�����-��l	g�m߾}4v�X��O�O>��>}:5nܘBCCM�������ڸ[.��r��L�j���#�7�'ӧ3=�CK;2U'���;�(7�pkP8����K~^}j�+CXX%%%�k��%լYS�O?�����2E���_|!� ����҇~H   %��Y��i���t3����~��&�2���Q�h�ʕ◩*�K�_�>���[t���l�ޠA6l����-[D[Dc�p��$�t�'�oaz��̅z]��g��bHNN�2R����3y�k�v��A7o�!^����Y�8 ������wL������V�o�   ��$��d2yt��	mZ���ݣc�ݿ�l����x
��={�,s��###EI�����صk�N�����9fJ��C�[�ɴ\�[6�%Sq�j.��a2��2|x��������-ZD�Ν+���s�wr���1;}��|��{�f��������b��)̇J�g�&�2�xp�w��  PG�`��fn
6dP��1�IΗ�đ)�w����k�� �|||(""Bt�8r�����ӂ4w۶m#S�y��^��D��xR����/�ȥ��$������Iי�I�&ѣ�>J/��2���+:}�����>س��D3f�����8��k�v�#^+��~y�@]����t�};~�8  h"Y�g��N��)l��qcn]�l�����!�K8_�rE��l%��!�믿3j?��7S�NU�\�.�^;�N�"ܿ���z����?��J�]@S$Qz����ڼys�'���ʘ�pT� ��y�=a2�y`��@y�����dLx��������/��ݸq�   ��<%�;����'����lE4���N���Ѣv���q���������e˖z���R�Νi���j�q��J�9���Q��I�����ԨQ~���U����"���P����j��̗,YB			��{��siڪU�諯�2�NP��N�:�=ƃ^��3�   �1���˹�[4�j7�=���n��?���F���3ψ�1S�3����*���rtt,�1M�4)�<;���!�W���quS�i�&1�偹��rt-E�j?����;ȝ�   ta�`?w�����فݻ�=�����d�xF��}��ggԌٯ��JӦM�������.K�<yR�c�u�V�m��{S������4b��H\Sg(c�\�Γ
rSj1  U�`�s�"�<;����o޲��K&S�3ݼU��Xc��_�6��I�h��j����a�(;;��������]�,��@��ې���׹~�qM:/��ڷoO��g�g͚E?��  <,��D;�D��oL7䫏o�{����/[�ٽx�w�0e����EЋ��"0_<p�և���N����)�̳�%�m�V�G~Q7�2d�ظ�q-:?�Tݾ}�ƍ'�l�˘�$��bl�{ �t��H@�U��]���r�*,4�d@��%��v�ڕ����l,�7n�ڻwo�ʑ�9R�a��?�P���}��Q��<��V�ŃA�����S�����O�<�仱(���={������/ܵ��ի  PQ��;0+?�fM�����N��z�Lٮ]��@U� ��'x�Z�j� �}ܹW;���N�^^^�>����r�=��<���5�C>/W��o�k]6�2��  `�*%؏77;:�g��r,&6���s� S���Lo���h��]l�Ｆi ,]�T<��O?��ݻ��s�W p�ȷ�~%!   &��v�	�^̦��#ǌz��E�6Y����"��8|Ϝ9S��hZ��w�^�T%f��C�{�����nfƏ�3g��c�mj  ��J��sԘ���CgO?�CE����| �l۶M얬�E�'J���뼨�?�K�.bq-w�ᅦǏ{8   ���`φM�ް�C`@�aa� �"�𼘔_   �<Tz���d��Wҹ�#ͯ]��|��S     ���`φ>?5�ۍ���p|B�㕫�     W%��=7z�����'M;h��K"(==�     �b�,س��3"#ׇ>��X�ח�����B    ��W���y�ϙ"#��C=����     <�*��z�͏��лg�c7b�?y�     ��Ty�g��3���B�����̈́T�ĤT     �E�gc��Z�Τ�C>]�4���s     tc4�����Y����>=��?�\N     ��
������6�|���ݹ���G     �gt�> ��Mk���h\�-��_'     ���=5n��MBC���a��Դ�     �e�g���o�\?��qCf.�,����	     �3�`��]ɝ��Ͻ�sC{ش�7     ��:�ϝ;�p����>����$߿�!     (˨�==z�����<�����j܈I$     (��=<�TT���Ϗ��x�Fʼ�E     ���lĘ"��w<��_}G��ؽ
    @�d�=K���Z�Ʋ���v���     EL*�O�<9���?ի˱���:'O_"     0�`Ϟ�~B����F�ۙ��f���J     ՝�{62h�����O7x�e���K     ՙI{6<h�'�B;������~"9��   @5f��^&�ɣ�g�oӪq�^Ovh�g�q    ��L6س������B����#�q�N���    @ud����;�⦰���ܺpi��Nz&    T7&�٨��~�\���!��Y�"���    �:1�`�,�Ok�@���!O�ۼe/    T'f�
����x����ؤ����K     Յ�{6l��Ԉ��#G�/>!�66.�     ��
�,0x��Qa�oL��E䷻I^��    `��m�"��{6b��/�����I�t'     s'��a�?���    IEND�B`�PK
     �9s[F���9  �9  /   images/915d9337-ea3e-4fec-8caa-7acd53f715e1.png�PNG

   IHDR   d   �   ,�*�   	pHYs  \F  \F�CA  9�IDATx��]|TU�?o�d���B�RD�4�b�]�k]e-k�om����mVY]�  *-� Az��������̝�Lf�	�Ā{�Ef����#|2�z���ԡCkJo�r��m��N�N!����I���R|����ޛ��7��YCzS���;��|���'J�����H��A��xs���;���o0`����%�x� B�嬡�6)������������].�X,��jyr ����J�.ϫ� ��S{hm�����36�R�w<_��Qs�K̃|_����p2kS�9�;����P���t�O���;_=�w|�\�6��&O�L�ƍ���2�$�������^z��v{���^��5����������n�;�xI��a��z=������$�b�O�Bqqq���?��ٳ�X��ЫW/����C�ѱcǨ_�~<�v�"��ɟ�>�:u���r:~�8_��	�hC�n���?��7�ֵ]4i�훶���r���_~9�y�4m�cd�+Ծ]*��Vѡ����.��~��}�Y�o@D�Rt��í�[�A|�cD @+&r���9�DL�����ٓ'~РAt��AZ�jU��������g��ى	:t�P �%�=������qM�?v�Xߘ1cxq	����ڽ{7�o2��[�fQqqqDH�M���;a8��H���ת�l�&qLs�Υ��:��O�N�1Z���1��丵B�w]�|K�'�Φ!C�P�6mx�h?���6�L6�G�� d��W#���$ھ�N+�*�Sf;��̤_~��'?5550h 	/�������1���qg3�u�����ϧ+����Ow�_|AM&iժS������A�� �ĉ���@1w��ѣG�#A��w�LpF���������h��j�F&L`6a�Z�-���1��]F�c�]�d�k���ge��}	UUU5o(dDz�N��X�^r8�B���hp

�ɨPj���&/WRR�+,0XI���RjJ<�է,�d�h4�s�f����{y�Ϲ�.�@%���ԱcG3&�cbbx1��O8�� ,X@�&M���Fh}����WڡC�x���Ly�����W��ŋ馛nb�-&�|gi���^�^Wn4�j���bA �N��I�K���e�Q��x1�!P���h���L%x6^<)�9�]jˬ6�^��Iq��f���ur"�a��=�����g�M{�졽{������e�<P	۶m�a8."�5v�Yo:\pV,���CVV�s��&n!S6m�Gݻd�c6f*e���v'J�1��uE�~@��������j>����=y����c��-H�gӖ�YJ��;H�,��*&��/���A!�.�����w����y�6|�]w$��mN�ۿ�|������!X���[�x��������rZ�n�8W#�%�xy��_Q2��LYBU[-�Ҳz���z���Ç�̙3Y8l!11Q�}��:�Wt�`_���}�6l�C}����yU�>��fJII�X������v�Xqn 2�`��7�D���*mں�6�`���!Pw��AG����[wکow#O�Ɉ�}Ǵ�{Q���v��k�����E]��5Xؚ5kz~^^���S�~����a����o׎n��V<�Hۻ����s��)�� �`����+ڳ{��C� #��	�2q�Dz��H�+��P:���sS�\����3o
����g[�P���@��-��T@��X�{<
O8�Zi��W5��Z޷�~+�}�i��? ��|�7o_�\6J}���"!ན�)��+/� ���[����������9�5WЎ]���'=�����O�
��;/��b�����U�ӧ����L�7Y	l,���'��!y�z���Yh��ўR�b)w>}�駔��F��v�<�.��%��Ӓ��2&H�r������׵kWz��Q�i�C���b�ݞ�����oW�J��� �I�*���)Ե���v<����r�U	�y��䖖�ȑ#Y��z�[�n���}��K�ѥ��w�V��.+�^����s��zwHY!_�)�{CA*iY�?��{�b��d�J�b�F��]�θ�.��v�w۴f��TWc��I!� 1�؝&r��L�r�,�`wD1&���k�e�_)��_��pR�D6�k���\��!A%7�>����?��k[:4�[!�hU�G"��4�C��j����v�ø׿(a��x�'}ʵ�)~����=�~��B[�lawWþ}�B
a�x���8�no�G�/�N[������m�B&G�i$f]B�\�au���Ua �:L�!m
���	l�8��l��B�R�@)� �ڷo���J��$Rv��w6��o3bh�����.��MY�~7�K9��!$c �b:��:�oG?���JK+�t�� ��},t�Ff:�"׳�Y`t������A�n�'�A��Bp[b,4����kϑ��{o>ӨQ#��p��TA!^��J���U)}J@ȇ~(�?Q�Ν�&T��k�V�:�fv��?���Z��h{���w6����!PÜE�wt蘓��u0Ҁ0���j����e�~�K�/_N��Ӵl�2���է-9��,�S� �tIIq?��W��2"�"_���g����ǋU���`4�^�:���r��;�6�h�y�>��Z��=f�.c;$�$&�W:�3�G�	v��~`c�{��N$<���t�ȑ*���_{����ya�����O5O�˂��R�lx�
��PB��ܶ�*�V���qq4wI�����P����B��W<Tp8�֮][����z:��V��䙫&��y�
)2�R����Jۧ�@��돂@��CQ�ֽ���1���NA1fK� � �b���o� TK]YY=���U_�}~�%W?:����H��R�u�]ד����^�O���)��b�|��� ��$�ӯ���Ks�-�iO�[�`�W\p�C@ʤF!��CnMU/ ���bm(5���-�Z�r��'��]�4��gi�ܥ����m]��˓Ͻ䁓G��V�#P_5��?�)���^R<!'�����L�F�?|���[F�?�u���&���ϟ	�\�p�(T�o�2�����dI�9�uTt�E��Fκ�������~�uӘR�|���>����%o^9z�ݟh RpN�ЬV����5�BZ�%�Vo!<�N�q��V��B�	5\'J��������'{�ra�H�����0"��$��8��=6�͊3W�$�R�U~�P˗%)���w�`��yƕCG�1b�`�;d�������`��v�7�B�s\�+�N�#[ۈU�u_��͛ӚV�xS�)����-+�+��q�@�Eu��p�dP���X2�r�;�DN��<.;�����R�d��n��U��1���{����E���o�$R>�/�r��lY�]5���ˏ�V�F�|^����cȥ1P^�P��&�ٲ���8�*����ĳv��q����;w�{�$R������u霑#�1�޻��<>K�m�Gns�`W?����"E �ů�����p��ɨ����� �5�=N�;���V��Б�}��؞'�-���UGH��[�	�4�ӧ{reB�o��z \#�V�!dp���q5~d�B���@"��}�S�W$!��[FJT�yDb��+iH�1�@���yI/>�]XF��T�N���ֲ�����Lh\�B@�:� ����%�pu%�k�Sm�b.{9�1/S|XW]u�f!�!ZȐY-�2�4�:B�X$��?��C�#�����LD�
�ѿNʋ���m)�rXX|�A�d�a⑟E�+RI�yK�B47hq�Q�_����}�b�_=��)Ox��C�r����B�.�7'gU�G!`92�3�o���P� � @&l#4|* ����RyYQt��ONN�J#$HD �yW��C���`+��"���oC����(	� ))�	�C�D� ^֨�2F�����ZEj4*�E��b+�J�/|\@޺u��|T#���.�R��͑"Tf����I�8����%j��!��<HX �9^�m��4l�0Nj��SWf:<�����$�F$��HY�v��!�`�*�IG��W��`a�8���٣�����&eo�D볲��!D�Y�#s��-��09�f�d##/J���+V��B���??@}�S��������(;;;0�`��������'��(����z�,�Id���E��V)���V^FW^z)y�8�ʲ��v�y��F=�p|��
+erK�,��wL���R���; ��(�jR��#�֬Y<ѐo�_=˴p���K.���Xdi�GL���|_�,�(:�_Sb~�RL�Y����!�._ٌ`1HxC-7 �L����8��*B�{Af�� �{}��G<q'S���aL�g&��{�;V+��X��,2�J!���S�$��jYxQ\��]�mۖ�/�*y��z�#E�0L�"'�VncTe�\P
X�,����������)�v&���Цd�	 2��,���z�|�0��� *I�s�	��q/����V͛YU���C��F�jY����{�Z׃l��`Y���"y=V6���#b*	85
�AD���4pȆ\���L�� (L�����_��A:�����U
��!�!�0�ËJ5���c��Q��$9|��!��o7�t3�2z�����`�P�Q�d�J��P);�8~ٺ�>��	��R
j'�J�]���Æsi_EE99��Z�tOQAz�8�3ʧ?�#f �gZ2���܊8�C����r@^>�j]�8߁�t��y!�G	���3g��5�Nz�C�\��^��T%"Ҥn�z$V�y�'�9�脄�})�¦g�6P&khN���n̪�ލF\��zi���XP�F�p����M��ә}Mt��XBfV6:@`K��4sn)uH7����9�W��{��{h��et�@3]61�wNE����<Θ]Bǋ�ܔ ����Ȃ�(
��>��lNV@ +�	5]� �p���B��҅�
�&j"
e��f�7�hM��������U�0syB�t}��uN�pFO�k�����ZT�c7�L3��j���z&}5�:Z�j�g
H]�� �WYe�7�y�Λ0��R�XA(�������s�1�r

�)-=�������X���dUV�x�O�ts�5&|�����8>|��'Z^(�U|K���b��*����k8~�g#4�j��ۑ�'x��:?�����	�ӊ�q@+��,�Z�|<��f"�+�L�B�5U]*�W�c��)�`�q�59H]/ʈ��9�c�1����$�ǰ�c�s�$�1j~���pWX��/�Et�/��&}Y�A�*R���8$�ͽd=�Y��	�U �+��G���B��h�7�å��؇�@-#��E2�������װ�e��B��ؐQs����Q9�K�:n�d+�������8�4Ν�f
�����!�Y+�z����4JPCᦁ����{F�OR�p�x
��-��(�3���P�wt����b�}\��P��ֈ�z�h���P��?!�<Y���d��t������n��Z�u4<7n��_�-
�d�(e�G?�D[E[G�T�:�kuu�����-LɊ wJ�y��4fM�L8<]�0@��j|�`�r�5d2ǒUhX�.~wE���o�˾.��gE�e�d@���"���[(&��ý��	�~���|�dw8�cy\��&�-dbUe%�Ξ={��dj^�	�W���US�2�w�-�;�|Me��{�.���Cj�P�a�z+B�f�?��%����X,p�~q1�s�I-�;y������g�+.��bcL4��+h����RaTe�2[k�i�$�c#%�����x��-Y��d������ǡB�ڻ	�"d�~�#�e�ތ�8C��9�kD2�������8ʉ�~Z�gР���jel������'�"���ӛ�Bj�^L�SiO���ș��x�R�s�.�O����2����tP{��׋%�@��B�<��A�u��䊿C��%�x�ۙ��rbB�}r�9���_�뀌O?�4p�ψh��6��D��jס#ev�R��ɥH.��l�ѓE��l�������1�M��)VwT�~��h�������Ψ���=!t:a'����S���-_�o}�7r&L��Ƞ�;��.�&��X|�@��,���ԘEX�U�����
��z<r�	/�KY>���dS�o��715�%����:��`Ih������8�ٳC�QQأ+c�tL��:���$adpFC��&��1��St�� |�h��I)�Z!5�ז���78 �#�����dpL~�5	u�LAT�DU�DlFQjPz��	�~e%͚_JW_�N����do�a�?�=�.K�\�hA�;Ĉ'��렇_8N�]OS.M�u}�n;M}*�F6�]Hb^�qq�>+=��	�h�6`�,�/�lvG����q�BV��m4�@f���"�lay+C=zq�����
>���?��M��gҼE%�Z`��>�9.�/��_\A߯����&V;/��,Q����ŉr�5�!@��M�3k�����9�qLa����?�f��u�ӻ�޽�z$&Pv�&�5u�ؙ������C�z�����z@yEm��WoBM�!�C��Gi�ZQ��N
e��B,��hY��KC���8��A�sZ��cƌ����yw���[�F����4#��{��n��o���ڐ���Fx�����ģ-, y�HF �"�9J���K��pU�2��A��Y� �d4J�M4��ǰ�Offf����X&^`�JX�' /@�X��'����
[�Ȟ&��n跈|_4WFb@�������~,P$r�1��%r��J`쬀s�%Ly�E
͊��:�J� �i�E���F�λ�%bQ qBv ��C����u�V�i�R^���<l�g���lv
	œ%b��5�ѥK����y����mi��6�������l���o֛@6� ��uz�?��kI5
%f�.�CI�W׽�4\3|�(�C6E}a0`U�Ș1cO:��1�sƌ�Bl��w�#��������t��W��7��~�p�hq>z��ݛ|����$%NCZ��<��]��J�.�D=z���>������ɾ,^/���}D@X؂�B)�z �j(Vw����l�}�Nyx.jAP��FF��Ub�i���E �+�+�@��#�~�=����D���?Ε_X��H2�I��IoO�N��J�NZ�����x��:PN��]<�"n� os8�u��C�
]V�\x &���SO=��!��ܖ�q�d��� )V�>���wЉt|}���q�*J��AP�S�?O�۴�cyy�C&|z�v��n��.�!�(���"֮�jP�-��JIl�D��G�YG�?	��顸X�M���o��nddoڴ)$RŲ�A`�����%B�K�O�Ǟ��9l�e�-6�g6�-��Wd��I&��?�HXø|�1.U�-�1FP���U'
���R�x'l E M��f3���0r9:e��X#CՃ����Ř�PR�Z���|�d��P�h�.����W�EY`k}ړVS��%G�*��d�-��}0��ΑBn��|{Ne
!������Lv��k�L���/�mGF?4/i?!�j����)~x��x]Md�I�h�
��ӱy!BCk�`E&jZV��x��B�~��A+^�H4ǘ#ҪԈ	~F]Ȕa[���KSyY�
�F���PQ%~k#&��0P�	`��M +��{���$��E�8�@�0�v� �f-�|Z���}������˃a�����3f��%�J��T����Y�1I�����Z�);%�%ԥsV!!�Bir�=!�T5!˸{�9�%�ɖ�V$���xj#Q֪p%�X��c�v]�K�9�^Cv���;�!*1u���LՐI�l���A��U�[Bjr�#��7��bk�:UV�28������IF�@a����3;�ז��.�{��s�$�͋M�AƉ���wԹ�܌���E��e�H@<�-X��� yMz����zW����]�ԉ����ߺ41�D�[y�F�eW^I'��+:X��m�5�����Pi��
b ���5+B{+q0���3Iq�&��.s	�؆�d�	�0�#C	��Zv^��� �wNj��d	4Մ�����f��'�uA�C�EM��_Y�F�G|`S?�
@�)�п_�ڶ�Z��"�)�5�k�)�n*�QD�t�,J$T�b��gY����;f�_���oǱ����ۯ/���ճ�ԪWUV5Y'kL.�9c���:_{�%�#xR%k����W_���n�HP�Z��3��B�/�>AI�P��3
�Z~6�6�;Kȶ��.��zZ�pA�qG!b����Rz���ŋ�;(��J|ը>�t9��M�:ұ3Ti�B�zJ�"�ǎ�1b��@t��M-��k�%�d�ʀ,X�?����j���W�8n��F���,:��%�M%C���d���!(��<yN���h���\�����Ι=��c��Y�XI��=���W��+2>!��}Y�t���;X��U���-����}�tr����\V��@ T���t�M�.keoȦbw�8���7x�Գkws�9��P�k��F;�>T��Uj%r�ei2��M	���Y�/�����NB�`�^�� ���,ul��z���\8\"-��	,�)¨t���Bn�Xbد��*X���ȢO{ �չ�x9�&�B��^Mâq���ip�e���pxq�@Y�.A.$�\z�̢^|�E����tP
�G0<�.��@uP,pLvC��<�lAM!��]��"X�R]�D�7�/��#�
W��7Ae����4֍������r���S�2�G�	��'�,pb��EA�������G��r!5d'�F�e)�@M!��" � �#l��Mk��A��}�Tf/�s��4!X��޷҂n���U�{͙3�����?ƈP4؊l/	���|��qG��I�` �9��eoΦ�}���P�c=2� ��a 8#Q{r�� ��)`>`#��Q�eed����L�U�/7W���M(���yMG�^���>�h*�Vj���;�d�/��a��.�A�>�� ��A;�z< <�!Էc�O�T��p���ǆ#P��D���@~��7�	Ra���単	��'�;�]-41�������&�AT|Y.��*���$���õ|Yj�)�!�%ży}}���&�e�����駟x ��;�C���?�˟����>V��T\\Q�<: ��+�g �< _�NE
Q�e	��d��g��}Y���p��8�!5)n�$d*Tl�!�ٛiܸ��WJ��(�N*)-�ٟ/fѰ�v��$ �
����/I�tU�^��λ֫n��~�;��?����J�D\���YM	?�9d��۠U�i#���2�"�z^�zP�}��.$?4�dٲ����8�;��޿&@m���!�w	�v7
!��PS�� P�㪮R4�T�IJNb�����!�Ы�ɭ�ɔ�f���]h�/>�#�Ӏ�����L*Cj����h��m!��-g[�Y�D�SF�j,4ڗ%�&�2)@�t8�T^Q�Ã�r8SSG�Tf��ہ�u����`cN�� & ���o`�6�I�K|��䲁��<@]N��&T47�����B���+�����;����#@�Ipn,�@�M�{��c�@�A��B��`��T4p�(w 2#x�F�,��Y��sG��7�歿В%��:O]���}.'�4H��Klٺ����|
.��l2 ��f�DJ�}X�ֳ�AA�}Y`W�**=�IX�*�?6G:8B��,K�x��'Z����w�dܷ�=ڑ/�T$�H���?E_�lBXGF���I�va�\�*@�M�UQ����Yh(����@��a�3�(�u7_���[˿�����ܽ,�;v��	l��l��wbC!�������ڮ��V�{���K��man@�������lm�U��r���Z�!Q$��(<�joz�t� ���D:����pђ�7�OQdԮ�/��B���2|��b�ڬ�4Ҩԇ������[���&΁f���
Ë�,���E��F
2�����p��W���e�7<؏
���ܨ{Q4���@��P*Ԋ�Lܖ�79p�@���T�uP+I��e94�H����c2K ܣ�pd�c!�lx�;����4J`#2T�a�H9N�lB0�؛v��e2/K��~�jo`���&�a�{ե�+ j,����{6@RF�be���w���4B0AH^X�pa��`��*Wg�KA'��Ϫ�����<TC��E�Et�o������yY�����"�V�(2r�M����Y$�H�'�t`�NZ�[><4q�0Ҭ<�d_�%�7c�ԣ{F�իX��2ޢ�c~��0'r�6���!����o/�����Zu
���Pk��oO �Iŷ!����TC�
͂�f�����k!����\;�<�Z�{�N�dS��_�J�Ӝ�*�kS�	.���T�қ�� !�bb`�A��U���|�h��15����/�B���X�|t�
l�d�anRPX�N���3�?#�=�O��n4Y"���n�އ�#)�,� ��i�2�f�#�Mф4{{&5D��O�3�f��t����N�+0�p!�PI�jc�I��[��@��V'��&�В"��P�������b���
f��?�
pZ!DB}�-N;�H��}���$8�"�#���I�&E={>҈��B� �>��r�)�	��P��*��!���\ ��T0�,�7�M��x�Av��wA�G��Pz��Qj&cu5�i(HgjEyw#B�+)^�޲�-����e�eL�M��L���k΍���֊7/V�Q 鳥e�׷
�d��>X&�~Ԏ��x4�D�i��kD�6l������ J7	�|US�U�.�69B��w��:t0r�TWV����%���Oe�1���ۤ�v��C��,���D Bx�v8d�����[���#����ǡI"�� �c��̶⡂59=�E�E���S+oԐ���l/';`�pC���v|-�'W~(6�ܧ��v6�߮mF��G�Hb�H��u�Sד��.&��A�R[�q��wxF���A��سn�:j鹸�>�('��UA�ο���<�>q��g]��@@9<Z�x5�}��Չ �XP���!Э�%g6ԉ�w�5��{�5�8~8��ݩ���VO�/����aW5��<zY�?���s2�Ɛ�J�Y��������袋�qC����C]#"��9�����4jD��3��wK�.*,*k_�)��]I��.��T��c*��rZ���N��M���^�H��+EN�"�4�E��#A�_�rd +1!��"�@�=���F�@�zf�^�4k��%��K"�BH��j�2�,�?Fn$����
Z���Lz>��PZ �mD2^�'Z�����O6E�Cu4Q�YH�H�J�j!d�@Ɵ�}��=�z���d�E���B��R�7�V����.B����K#��;\�Ѵ�a����TR�� `r��2��������Yp�B�y�Q�c�K4��3��z/^�nщ �46�,4)G``��9q/�n�s��i��JV��J�����/�<��wY�UR\«_�\n���+������LFŗ�(=�����#t�ԗi��3�W��}2�h e ��&�L��c��h�b�B�2-�'(1Y ʤPr|5����w�ۛ���Hp����}�� �׷�}m#��s}�Y��!�E?v#cɲ��N��;���Vׂ�
�-�]ag�%g�hr��"c|��xٿ	�:m���X`R&E��:C��"ɢe���?V�tF�C���Oj�o���2Ae��:���s,"��l�ᾺXy`/�PO�ْM�%,\�%-5P%����DJ.W2���c����/2J���|ֵ��i��G�X�z65Z�!�Nv��ZG{=xP��B�ʓ�E���h�"f!�
\K� ��aWo좐�G�q�����M����`�"A�sj�k�����D㲒	��Ѐ/���M�:�8�ju@c���+�	5��X��\�MFK��g����u�q��������*Xu�7;x� ;���&�J�ݹ�4���h��/�}�� T޷�Ӫ�V2�t��{�rkV�lT�#��-\+�n��Fe]���ء3ڠ[��/��(m���S}����5�����{o�>㭷���u)ر!5UC��]�9�	d�ꩧ�V:*,v1k¶@6c+;u�{P�a�4��/���r$p̘1��o�-UV4tV�=98�VR���C�#Jְ�qFz2��UQޱ"�۷#�'�`ׇ�l<a�L�,�bL�څN%�+�T�*4jH�=�L_~_���!䊲����������{�9ڽ{��I���:�WD�Uv��_�BR4�T��8�A0ţ�(�	V�+���^���}��.��\3��*5~�����ݲ-��Vl����}n_3_\�C��.��&Q���Lz��e�uu[PV<��N����77��1�t޸�'�F���'����t�/�K/��Eˉ�B&+�Ġ+�ĉy�d��Q��R���5��UV���w��}q�*���x<N���'�9�*��2������X�2P�����e_ 7%9�ƍ�[.(����F���ȸ���ۺ�4���t���h@�(��#�<«�"ؕ��l�:�$x��b�Q���lJk��l�+ɢ�$ߦ>�F�e� %q����(�^��=L&�`����*��*�����ٱ�o���j�!r��^x!���F�9� ����%�Ř�Q����_��� ?�b��?��%����d>ߏN��>� D�hQ�ۏz,8��x)��w���~��-q8]`<����@X�PzI1a���?�l�ݳ[��E�b�6JJJ��`7 ̍���~UFݖ��C�F��0��5�VZ���iBj�����fzl�8��U��_rmjrܵ;v��Y�yN����a"[?`�����ӆ�}\���OO>�o�k;���I�4���.���χ��gѡ<'Y�r�*R��I
u���|��/�~kr��Q��~����tѰ �ZN2kN5ɳ5~da"��n�*�&����+A��ݙB�=�/�b�Ç12��3|�p�ī��g�c~��O'�);�/�ͣ�ؼy�]�4�l�FE%��'7�)+��`7��rR'�!n�Pu]B�茌���MtV3�;d�40�u���\�"��@�%L�6��X]:�Sr���:A�	�ش{�����B-�`�����kX��֭��]��u׌�LL�|�ry�.�)��7�ֱ�_Ε����!PmK����iE1�Uoq��K�(08��'� ���H�q �d�8QH�?����W��攔VM������ul��N�]��G���Q�t�R�l��⨳zQ�Ԅ��������~��]ɾ�VU��z]�1�!��C����/>;�,�	�H�lֺ:��oJM��g�(�j5�j��ܴ�����5}�b:Us��]�V/��U>�P�&�j;�����MP`����S(&ǦӆJH�Vk�B�5;?'W�Ai�Փ��&r	rrð�� |IuZ���r�u�%�X����tSy�~r�Y���;2�Wl�M�Y�R���
#�����k6��8VP�//P%{ 7�c8g�#�y意Kț���@u*���P�4�wr�J6��|q��*��dm�Cw�i�T�����t��qw������~��12��w��4c�L*��j׳[�'
�iݦ=,�� �9�x�/����GZQJ�Vh]~1��쐯����5U���"^�A��;�H.�1<��'�~���q�)q�v�>J{���ԩ��9��-��ߚ[>fԀ)�������<Q� g���t��wӋ/����&�x�n�W0�Ҡ��Z��J�>v����~�u�F���ak�wL6�Y�hMj�?B����вe����fZ�3��U�4V�g̘qZe;ꮽj]�t栾9g��|ۺ�;�X��@.�����*��cp���O,�m��e��VkX�`[`k0A��ݜ�R�,�5 9V�]`8��O���� M;���2w���n߹�'X�L}�}�8% !����x��ѻV�+T��G _k�`D�>�7������o��������ǆ>�����.�'I7J�!ҍ�}�T��,�ؕ�,ʢ�\B7����ߞ�ŏ��E=NGղ%�/��F���}<�z㭹t,����=nۘ�k���4!7��M
�UR���FG���    IEND�B`�PK
     �9s[z|S�wq wq /   images/b949fd05-6e10-4256-9d1b-e11f1f9900de.png�PNG

   IHDR  	�  �   �]A�   	pHYs  \F  \F�CA  ��IDATx���`[�������cK��{oH�0�����y��$6��6��EK���i���Reo({�Bd�v����{�Md��I�XwH�~@�$�W��{u|��O�$	�E�?�t�:R��t��p��bHCI�             a�!r[��sq�`<%+w���D�])�Z���y���MUw            H`J)1����}�`<!0%�<��ϕ�)            ���3�}pUp��^���1��/             ��xE��ɞ2�����U"-            �1 ����y�ܟȪx�u�             ͳ?ܗ�oϜ�A�#�Gu�zFyi�fc�Ի            @�(���@N��}���[�O./�x�lC&            �(#�/��1��ʇ�ƃP            `�}�`a6?1�\+            p��#��Cz5����k
u�����l�����7�0��~u�X��* �G�ϖU��B�/���ZN�98,�t��            �k`��r��Mz����+!�6�WZUS���}�R��ܤ�t
f���F�ߧ䃵�	�9�p_,#��*�ϟ�D�	            <�&���Zw�Ǆ�o��+���{�лf��&��c��h�.X.���s����{�2��fO��)��x�%;K:[X!�>\"O/Z}�G�U�`�@����F�           ��T��ʍ��zT?���T�^�Q��].�G�|�=)��>��]q� �kIe�<�t�D��'����[�@�}�:��D2�GG�tX_����(�}��`ld(��{��            ~��t�/#%Y.�[�-Xq�ǟԳ��m�Һ����RQS���������EC{�i}��{k6�Q��b�>�&+w�yJ�P           @�x�����B�d���'<b���Q�Gs�	�z	���ġG�i��b	�>��g�o4�           @����E��㎓���H��A�zwQ��MKN�K�����ٹWl(��z$�}�}2R�#�+���&�Bb\,            �$���ʳdP�6�2#U��Wʊ����W���_K�0���^��
��1��<~������>�a}$��b]��eQ]����!�B �nW�Q<�p_, �[�$���J            xRj�_�5��v��Aٵ�uߢM;�G^��{��ٯ��św�q]���O(x�Si,����j�a��Q]���2ک�@doy�Q��>�#�[(%g            <���V���kY�}�lܻ/�7�s;�|D?i�"]Ftm'����rf�d{Iy��xt�r+�׽U@N��E>X������̒q}�X��X��!�c�E�w��O��]:ggEq�����`�2B            �9�~�\f��@ʪj�?o�
��k�߯�`�Ⱥdg��.9U��߯5��'�X%��h��%�����]u� ��zM����W���?��ē'pI��}�>�"�[(Q            ��nW�!�W\Y-���%y��+dh��r��r���ˎFF�+�����Z'�=��\<�����uaA�����ix�Ͼ���W��"�}��[�O���}            �-U�!�������Z#�س���tm��գ��`_��d�dXk�?����W�l��_���PX�e����`�.�*�)5�T ����l�W�a�2��R��U|�R��C�r#�g~Q�J��qYKeH7�g��?�߼o�y_k         ptc��Zm(c�2��E��D���b#$�a�$��h��F�|\�y�g����?�O)�!��`w��Y-��w�l�-�%��ל0�.�w���u������uJ~��ɯ*�9�!���!�|��a�,  ����<���;�zgϬ�-�Y^��3�|����3Dg�'         Аa�6D�Qo�E�S:s��c^�ԩIYe٣T�7^����8�\n���Eʷُ���C>.l��r�٣��^��G�l/.�K�������YY/$�S�C����}�"؇�3T�O$$  {�'J�%��HѦN�ȓWD��ݛ�����/sd�?ҲK��6��:�Y/5��Hm         �U"�1�e�}^�M���b�M�-�X�]~������K��%g�Q�����Rw}����>v��+�γF[kz�����E���b}���1F���x0���ʴ��!� @�0D6��gH�߷ϸ���'�vSe�ȋ�[M�ѹ���C�j��          q�2�#���Y�{�~�������/}�ʙ�OI�.��P�"钝%?>u�u���F>�f�a���"�p�f9�w��	e�}A@=��ӋVb��`  g����ř{џ�)qa�O񛛙3��~I�lj2?         Ĺ�"�Ҥ��3x�%3'�T�Z�L���;�@���5���?�����/eٶ]}��~�$�{�eF�u���K�a����g˭`_�V뢽�t�WFg`C��iy]E�  �2j̃���V&�|���J�Jgޡ���i}眹��н���         �!a�G�)�)%�N�]$��;�M�۳�̛��9��s�uY)~���IC�KAq���Uh��R��ҿ}+�̬{��u��o|֤�>�t��w��uS�jL�"����Ϙ�W�c� �A�y�l����7e�x���&n5�\��;�?��U)�E         �g��n.�/���&�1���#�je�|�z��]ƶ�Rk�����!�ºhWi�<���{{�T�BMZ��v��%��1C�����6�Rʐ?s���9�  ��T��9ť�w��ֈǕ̸�嬟�9NՄ�e�<_b����Y��s=������7%Z�g���q��g�zW�}�d�Ϛ���d�:�z�C��K���k�����/�%Z�g�Ȩ��?'Z�N��=E{��I{e��h�7��+�<���Τ���굅a<0B�n�/�B<�x��y�����֘��w4?�h�9��K�V�߮�����ooy�|�u����RU۴@_}?a��z{�u���Z�~"^0r��� ���۫�gN~Cb�~�<��0�;�.��o�#:���ߢt��]�^���׼�W��O��w%Z���\��-��M���d��"l_�Q�}��y��^�g����O���jd�◚�'�Y�e���z����Y{$���D����5/�K�߰R�d䥒(|�_�B���h��D����>^8�H�z���h��R{e���x����a)C��h�䧽0�nS����2u��`i�_�U�T��v4?�qO�u��Ҫj�*-�A_�!A�v'��}�_�Y>_�߫�5��Ba�[ur���T�<P��J���JF�s�>  <�<Y�`��s�:��)�h��!����aCS����yf�?;bi]��z���7�o�ߚ_/�     	�0
�ϘP4}�b�EӦ��ܝ����'��ET�۫����ky���Z9�4h>��?��P��B��{���@�  �"˒��y{�8y�ĸ�铞Ϟ�?!���RA         <�0�����7�H�+�1鑬���J��(��p�dx����17��'���C�  �,U)ɧ���{%NΚ�^`�_�m�h.K          �1dM�/����n+�8Q2s�K�S��7�xM�J�VJ)C��ͫ*�1���#� �{�׆C��;)nB}�y?NɿD��y@�*         �G��U)߹���'�����Ϳ�0�Q�`3e����@n^*#�E/`  �`;#tny^�6�SE�&�șu�5o�         �*C���	��o�Z�T�I/s�dV��UM [1r�]� �4C���]S<}�Z�s�3���<�j��\          W�O��O^*q�h���y�̫�#�ق`  3�L+�~��� �2��2P��$��x         \bjfьI�K�(*I�fU�Q'
`;��s�yB�/:� � C���=��D2mZ8iʌ�Cʿ�<�k+         �����4�nI$�Zcܑ����J�� �cZ�h"� �C�

ݢ�n�`���ݒ=e��O=��:�!�pH����[�a����m���m���?~�_�,���A��R[[�ט���)��<��-�n�����S��y��[��y��[�]oTR�3|7렛$����r��1���0���Q9W`Zި!� �c���r�K�*�5��@���c���x�p8,���RQQ!^ԡCGk�e_�f���E�T�>j׮�u2-��?�7�t�^ܾ>�Oڶm��m�0�g�^5_��W^�����L���/*((�ޛ�B�^��&���;�mѢ�u�"�m�`�U�Q���Kh��G�?{
�6����h�=ƌ��&~)	�8s��`i���=h�xHJJ��~Zuu�x�ޗ�ٶx�^���-2��4���}H8�I~�0�W��{m�z��=�O�h�㺴;��=e����r��ee�ɽ:7�o閝�~W�1/sd��ҭUఏ������j)�����*�ZX*�Q�dŠ���_�VQY���r�p������$����{k6����C>~L���1��������$|��f��w�N��.k��ٴ�D����r�$4e�U�İ��r�$))Y���S�}H۾}sݒ�z��!����υ:v�d�[UUUԖ��z��ա����o��ٟ�r��}u��޾Z"m_͋�j���(�3�U����`��TV�;w�Zg����!״���.7����:�ؾёh�F·eN�z��J4��Ϟ@{��Ϟ@��QI{�	^=�0D6�V&�Fٴiac�(_�����yF�.]d��͞{�Jӗ��D�]���y�^�+++�b�O#��\��p��R��Mh�{7?�_yrѪcZ�/'�$�9��A�/�P g�yB�խ���3G5�k���r�˼y�0��	��gjBaYQ�[�l�!7n�ז-�e���W� ��8^�A��.Y��D�_��d����>k����C����F�EC{t�{]_���ǧ'����2C�|� ��'SeΤ襘b����
��?�Dnrk�.�t�'''�6zξpA�gꍄd��0E�^��o"���ؾ��g�ot$y,���o����st%%X{�5^�̉tj�%���Z��7���b�.�u���&�J�7\��7�*ٟ]E��UI{�*/o(C~�s�m�����&~��ڼz�x���nz���2�v�ջ/�g�}�A���у�)ؗ��*��-���)��� �y�{J��t�U�\�X��'�:��.׍l�D������¨��/~v�yf񚨍t�f늳�>%��'�5'כq~�V�����y�^;C}^S8[or����ؾv�T#�h����3�=�����t�8թ�h���+�g$���B����Q������^%�Dk��xCc�:�z�A{��+�У�g������귆/�=�Αx�W�nv��"�S�����}�*�����>]�kˬ����{#�KZR��)��u;h�W-���������->��=g`�G���;�����7�DO�|É��o.$:�;�6�V`)�>i]07_�ts=���+��N�
"�S�S�{a
����޾N�dh���h�l��uN"��"���q�S�z��t�nw�Q����Y�W�&�gg�^٫��IG�?ۋ��,�o�iӼ1,�κ}I0'�Qr�x��a7�B}���D�/�p߱H�ww��*kCRm^i)VXMOQ��7>;�e\3jP��%��.+:�׎\w=6�Q���y��7(j����˹��O�?#%Y����'t�`^�˙��KZræ��a}d���K�V��,<��f�j�y��cZ�ڰ��������R^]#HT�΢��|
� �3�(W�}���n�
"�S(�3�m�R�l_��[���L;9�ف؟�G{��+���^y�[�9nuj�5���j��}�ꬣ^gP�3h�`�gg�^9��Ig�?;����o"�-2�*4����?��in�ݜ�E�[�S����!�̮,�y�?G�;�Hx�P�
��x�붞���7?3O\���:��]���~�U��F4{�Ze��y�z��~w�F�����{Y�wlc=�M;��\:�XXQu�����E��p}�vs�z�`��rƟ Yi)u�풝%/��;rz��V��hT��cUEM���?��ʐ�;Nf��@��y�O�x�����e�l��^'�n�
"�S���`��G�?;���>l_��^�����8�9�v��ӝ9n��������733S�P��uT항

�9���^�W��J��Ys*�U��u핽
b�xC�<�mڭ�^I͘�^ '�k�TO�(��nn��"�^%>s
L��Z<����E�0�[��.ا�O۫��_��I?{m������˛�6D%�w����Zoz�'�Xe��	�iz��h��ƞ�J������ҵ���dh��u��̔�W�-�{�yId�_"Oi� ��n^��GK�*����Կ�3�y����N�)�*�p"\�P�7���k؟����ګ�S��ɩ��tjP�=���S�����p_���k��B}n�b���#��u*�W��u�ڣ F�7|���P*o�y���aN����P_�S��b�G)��%0e��;<�}���d�νҷmK����6)ا�Ž|䀺�O~�Rj�F0�O�[VU#/~�NjCa+X�G�Ӿ7�����ֈ{N[��P.��3���WJ���u��5��5��k˿�D��`�5r����7�tƓ�8^��� �(�1i��Q>���!���n�:L�Gq���'�ۥKWOu��pA(Tf[��;w�X��n_�՛h���z��tr�ϴW��δW�Gwn�6�HJJ��ƨW�]��׌�Nw� ]�޽{m�X�b�EEEV��^�Wwjlٲ%��gګ�I�����n�y���z��k������,����^EO2�'����ޙ�>�,8X�g<�+O�4�~��իm��ljjJ] �:w�,k׮��|A��v�7y����wn0gv���>`����_��u��a}���ޓ���'���S�f���~�\F�z������dH�6u�_�j�5Z�����r��a����T�phoyʼ�z����|�{�r��#�%r�O����w��W�{������K����9��&��5�!θmC 7���صk��޽ۖe�`���ٳGv��i˲;u�,^�����v`����z��}i��ǋ��^E���+V��e��`0(^�ے�˗۲l�֛H�W��vm����Kvv�x����l�2[�=p�@	�%�W�3��
��׮�j�G������l_��L����*:���"%�U=2��Q%�MY��_o^�%W\\,k֬�e������z3)�M�@���:�g�������z�iy�����B��q���[�R~~�I��)�HI�K���G>;���u����WO���`�������k�-W���n�/\Q���t�n���;�Z��]=j`�}'��,�[dÞbIT��.��?�J~p�m���$w�5Zr�yG�81���~G�3�>         �%t����T�<�C�#�wX������{k7��~ݬ�׌t�`_��k�و�>��'<Ғ����n���7�+b���j��߾�u���]�k�,ٴ�D��7�ig�!~�T��7X�K�Ӯ3X������"A0�6�F�/8<}Re�D         ���pHj�޾~��6�}�D��GO�	��أ��k����1W?@�|��Y������5�!��eFZ����P����/\)S�O�SJ�>a�����-_m�)�J+LC||����G��t(�,�)�O�n�iy�>�D�e���|�~�gΤ����BUj�?E         �(1V�μc������*Y O ��(�}@=/~�N�+�%��/e��ʴWO�]=���r_[���.���:\s�4��z��ݳ��Ⱥ�����6N\��w��m2a���i�R ���B�餡���j�֣1���m�82�)eDg�8W:g��`N�n��Z         �f2DV
�h���́��R%*S / �w�}@=�5�����r�C��:����>>hļ�u������Ei�N�L9�O׺�+v˗[w�8=m�������vo�Szw��n�8�l�i�TW��g}9}�7�Y�P�
+�d�;��FX�ń�䪇^�7ÐU�&Rz�ӓ         h&%��5�2��_m��F
���}ٹyF��K�#���W��:ZXS�rC��\So��%��֪��?V׍T7
��.�A���`_d���� [}�2��ws?X,7�&��>�pޠ�2�wg�p�AS�04�!�Z�        @(��L)��])�}�%>�Pe��I�������m�f�^�*�kGn�KKN��׷��_���P���k\X#F�C�����/~�NJ*�%k�����#w=��5�����S��ܚ�K�H�3��\�����~~�r�ܧ��'�VA�(16Y��         ���&A��6�KO"�g!�4�+�Nգ������WZ�/��
�E<� :�����Ez��ݞ�n�l-*=��+jj���k����FLON���'���+qCJ������P�C}+
v�W|sL�[n�b�ß,���:�n�ܫ��=��A�A"~��D�T��         ���{j*C��E��`�=���;ɚ75�/���/��_b}/��m�a�Ң��r��90�����?���u+���w#AȦX�y����%�U�B���?���N�}��`���j�5:#�a�r��D���         �Z�T�$���t�W��<�G�hĶ�Ryo�&߯�u[�t��k�,קK���<:����t�T�z4>=��|�~�l�S,�[��'t� :���Q
�V��E�/Q評'�~���ں=�c�tx_yf�jA�	�����0����        ��RR�Y��|������8�G�8�y����un+C;����������E���\�=��5�n��K�6�M�ُ�o��i׎(��8_�6�s������#�����屛.�����(/,]+�� �)I7�R��          g����5�} D^�r�UTI0=պ���=g`��￺�룚n�p��wl����䫎iYW?P���Ԅ��e�$���mܷt�N��^]�^>�f����Ѻ��z���w�P�}�BU���QF�        @4TW��M_���x�"�BemH�]�Fn<q�u�N*�~_���5����)t��mf��3����Ց����$���}z$A4��^�H^��w�n�u�hy|�J�������k"eH�\         �����k"% �E�8�yV�����4�o����f� �6=�������lp���Z�[�Yи�m����t�nw
f��c�ɜw���8ah2�	         �C��8�̠O�0�}�a|�a��ٹW��m���'�X)���Ou�ÂW?��a�|���ewY�Q-��S��-�IVZ�u��=�}V�@��M'�a��6�o��+}�~���rf����R6e�	�0��ƕpH���l�:3`         �n�&Qbt��<�`p�-X!�<���=� :��=����ʨ��`�6ykձ��G�ꄁ�u=-�ζy��{u�?\zZ��*jj%�F�;�%[v�sK��e��Z�[e��m�������&Q����         �#�O�$���+�� �"����3K���6C6�)�ʲ��p�g�>�e=�xu]�O�S�����������������'���Dpd�{��hho+������x�A�0�`_S)~W         �C�{jC���ǈ}�w��@O)��/W�ԧG���£���M���B�f�[���o%��w������$�tx_�Ѹ�2�s�������������4�������n�HM���;⃡���#j�;�lLjZ	         J)�隠�O�kU� �,�}�K�T��~_����n�%�Ǽ��pX�[�Fn;��kFlR�oh�6r�C�_͂i��&3]���^uh�`����IO�%�q��>�K;��c�X忳P��WJ,���O�
s_HK���4+�(J����T�X�a           :���ۖΙ�SpH���B/�m� ��r�{���F<�hU�`�w������@ʫk�sg��n]���v���˳�mp`����X���/c6ط��T�p��v�HA�Q~�7N5�� 8�����         �������'�F?�y� ���A��v���ڐ����f/���d�b��*`��JK������?_!�6��������E���\�Yo/�����KX�B���)         @T��B����B��4�}���p��7V|#ŕ��^����ūe���}�Q�)�WQS+%�:�TU[_��]$K�씥[w���;dWi� :v�Uȟ�_$?;g� �(Q�/S����SwCjx�A)%�{��=zز���4�]oϞ=�[�n�,ߋ����K�w?�j�ī�ڵ}����Kq�����4�+7�^E�׶���QϞ=lYvjj�x�^��={ضl�a�Fw�^���5�l_�%��M4��ѓJ{�D۾i��Q]�װ}���X`(9��W�!8H�Y�R=%�l�R���o˲[�Ȑ�Jo�تU+����Ȑ�*oՋ�#؇��i�w̶m���|��Oz�m�b�i�|d]�G��a]��?�.^���=��_����~�{_�Ժ �(���U<c��A�F�Z�{�=@��>)��ζ�y������V�F���J���U�l�b��+����ګ�+�������2�K��55Ւ��;7<q�+���׫;s<rHO�QV[[#���z+++l����JRRR<S/�Ut��^�Av�W5�Ϯ����Z������*z�כ̵�}�S
����uJKK����|���H����JJJl�WתkFl � ��̓}PL��J�z�M�:ٵ@ �zg;����jv��Eؾ��^�P�;h������ݩ�g�n۟G�����%n��zw��e�󔖖Hff��9�k�u���U&��q�Vo�qr�r��<굇��g�������o4���`�Ae�������ꫮn�̇G��n���߉��۟'�W/��@�  {]%S��!Ӧ��C�rg�1O���Nv�G���N��s�^'F��/��u�ڏz�C{e?�}9թ�vg����ݙC���^gQ���v�x�^��~��l/�u�_{����qEǩ�O�6��rA���٧�_z��9�p;ܧ�u"�A�/v� �V�m�����!у�:>�Mq{��d�p���z��V�N�d"ؾ��^�P��h��C�o�;5"��r�^�:s�����u��o8�ׯ3؟�A������o��,+��_����|r�x�ӡ����raa����V���b�>  ��n�:��2mZb���ug^_	�ss�}7;�#��l�^�9]�[!���}��y�k�+�%z�ϭN��;�ܮ����u��Ө��}E��J�zM9��rz��(��rP����k�r�+Gy�xøK�N��ٵ�	�1�81�	nO�}(n��"���W��}n׫�}����4�84�}  دW�����"�	D��=��k��N�':۩�=N��vH&��}���>�+�$j���N��:��R�S�//��D�U9��+m�:U�۝��W��r�ω�^9����ծ]�So9��+��������^s��,ium��C1�=J���s;���}���n����R������ � %�_��<+�n���rʜ�a#|�[�^�d��t����D}�^�׎p�J��땐LD�����|��>ګ�I���E^	�D��Y�N��D���L9��Uvo_��WN��N��g4G9�\e����]�����]�W�rk��0�������ι��J��R�\��M䙐[�~?M�+��z	�y�>  ��T�@I�O�E�I�2Tȗ?G�r��Ë����@(G� ���y��h����a�D۾�>!m�@�W%X{E��A{-h�z��:5"��܈.�uZE$Z����h+���M�z�ھ^m��^�+�r�y�]�_�+o��Qt��^y�7(���i�zF��I���	�����_�O<���̓�YE�}�d��B}:ܧG*��� �!J��Y9s+�9q�$�`�����in=����w��!��z�[�՛��$l��E���O{�7F��u�֒�V�W����2h�'��9��^�7�o|3؟�$*7���y��'/���u�m���1��4/�2��������כ���z�|�  p�JU*�\�ę��!I ����
��\}
%ί=���Bl߸E��͠��k�3��'�[]�ߨ7�Qo|K�z���9�Qo|���F�8"%IFX= ��?N�ջ�*dݙ�7R�����D��ph� p�uZ���_�L�D1ujRm�1O)�F          7(Ȭ�}���(&槪�<��xo�d GD�  ǩ{9y�gN~C@���oD�q         �H)#'�3k~��)�I��̪G
��D�  �)�)�G��5��)�$�r�2��%         ��2�<��?�h�E�Sf�*b�H �,�}  �B�U!y�e����μc�ġ`���"��$         <@�
��eݙwJ�}��H�Ιu������]�  p�R�K�H~)�������G�y��xά1U          /Q��/$/��=o\����%���7#��H� �i�  p�R2L���̙~^���̝u�a�sfmY         x����$�8�μs�e�>=R_X�ǕRi �� �mJ
Id�9�<i��JbX0g֥b��8Y         ��)�z��|�ɟP4s�"�a���7b�M��/f  <�<i�B�aV���Jf���Ě�S}���?3+��(�	   EF3^�s����@���^�Q�}��y�T�R����!o-��:�z�C�΋�zG�����x7���������Xs��Ɂ��{��j� �+�  �
�Z�$��y�0��4�y�������K��������h%����Y��#�3��	O�i'k+3�M�V�f�c�����l_G9Y�f��*پN�^�P�������?Ys�wT��>�&���=3�GF�H��9��u�|�)�+���7�x�L�+�<E{��_��Y��w&�m�Po4)Q�'�9y�d�[7�ʭ��2gzװ�xܬ�dw� �)�<o�ۃ�Ǉ&ͺ�4�
������Ws�;I{���uI�V�;f���}���7�o�'���ר7��U�ʺ$�D���5ē�h���U|{�㫸����R�K����97�M�\<�Pٹ�ׇE�4o�с8E�  /Rj�?I�s���䯺g�}?-iuW~�P��;C�:�<5T:         p̔����4���hHjsJgޱK<$+gN?����u� �k�  �,��G�	�]���mQ�ʴi�n�Q�ܹ풤fJmH&)��         �7J|�?����s��yL�H����J�\��Y=�������Z�� ��>  <N)�f~�?P������tU���w�9�z��ڐ�!F���
e0F         �R���W������7R�sK��U����3�.Q����d�:�� #�R]�/�+$������C�G
7v|E��"d�N�GZ���"���s�5� '
         H0J�V"�����s�_W��~r��
;�.���-���r1��E��uG!�> ��  Ƙ��z
����m���a�z;��{k�}����rʟ����3�/�Eg�'	�u�
         $2%)�>߅%����+�x�
��7/g�1/w�Ԕ���c¡�x�I�KM�I @�#� @3�;���h~��6�@N���*�[+Q+�R�����H�-�*5$Fց=����|\?�z?%���J��Y�$         8$�Z*���+���~	��*1V�>:1�UJT��Qb�>��oHr(�2�o?�!����!�U���#U����W�`  q�<��n~їs�����<SPa��*>��Խ���         p��H���h��h���ה������=�A�}u F�             �1CT�t�h���}             ���"���RUU%^��nQ[�����B���ŋ�ᰴh�B��             8�s�βe�υ�t����$��>=^�.]d��͞���!)++#��1�             ��k�H��.^��B!)//x�>             ��J���P_�W�}����`            �ߧ�M�t)����ڐ 6�p��a7�B}n���y�>            ąkG�_L8Y�geHEM�<��W�˗>���X�V��0�RZZ*Ns�^B}��`            b�w��'�⬺���I��q�IzJ�Lz�mAlp:��V�/��z	���}            �y��1����5X�ewY� 68vs;��T���b�>            ļ~�Z5z�ߧ�W� ����n�W���
{�[jj�TUU�Wt��Y֮]+���,?%%E���S/��`            b�O�C~��������e͚5�,�_�~����P�>ZXXh���п?���S/��`              B�            pI����H�ʚZ�^Rn}=Vz`��L	��Hyu���˫	��C� �Ӳp��T���Ł�R�t�Z��F�B�⦽��JuJ���㓰�ݱ^$טg�;������L        ��t��	�{ʄA�dt�����Z��Pؐ����/V�?>�JJ*���գu�\�����dD�v���R���PXo�!�}�B�-XN��!��"!���M��0.�P [
K�n�1�pvfں�pX^�r�aӻM��ܶ�}��m�]�������j%�#n,�M{K�pt�|��Q]����?���\&�#��+iW���Ր�[�˺��$�����k��,*�uܶRV>K*S2�{��ʀ�oJjU�������b�ل�         ��O��Ni����O��Nm��-���y�5�löC.��kΓ��w��'�}2�{�r��ar�#����{���ۊ�����ɠ�߆I��߯�Ӌ��M<}�\8���렇��p���>�����lp߽�j]�կ.+�uiWw����.�/\y؟)���kF��|�{m��r�C/�z������������\+ ��P��Đޫ>�5��P���!��M��}z�>������J����         �>Т.�W
��ˢ�;d[Q�$��rB��r���V��Kv�<w�r��ɧ�4��h./���V>3�t�N�QZ.��Irr��rZ���s��Z^��w�?=%kv� �FO+�Q�2��F�Ӯ=H�{�3k�]��SM|�M���k�����t�P��]����w��B}U�!k�N�$/��"��y)�aW��
�}���V����_)�֔ ��vay��&        h�ͅ%�����}�Lv�<���hލZS�����^u���㿥6nty�w�?\*�-\��Խ'��$��p���L��-�%���r�ܧ����
x��Oh�{���Y2�wyw�&Gק��L~���r��ϩ���KN�����\x��|����������߫1�/`#/��"��y1��p�WC}:�7�7d9ᾘ6�c�lx_9�Ok�ߴ$��Wֆd�����-�����d�  @��)%�Z���U���R     ����g�nW�a�Y�m�\��d~�Ւ��K�6�2�Oyg�ƃ���;�j�k��C���r��^�W~�]�ů_��V �w��
4���^�d�O��C���E��ȫ��1=БƦ����u����i�߾\�=��`����+墡��)�JK�9W�)���s�=H��&���u�?�f������^�ED3��k�'��ED+���P_D2ᾘ��o~�8�o��)��~czt�.S�8A���k�������E v��Ӑ�mep���4"�2Ҭ��mSYu�UT�ƽ����Y�i��W�H�j��.m23doy������7y/�GN���]���Z�m�-/~�V6�)L�K����4Bz��1�e|�nһm�d������5���M��O����7I>���ʨ{�,)��E�g-R�e��7X���������lC;��F��^R&˶��m�}��~�7l�k;d����}����}W�M���5��u�Sh^V�6����/.���   ]S�t�q��,g�7����m�"4u���o��v���?�O��6zW�F�U5�����~�[����c��Vu��h��7���i�mݾpho�M��>ϱ����2�{Gk�`�~��Nj|$����z꾟<�����苅P_D4�}V��p�Ă��b%�A�/����~pq�/4�؜7��u,s�?^�> v�h!��>R.޷��G���Z�Z�:����Xq�>r�9c��p�������'��ҵu��OX��T�KFL=�dy`������I�D��͗X����;����Gt�/^� ����o�� [1�����S� L}�~�����t����|$s�_$�`d��V�2�w+ �߻г��E2�f����|�@9��v: ����zM?l���w��K��%���#�[��z���{�]-rὶc�>+C.�ך�+=9I���k7˻k66���å�Y��;K+����x��u��Y�[3���?�ˆwn'?=g��i�ө����תjCf��������˭;   ����ꝯ�-��u�3�� �6zV�fԠ�_��z���sO�n�7,�;�_��tѶ��B&?��̻�º�~}�)֧���*<��56ﴗ?��}��hN�/�B}�P_�ءG�x��K�N��9�ܒ5�نٰ�H�*�E�HO��-2�[�`H/��&�n���Er��G�r$ ���㬠Zz���=�#3��գZ#R����V����Դ�t�����_ן/9O�#}���g�k�]n�X�=��ON!m2ӭ�q0�	�<���KO�ז��B~��$��9���=�
�ꑞ�M{���j�;�~o�w������ɋn;�|�'���E����&�s�I�3~T���FpA_���R�������A�gn��P�e���O.�=���Ƕ/��u��Ow�����)/��Ӳ����Z7�4D~{�8��Z}��׮�Oy�m���#��cw��m�x�3����]|����a�5�PtPϴr��^r��%��Km8,   �m=[����J�6�.���? ���ߔ�o>F�,�-_m�e}b�����wut�ύ`��ʲ�ִ�W?�n��^u�\0��C�����|�T D_,��"�%��������j�/�p_l���S�B}��!���˿>]f �����S_��

������}��T+ q��_ ����Q�������#li:���ϖ[mڈ��dP�6��)k��)�O�a���5�x�j���n��N����a��(2��*`�w�e��G_o5/'օ�^_���:�UZa���G��#�k��y����th��� �E�f���Vxrc�L�{r���W=]����@'t�`g#t�:�G��#��0���wi+׎l�����=F�^�Q>��cr�^�����>�`�^��3Gt�����n;L�jk��9U�����>Z�z	�N"����%�rޟ���!��pq�#�j���ȍ�I�=j�FB}:Խpc�5���O5���k'ȅ}ڳ����Y�����t�Q���h��B�uh��^u��P��-;�Mۭ)����jÆ�>�>��?�۸VHs�yѯ���Ѹ㤳���W� �  ��dg՝�k͝%G�����}=��g�0��u���;]������M{K���[el�}��1C:��Bn���w�s]"S��أ��z�q��ix��z
�3/`�X�EM�/�C}M��z�/�
���.7�%��=�M=5�V
�wxN>Z��I?����Q�t'�ۓ��:��1��EA�Ly	����P���_���}�����0ҁ�Q�y�ONa���?X�?�|˼�Z�:�w�C��Ғ�����\y����ŋt�P5ě��[��~��W�m������2aо�mO�i��ӡ��F�ٗ�i�n9e8��F�Ф��R�N#����_&�6R�^�Q]��
�y}��C���6�C_���Mcr�<�.䥧%��TeMm��|n���aǻ�m�,��c��U�(�F��i����߽�����k뽋��z�C�r��}��f���eɖ�5z����.�>0(�G�"=����G��5��/�i����ij��v}۶��f���������[���S�t�}����ٻ�(έ��xB<�� ��ݡ�B��R�W��[���u�
-�P��!�G��qw7�=o��"�ldv����_&�͔��ʼ���{�.��~2w������A�������R���������v�B�KC<2�G��I_�@�e����������:+�/��+�~�g    ��L������iM^��+W��	p��F  M��
 1K����rH����uE��-Г��y���j~��ôm�\Ek���;n(]����;���m� M��>9U�}��S��z��b�{/�iK�ON���:�7�*u�y���������P9ԧ�'#<��������A����
 h���W��������׸�/����7y+х}{���d����@p��-�s��+�JN|���k�z��p�h�Wg��mY��F���G\����ؖ+�u^�_Jc<]i~O��I���p���,L�^���m���x }����q��mWo���x����ly��~m�7��Ә��<�p���u�p���'��K'KZ��K��k�5,��A`�	s�V��r�<�q���וߗN!����?z�Cmk頪14>�_�[���x��g牱�w��<^�t��{¹��e졽O-��9)�����g��K�7��)�21�7&���|�q�-�;ꋶ�\+}���8�:s�V��B�ŕU�;q��_���,��#� �   �����]1>�yy�q�&��D5yր?;J�= Ԅ`��p;%�R�|A�[��m�)Z���*x��=�f���_��Ќ/�Z<�&~�QѮ���<X�[ Z�47m
����ӦP���];rO�O�B}rUᾃ�I���	���տ���\	���q� � ��
4#���南n�����.Ҙ�#�D�O�fZ=��^:��"E;����<���\���q�hߵ(Q����P�߄�f���6[KTS�CDZ6��ǟ>�w�Fz��*�ӽ=˸�!��o7R2i������k������53��w7�P�վ��B��)�㓃}|�v�WD�${v_y[[w�F�O��ܦ#4���h�+�=��*�?��B��	V)��-��_Z"��<J_�P��򊆏���ա�;x#�F�O���DXJ^��K�{C]ch�Ί�IseF@s0NJa8�����&�����C}�?�s��#a���&�c�_��y�AT>.4ɍw��]�RS𘰼�􏧮4)ԧ���>9H��-:��ߑ'8    ����jG?,��(��ڎjU��Ɋ�O!��T�'��+� @���� #sf�������H�������'��L��#��������B];Y����؉6E<\[^��s[��$OC}r����1�'ww��C}=C��������V�۱�y��j��v��vE�`��41��  ���ڂ���+��XE���>~��k�J����J��q�sWǕ����i7ږl:�	`��f��������'�O�s?%�~���'�8���V��2/{kzw�pю�Xx�8��-;?W%����[�*3��DȢ�����d�y���1i��i_]��HXl�����_��P!$v䥭���yc�1˕��9�q����_̔Z�r�Qy�J��s10���C~.r%�i��M�yZ^�xB-��%�w����E2��
���עi�[hۊ9�b�#r8y��%������ܱ��l�|��k�    4Go�N���9��w<�cu@H��7�����4E���v�� ����y�x���{���'���_(���{�i��/�?���yj����k����w��}}�)I�h�����q��KD ��A6�1Z��p_���t�g2�G_ ��|�p�{t E{!h[� ;wK��_De�� �h  ��Z)��i� _'S��3����>��X���6R��x��B{�R��fPU(�9t�o>�:vQ�x2W�Zԯ��}�� N��E���|��U�
�����<X���Q�c��5�OQzn)��cfx�q��%�I�+��NT�w.ǧ*&0ڙK.���H�"���#���4��#�~q	}�2}���V��6U:����
�Zz���ݒ��<�}GJcXГQ�JGPBM�q+�xb�����I��������V�ң�sg�wY3���,�:    ���֒����8g��L���d��7�ݑ�<6[1����3���� ��> ��J.J�3w�D���/>�|&�/�6o�p6&I�x����@W�v=9OQQ���?�>�  j�S�>*`u�]u!Z�������K�rPKҭh�)u���!ܢ\EJy�  M��3W�S�G�;���K��̔�tekj"�`_vQ�b��4�:�R�e+3J�ɯs�ʏմ ���������Ӣ�1��8<%���/��O�z����IJ�����xh����mj��M�/aD���-z��P�[�2nY�%��[Ct�Z&d�*2�<���j����cI|�n�F�,/.
�1�]��x�.�j�d���;��������/$-���3��')Q~uPn�Q��4�-�s�\Q�r�����Tzx�>��m-[����Tέ�|����o��LR��s�3	��>��D��JۚX��    ��|�������\���m'����n����٢*9���y�u 4�} �tP���s�z����r���q����@\9�-����ha��`��w���sт  @�̕*�(J�*G)4bn$�ߍ�Ս��X�����RJ�v����A?[�q��v֢R����[%�TPZ.�ᰔ,
IJ��q��C�"Ӳ�Ƹ���ШgQ��J�\=���P�����TZ!���,��re������O�*�����&&]Յ��w4*��-Ov���l��qK^�-���K=��{@���9��e�h�[�i|��z&�>�5R<�6_��u)_pxe� ��!U�qR������������U�z���Zҙ�����ڤ����~����>�PT�|s�)E�MS)W߳7�H�AGG��W���؈��ES�B�V�#W+3�ڻ+���Z�f7I]Pb�g�#�
���A��{����l���ύ�/>��g��� 盓����{~|�f�   �#��ɓr�?�o�F�l<��q;_g[��W^�����} ��> 	�21�i��*�O�/�c�qu>~��k�`[:�7}}�b��x��������ށ�c 	  @ڔۙ5�E���;�͍T�Xޚ���]D�!�ԕ��OWRiGPD�
&�^�C���qџ/�q��ǓW4����
L�l�P���S@'#�E5U�2a �v�D�E������>4�Fvs���7IW�~~l?���]1�W��\<Q(I��\��J���$��I���h�0��Lp������&o�TB�����	9�:_��M�l{yFx����G��W�덅���9����\TG��M�N�
��5�7��#=>�O,s0"��}TAn-7R2��=���gEh�'�����&5�>w�z����igE'_\B���۷]	ϓ�O_�y}�� 7ڸ|�:u��8R��%��,�׃^��?ZT�7~�ƓbcjLc����snO�O,LUZ��g���"�:6�U��[4A\��V��5����ܔ:~��q0~�w0��}�bl���V�B�7K��(Rۿ�YT^Y)B����1�ϭS��,�k�D�<��љ" .e��i"����=K;�Mֆ/��q���!��ڡg�G�����רN�#ٹ˼�����dW�y��zoc�5   ����O�Ut��);wr��z��ׇ��7?6[q�Jv��֮� �	�> 	�A*�h,��r����s�hg�Ve��c��Z_��ǆ�*~��8�   ҦwW0�Y׭�Z���*�zh:���O�X��N��J�<�����|Q����i�wW���ɇd�{{З��*.�);vK�t�J!�^\���/�q�vܦ����9������I�������#�������g��]��V!4b��KS{u��d�!�i��.�>����l[�T���w'.׺����2nO�Q � �^��ӏ�#d|\v�d�d|v�<�,uv��'ο��Ŋʌ\=n|wQ!^~��!h��,��mm��}����C�d��w�Z<QT�;K�Rhu@�X���+{|�)������G���D��E��rw��O̭�~oGՂ���[Z�M����h�7��ӣ��듇�0#|������3%U��e�Q�:�_��ymv�D��*�e�������P,{}�*���tT7W1)�1�/�p;��-ow[+�!u|��q%bm��ы�����N��?�;�ޝ>��E@56+��s���R|v��+�Y�?߻Y�Q_��[+WK�����e    ���s|�ڹ�|d���e����f�ù��+�)Ɓ���;��� ��} ����mx7\����l�pC��ԫ̓}��W)�hS   ��m-�?2�F�GWX��_��t������lQ����\Q���?�?����n;�Y��h�ҩb�ká��/,��7�AA�|9�����/�^�K��̪�z��@n7�{�J����Bp[>�?�9�ܬ�D�S���دg��&x��[}��Mm��=��wyҔ+�p�����@_�����v�o�.����' �[m�%�o�A-O�-�92�m���cA_O�3�5����Ն�?�)�p�g��S�M���96�����zݸ%{}-װ0�/��z�F�����s������{ϐ&��*�}�����*U��3����������gSt�{�'6W���ھb.�r�fUQeWe�W^��+�i;���i;�-;W����
V�Ý�dD<-�c�$�e    ����X���;|�=���&����O�Wt��ɟ�o:J�����hc��Lyp*<5KL6d˕p�h�HEՅy~��ڎ�b=    ��A�J^��������x��ա�>��b_W;QQya��0���簢e-�@� W��4��pK�C7n��ph��E�>������E��[p؋/��l���ɭ@3����q7����� 
MJWy�,El�?җ=V��	U���m?!*(>?��8v���?��L�����~~nl�&�wKs[�3�מ��<zfL���럋7��m���!��l�n�}�T�|��4�rq�f����+{=�n��rd�U��.?9T����U��ږ�yR�s�n����q%,�Ŗ��ZRM�f��L��̑"���}Hq�uy��^6�3[Sq�4��ڧ#H���F��S���Ǉ��oA��@�*;Ƨ����>>G|敲��^Ο��m����%}���J	_��*,�����!/�����������ˣh��pIo+   @{�]v>1�����G�ci�ݢ@Sp���+�(B}�/\�g7њτVVVԣG�Y�����J�c���un��l{K4�} m�R���I�>.��]�O�!��2r���F�G[% h<G;��݉�KԿЛ_�G�撔9;X�OoG*.�S{]y����8�2W�N��ӎ����^W�l{/H|{A}!o=B�J���"�z%\����EŲgF���g�n9�U�r�Z�r����#�W�c�d���O�@���.qAW��}ȶyJ�.���&S�㹵'H�_Ƴxy�����F��C9o�:Eۃn�
>|^���~��q��g�Ka��0_��U��x�_��ȡS���{@�"�[���Lza�Q�:~��p���5��#u�hLI��}�]$~��:�j��4Z���.�;�	���W���j��2�����W�����(Z9rKG�L�����TPRJ��Ų�M�h}�m!K4$ ����Ͷ.��s���"M�v�M�^8��TW��4��	�����N�&f{%�����ωꄌ�Қ���c�~�.��&z��-U���h�dh~�����^{9XS7��v��j*��fl�OE�e��8�ϛ��t#%CTx�z�    ��+y%m>G�q�mHPB�p�yW~v�6�<��ǔ��?���q�g�1r)����>���۲�nn��CR�޶�`@2��U���[6���5�ҁ���&���!_�IE�Mo�RXT@i""�I@:z���ˎ�B+����!�����.�j������t5�6����i�M����8���XU)�?2������g*�hƾ8z�F�O_Կ��**�p�Fj�}\�l~uKEn���P㶜��%Z��g�(Q��)C����Oi���-���|��9Z�*&�ܤP����#���ӆ�@7G�
$�	a���ᆗ�S|ϕ45�-fcp���*��9�ƕ�Au\��Zx��7�n��Ŏ���s�&>/puv1�}~�_"nR�����a���9D m�CP   @;YU�?3�]��K�������;�Yw}P5o�!@)��rȭ���u���-,,�ל�����Z�kn^E�O3 �І�{wev���-�� h,���xPpp��}�KIϣ�RFG���v��PjR�/��Cn������5���֢@���Z��s�Ɉ�+O�@F`L��`�^�?Hs:"A�̍��ʜb3�S���W>@ĭ�k/�� Q�l���E��7@�����m*����[
������*qX��}�<q�0�t��n�� hI�>�-;    �;[Sc�ىz�[�ʹ\ݘ'
s&���
��)&#Gt�	�����;@ki�������m��i��[kn�<���>� ��{5�:���E�  ����дp������+(ѡ��$Q��C�	�5u{�ueۛ�q������j����b9>�����A9no��� ]r^�b�+�I)�ggv����mȑ�[��ם�ϣ3E;VnI���K��8�q��큱���yn���Z�)�       @�p�<?Ozl�/rw$]�ƿy��R\
�>,&�VTb�g�w��u}��&m�ڡ>9s��}�٭[�����>̀�z�6�daJc=��g���'��h�I�Y>K���=��g� �L���=($4�JJ+||^�f���Dح�=_ץҲ��WXJ��	"䦉�������������\�\R^^���w���~��rk[�I����b�B�����x���v���lQ���~�r�<Մ��<پ����o]��N�~n�}�>�N�hw+5�6S�����)��~n���     �%�yk_�9���<�@W�R�)(!�r�����]�wu���t�j'�5�@w�ŉ�����0��'�����,(�Фt1&q4<V��hwksZ�l�Wi,�w���G������� @}mr�33�jS�Zᾶ�^����>�6����5f}��I��R����	��s�0�q�nt��- h*n���hM�i��O��&M�|��ꐃ�%��&5�ش���5j{3K�U��ѡ>4��Uʶ�ѿ�h��r5��[$��ˬ�b�rc�Ӟ�I�9?m�-���|�y���7%���dy����B�9Y�JC��L˦��"�&����e�j�����e^���O    �vq�2��d���x��~�K�啕t4,�>� B~ �:;��ǉ�+񩴡��C��ϛ�iD�Q}鑡>�`������IAIm�N�
l��t���}O/�N�Ɗ��VT��z�Yyb\�;z0k��h,�&�v���ՎL�}=l�г�h֪������:�&��>�4��Ӳ�>�l/�}҆`@���Y�g�/�7y}���`���  4^_W;��׽��m���^�6��Qb��'�zr�fP��t�Nϡ�7�H���f�x,�����fZ�|�Ϟʕ�T��Df��F�V����&}ҕx;n��3۷�X�q�v�O��b׆���1�D5���-�׶����Q"��*ޥ���ҧsǐ�����߲�V�F�V    ����o���U,?��嗴�߆��L+�����<Wg媑�\h�C���ذ���d瞓zva�g72m��\����#���Pz~]�O粚ԅ�+�����9B'"���U�B{k� �/!'_#Bnr<6����*��Ɓ����~���]���s�$U\x��%���[���ɡs��j�0(_�D��������!��_�L#?����� �^I%�&gn^U����}R�^����>�6�'�];Y*��g����M����i� ��N�y�H��..  h#C�ݵj��Ah�&���'*���^um`����ͺ�����IJ��ɍ�1kxLw7�ֈg�*81�f��J;��+�����|؋��r�ζ���{����.6�biF=<]\08Gb�����J��&zdkj"�}]�i��k�s���P     @���h#&�����ϒ���1�����j}������g��ѝIrEe���I%����R����?,�(7щ��&x��;S��y����aH���I��t�>���n�N�k]xd.��E=�IOW�"R�D�Ty����Eӽ=jt��ȡO^��g��ߤ����+狀�\J^�؟ܖ�K'�61R��W�5:O�l�h���p�\~~�p<u�hL_�@R4��E�����e�ʁ>9�-�݈�/揥�{�*��{u] �q�r��p_s�u�.YR�^�qW7�� ��ҁ�j|��J�Z���b�Y�O������¾������O��l����Y��Ĝ|   ���M�;;6:�V�՟�xv}�g��-�}ܮu�_7�x)�Q�#9�����v��'�u4�b����i;ns3�-�i�,�v�$~�liFK����
��).�     4��g�R������=��ǹP*�>�s�q=��sǈ	L�=f�~����[_~�!2�}=y3��so��{e�@zc��zC���j�D�ő^�|T��?qYt��I�]|.�������~t,<�֝�&*ʗhx�������AS��=;ӓ��Ч��ω��9����]-"�X�t�hQ�r�{$y��A���J��w��s1I����ř>�9���ڋ�a'#����~�������0_��}g�0���I�dǁ�L��E|�n+�>��P�2������4ɫ39Z�Ҕv��������f�Z1��neeM�4CC#�k.��^�f�^P�} ��?���V�g�.7�km6_	S�؃��U
���)�`k��)>�  h��^��攡-��o�_�-W�I
8�7��C��s���J�����RT<c�Q�$E{C���q��c�}�ci�4��ʹk�<q�A�x�˞�H�gn*h�VU�l=..:� mII��㓿�DO���G�����?}w⒨���`6     ���\�)|��Tv[<�KL�Q��o���V��R8_�ixR��Ț��\%���[4��Mt���A!��6��������hWz4<���,س�XoOH�J���di&Zx��_��9�ձ�$e��#D�U>���!&�qy�1�Pȷ���v���nw6Z�.r��g���>��6i0����篋���P?_C��E@����A1����^�v���_��\���kv�S]�����M�n3mX>��y��W�ѩ�16�c2�n;A���_:U��EGd�i����XU�ג2D�u���HXl��6���'�e>���J+@c�� �m��he���QƚKp_�KU{�ۮܤO��gX/�ɂ��]MP�   ���;S���pfk���QK���yqk���DD�X�MRt).�~�����hebDY�ō^�]��j���`��K�y�j;��5{�m]��٤	�������%�Չ�z���_���Xu4����Y�챙Et3-[T�;v��D%��     ��tw�u}4s�=?��P����EQݍ۵��S�����M��]W������s��|��wBa�zm�	qMH����8~���a�W&���_���'rź���.��oцV^����P��o|�r�aM�6�����;��+ح���R}d�7�v�D�M"��Wn�`�Zu�
WW*����|�����x
�ޗ��w�͘�T���MG�m�!��6��7&}���SL��ju�ъ�~�fmN�d�}�J��^UD���'TO�4�G�  ��Y Z��z�����7�e��E%t4,�F�=�]݆`   @K��L��IW���́�}����@�x �dD��     H	O>�[x���s����U�|�+�I��UUE{9q���M�꬘��ݏ^�O���-��T�$�g\���s|�K~�Aڎߌ7{3��Ǔܻ�>����7�ײ�����H�N2�V����\�z�������?�gј���i������/&�)����SW�~���	���C�}���I�ku����Z���g�QXJ����!W��N]�>�������Sv\r8�9�ps��n  ��`�K�>_�l���hu�?��M�R����ǌ�j���>/n   �Yx��9>'�w�����h       ڻ��zR�[�T���*g��_r�S2H�py�!����ϕ�oe��h򀕔8Y���)�����tv_���v���1ʸ���a��igEC�:iT�OYJ^��X���+4��3=8����h7��@߸j���m�Zjp'��6�'�X"{N����hmil(�#�t�j��[/{�:q�[�S?��[j̪�����;9ť�����; p�MnO��,5\���rUɷ��7v�Rk}��{��mv6FZ�E @�!�     b �)-Z��Z��S��L�n��:�[}D'      @{�-W9���:�X�e|*�����4�i���7w����.mHyukϢ�2�RE^IUp�POz�3�*�u�ݴ53_��sTj�ʹ�3Q	"���%��÷Wd�=�k]<��"��8�򄁔��O��	&)q��`Ǖ����I�e-���,�~u�`g��o�!7)�_�������k �*�Fw���������2����A�)B�O��+&(��/@����Ĉ�۟��W|_TVN[.����ӭ��d�	  ��}   I())%C�>��̘�s�����
244k�q�f(;��Y�R���Z������-���5q�����D�x����EkU�      ����D��:�r�X�Ý��u���n��=��ǹ��3�&<5K|554a����PWW|�b�1��MG#^�;�YTZ�}%�o���2�����6�+.�5gCĭ��5�?�'-؋:�J/�%��@_|M�Ϋ�1<ޕ�_(�Y*��Տ�h`@R��.^�\,�hJ���/4�������=㖼��6�,�Pz��5��[�ѯL����Is�<)�V�G%�m��̥��2E���@OT6��������hd72��U���8&K��^]h��  �	�>   �Gjj:UT萡�Q��uur��
���,�T)��TY�';	o����Ft�ҙ�HS%�����&������<����j�ϾzЊ=?��h����<'Ɂ����/�@+G�՘�΃���D?��R�Lem���ut�����$�۫����    �4���e��|>o��\������6�*�o� w�?Sn��ˢU��e]]��SR�H��cH����O\�q�|�v�� #=�{�)����Z|զ�q`��=���gij�b\��Bz)ע��C=��x�˫љ6�N���p�J��IoN"����&�}���k}�.N�����\���1��ꪇ��W�l�/��1�/�U�R��Ύ��X����9��_3[h ��!�   5p�����Q���Z5P���>����x�g��lN�eK�	�ix{���$�RM�ަ⁜��x7�8�T�O��j�����=1�O��,�-�KJ��3�����b&v{�ǲi4��]T(��p5i��M�q�n��G>a{�͟N�D���    ���Wo�����!�L�=����%b�'.i]��G��?���;�`���ٚVM�L��xʾk�TXZF&���A�7$��6m�FoO*�t�/�p�2���َFz���Uڄ'���o����0������RKm�>(�����^T���<н*0�J;��v#%��^�I�z����YH�e����[��G:::�=��4��]���1���v{�u��>��&�k^�+������R��ʠ�8�w4����9���[�R1�>���ϯ�  �:�   ������\��WM
�%��Piq5�޻;�CJHԜJv�1����D�����r���&�1[�g0sh�(���       �^�Y���2}1�h��������ՄTj/��!�e�gZ�$�{�L��x#Op�`&�5�ۮ'��c�1I�~�0�{@0=6̗ޓ�gnɻ: DTH�۰�����)"Tā��W���h�J	��>�Lˇ��}�ᬑ���5�g��ߘ<D,g��2n1�A����,����FR�▣���I�;9����i�Lj�6�\y�6�}�)���=~��N��#ZCO��L��E�]�2ʕ�-3�o�l�a�X�s�fj&]�K�}��1�;Q���?��󛎪�>'[:���  ��>   �	����D���m�K� �KM/�Rrk��ѝ��3݊�ER��P��b{;��Ɛ���#a�-���ƇH�bJ�.��̑bPK����֝��u-�    @::�XPg���MQ*;w	MJ�-����!]p{W�f�
W��}���?���?yY�'-Q�e�q��6�� ��
tq�o�p?���Ҝh���+��٘��biF{�^@�nܢ�o��l��۟��Z��?�7���_v�d�Rye��7�Å*�-�c 1G��Kۓ����?w4�����>z��g\=�ߗf�v�'3��}gD;���!#==��\�콧�ý0������ER���)�m�oM��>�>�Xx,=��P���_�8�x� =���_�.nچä�r˯��Nv  ��>   ���B:z�yx@�Ļ�$�dɶ�f����JILL�c�ͳ��J�js��q��U�tv�wg�_��9�3(���@Q��     ��tu��eSh��5���r�!q.��f�v���D��U�u~��J��~B�c0P;�p�e�0�v�x��dI/��/�4uU�����lqk����E1+�������--�}�}h��=�䞝ōq��B�@W �
~u�N����DR�?4��|�A,K��jsኌ�?K��=J|��խ���~&�֟�N/�H�Vf�ټ1������%��z�Y�hY��^n{+U܍c�{������F�����X��Ɏ��q)"��P��}/�W�_���1��ц�uuĤm  ��   ��WRL|��	ZVVN1�)�^��U�����t��MDs������q���Ӓm     �ቑ~��c&��j�D:+U���@?�7Q�c\�,8!���h.��7����ԡ�b����Z9���yEF�r�bMP\VN�~�!�/�3mY�)��e�����M����!�$UR�[{���r���>9�O��sպ�U6Y�����#B|�����ުh�9��c�	0�Y�'��`���.u���kI��  U�     �+_7��[�2�;�D��=#.8h��,'��^���1�33��"L����^    �7X�jxs�E{��I���p�D�h��}�)�%\�4��^�q��\	�o�'/q~��+�9B.\�����f?W{���"Ҳ��W=/�����~}]�����I�v��5�z�E�笼���d�$�؎�n5���Ͽ�_����mw�H���=�wW���l�V��[M�+�j�	  M�`     �8O7�g�,ъA�J|*}�/����"     ����Ѭ�XqyE�5O�����p_��\�}\���&М���%�����6�K�Ң~=?�@�Kc�������e�Q���dal(Z���SAi%��6��x��*�]�'gЄo6�9��� �驹b|������R%ˎGv#Y�j}a)���?  ��     �y�[�jn<�z�f�����jG����嵁�(������̤F�/)'��&��LqS��+�b�9     �*�=~I���X4�:�>vQ�*%q�w���1���ҲA���shɫ����Ίh>�d�jV������C�c���D/w�7�H%et-9���FQT�j���oK���od�a�V�{�$R�-��7�  � �v��Ҍt:P�(*+��|�w �~O��+.��i�W���1�J��ꁚ7w��=!�u�opg'zw�p�|�z���}ws�0��{7˺x�T�}م�U���D�>_'^����}hXWg��,��r+����U�'Ґ.N$U�����&�Q��C%��   �~䗔���i��D�Cu�$���ϓ&����>�9����%/h�v7���X��Q�h�b8��M,_�O�mA{h���1��˦�:������l0���_�L�����q�˶��  М� �v�PO�ł}eh����5�su�3.���%�������k*���l=QX�^���˶�[���v4h��-�����ʛ�ަih�   �5��I����h�?��S^YI�l<L������wCK^�F�V�f�T����'���i�H*߿/m=F��	&�nJ�ߗ��_��Ԙ��'�RO�Z����@��]�i�{("�A  �6�     �p+�^�|�E��䤂g�sK/��lK�eۭ͂RiA_O���܉.�j�����¾w���ooP;�^   h���/Z�q������y��J�D��wCK^   �}8s�"�ǡ�ף�8������J��}<Ax��i�/��8  @kC�     (2=[ܴW8��q�%m���|��H�)�����ζ   ڟ��rzj�!���Q9����G.�&iL޻�%�v�bcA_.'�W��B��Eh����髴/4�@{p������ϲ����M9Y���A��2waZ�Ǟ�^Sh��}6w��u25�]+�Ѣ�vJj3�6���nG����|kN�m{A=�    @�q5>U����R�p��*U&�}�N9���o{�^   h���/�Wi��>��=Mm���-x�ڍ�F���*�wGh���'�Wۘ�+�������o���˟9_kP�td<����N��:��'Y�����}����g���di*�3
�(��� ԡ��O%%%�&E�e�MLL�m}T\\,�����M	��>     h7��J臓�E���r�/�=�v/���P�D��e��51��N��3�5e{����~��xn��}�Oi�   �~���M�ٹQ-y5��ۍl�{7n��� o��\�&��eo�l��
g ͽ���b�_s��.������Z�Ղ�?~���q<��غ���[@O��+�_6=6����M��cIqu��7�&z���l��x���L�!�I�2~�Cv��z�~��ʶ���T��᜝�)!!Ara7����5k�O�����TZ*�`,W,((@�Ob�    �v��]��m]%e$uo���6�&lo{;�  �}��O�?D��V�%o{k�{�g��#a�ВZW#[u�$�4���x��4�Ӎ~\�~���iU@'9�@T���}�&� ��d��G��I���C7n�&�ҫ�Y6����DDxrl7{q{l��2��0����䡾����"�pW��PH�}            i����g���d-y5���j�����ց�~ގj�   w�O�P����{FT�{c�2�ӥ��A����6�R��ԉ�<8M����jeF���/��9�ʿ�6��k�P��T�}�I�}     �0�����Ս�L:�x�cܛޟ1��u��֬��     �}���:S7ۺ[8jb^k#z{��f]'WO{``/ZJ�68���0�f[���!I�r�4����
��Z���.9YH�ܰ�δbx;ڿJ;8[���ܿ�����+����ؿR�ʫ��t4&]]�'|z(P��x\���?�F���OQ�9$u�.�����̥������@�F�>3��	K3��ա/�#s#���%hmݦ��B}rm�"�'e�    �`kjL?<CTw�/)��_���qFzzd��#����P
K�$      uqKާ6�ݒW[𲾮�djh�����	��6�feNs��S{���X�EOʞ����؉�_ZBR�fݾ�o\֝�î�zv�����lK'��~�*7+�v��<wG�ʷ��q��S/Jw��H���[;QXUv+-����-B��/�J_�HR6���쳆�X����n�ԼB�����3������ܘ�ą9�ȟM8 ��*��ڡ>���^��4�}      �0v���wv�St�z�M�tt�Q}��MG	     �9����N_��k���sMm��ne�L���i��ZB��E�gnmɡ-�.��i�j~��OPB�ڿJJ�ywmT���:}�Jd�7>�7V�_�0��l���b��'k������ӥ����Id��G�N$����4����U��'

����fb�^��4�}     w��1<Q�}zJU!��?��;gt��1�no�	x���!����U�?\-��ݍ�.��{�\?O����bp     �9��/��;� wG�=����yJ�Z��E�e����Ϊ�W�Wt��L�C7b�Z���)��GR�W\J19Ե�%���-��5/h�*��{&*�^�Qk}R߿�^96+�ܭͩ��M�ڗj����!�ע�Z��yGZ9�I?9d��Ƃ���~���I�x���C�铃�DU��XB��e�����f)��,�ml�hGP�h���љdb�Oύ�';t���'k��h-���J}m��6ĭ�k�#4�}     �P��,n��v��H�fU[��U*��T��r�K���ݾ?qY�̍hxWg:v�      �O����Գ9����ŵ��d��=��4���D5��Rߑ��:��	���9&����+5[5rkK)�W��`�\z�����۪�z���-i7���}���;����L�rv���_o�N��1޿�����\�k����t�z-�S����I��_k�z6]�
����K&I:�'�N�-Pi��dD<��emZ>Ktw�cWOW�^�v�>hv�������Y���~�U�S���ݼy����[d���m�uC�@�     ����by_�z��YHR�����1p�G�     �_��I��r\���vO��8���lG����u���S�`x�U8y|Ajn�*�_�o]ʂd�s���X�mV'�WTzg��Kr�f��f��z�g�&��,�nb��Y�`_QY��󷐤�3A�\ݒ�65=���J���8��]|-Yz�(9����щ4s�VںbY��c�|Ew��7%��֡C���a�����Iz�$�^3��=<IWW:�C�    �ګ�N�ۻN�Ⱥ�JZ�T���-�s(*=[����͈�,쓯      ��(����I��Վ\�����H�7�f/�QTF�XS�x����4�$U�����L���֞�l���"(�������%���ݸ*c?W{rn/�������y=R޿�bl��5�h ��I�U�6�M�E�>�2�
g��im[1G<��M�t��W	  Z�}     �x&.��#��F�kRNA��S~��~       ڛ��T�b>N�D{Cm��'n����V�'nƑ6������+Pr������������mO���kv�@4��3��R�w�y���v<1OL�^2��h�-���DLવ)y��+  �}     @�Z1�6\Yp��p
��$�K��|�nf�i�       �-��lߪִ���
�%��ӻ{�Ų���V��kk�V�����I&h{�孥���N�/%�@�������hx�byq�F�ص����fڹr.9Z�� 7���`ޑ���BS{u���"�'�c�ג�E5�5gC(�X��@+G���=��q�ɡ@ �C�     ��FԐ��"qk������[,�6�       -��s����<��c	��W�����m)*=[�G�aoMӽ����)%��7j�>{���#wks�}0c=3����X]���d+n+�����79��igE���Fz����$� h�     ZϺ{a� ���*E�e�TeV��-MI�C��}[�u�ZU�d4         ���Z������#C}���^ǭ�\�����bcA�{�P_iE]�M��񩔔�O���4�͞&��"~�Vf���94��퍮��c��,_#� ��>    �`kjLO��'J����gCH��C.����F�{.�f�ٛ7%h         �f_�Hۯ��%eM^O\VM�n�t�߇�f4]|v�v&XTͨer<������lcA&���}i������J����!]����o�F���  �,�    4��}����x��{��;N�����z�YwD         @��*,�搒W(n���Rdz6UT��9�ZR-�m'�~i	��R7[K�ͅ��Ǫ���J�L*�ם�Fщ�h ͹� �&3#272��������J  ���	,�CC�8���	啔�vG�n��{��5oilH/OH������Մ�Zg�IIpb��q�'�����5�u���)=9��XN�/��l           ��T�vȏ;q3�&z�����mU�}9�� �[�N�to ̓` �z::d��K�Ai� @�-ؓ�Z0N̂S�eoM�{v�G����_v�R��O�Z2��M�j<�Bl2��P �#J�KY�������d�+nxt��q%�4j=��w��3�¸*L�݉K��           �aI9��e.d���z҄�0�ێ� �C�    @��.N�ݢ	�ӡC���aoM>4���-�[� �6:�>=HGU�9'�������I���i	�{�?m��`8O_W�f�t��g�$��g�J��3A           ��݅�RUh�lgf"����H�A ���    P��Q��^Va1�;�B�2D��>.v���u4ԧ~���������!��_�=�'�dD<i�Ҋ
Z�f7{�>��h,nr|�:KW�SE��l�߅��@���b���"���KJ�5{����           �q\,�hXWg��щ�ΧsF��B9E%���� ��>    �j�j����X��ȡ)�o�ъvm`(}�2�{zٛ��[S���s���<K_�@e���b3si�l��xp�t�?�A�}=�M	�y���}t#9�           ��ޙ6�tu�
��I��Ĵz?�ۃ��u�o�>]�� h&�     ���X~c�ZOz�ҳ�}gD%;��w��U����O͢	�n	��!cC�~�����<J�
�         ��>]�ϋ"ӳi_h4�-��C,��W��{\d�.<����1b��
q� �|�    T�bc�X>W�㎇߹/:#�~9Dچ[辿�}q����JC�:�@7G�15&+C��#�{Et9>��D%О�(�=         �6�*j#=\��!ޢJ����k�	h�Y��&P��b}�ڎV��p�r0�HEe������ @s �    P�ܨ�2]Z~���%)7�J+*�@W���J��J�=C�/)�o�         @{��`C��{�{���14�^�6���9db�/����ZR����BK��8+:�v@�    �������W\R��8�WTZNƺ�RK�^          �6�ia�������d{��\!������' ut���m+撵�����3A���������}�p����U�~<y� @{ �    ��
Գ       ���Ȁ��m��ȴl�,,��1::�,�n4�ۃ\��D0&&#���F��1h!(qFz����D췌��F����p���Y���O�=��ʑ}��H��D)�ڝ��UtoQV){�
�mۆ�i��p��@�,i������D|�^vl������/OH]l,������p��++	 ��}             �6�j���4��g��d�ߖ�"�ŸџM�.5W��U�h��$��k�Q_�3��#�6y�<q�����Π��p�XnH�N����b�����3����Ԅ^�_,�g�i\������̷���U��v�z=��0��p�k����Z,�g�Qz~ソP;7ksڹr�ƲM���1V�Bʽk'K�������b�+P����qY�4�� ҄`    �]�t���]���\�칆�n�dRqY9       ԇ+�9X��q���B��Ԍ�uV&F���y��`s�}�=�i��h���PrNmy|�u�{<epgGڵr����)*!��G�z��Ɖv��x|��ᾴ��=���h~�Z�ד��U�kS^q)����d�8�J�n��>��֊���X,���8��D�'�{��'撳����_C�\����|����P���5���"�~ ��}     w�h��DC��S�2��ut=9�       �}���\����`Md�E�g��kѢ�2Ľ;m��ᦨvǭ\��O�ST�����Y#�w+3Wlc7[K1����ޚ2�NG�+�3i��݉Kt-)���D��#�D�V���g��7%��
K��8�QPRFa)���@%�*�>Wjz�p��6�	�ER3��}>o�=�>efF�ǲi�ّ���� �*\����ݧ��s�m�����׋��پ�D%:eʭv�zZe�mE�����Ǯ'�Qg���HZ�n���rU�?L���s�j���ї�R�r�.H�}��\:���*oc-�������)6��nkƤ:           hSzu�O�>e�Ao�:E�N_�O�ٙ�<8�`	����>����C���\��hQu���l+���o� �c�|��9ch�l;�T����ܟ�Sai�b='n����a"�3���� Ɇ�d��Ù#�ѡ>"$���S~�?��8���!#C���],s �HI
o���)��bl
�%;~/�&���>���JϏ�/#��W&$s#zm�	\��U���py��q�j��>�¤��2��x�6]
������~}PW'Scіܣ�����h�_���B�P���e�A��=0����*�w*"^�� �ûh�����X������+Nd\���O_��2�fh  @��ʣ+�-�n��      h_�tv�?�����L_W��;g4�d�RHb:��t�"4����DhL:�u������H��Zf�B�{wU��>;X#���.n���lGK������S����HɤO�g������lI������t���^����j�8�Գ3�\�r�KISq5®��>^g�ڪ�w�*�����H��p���wpQ]i�_�ޛtT{�$�DMli��kʚd�ۗd[���l6�h��M�{Q�)�{��{��3H`�3���0w�s83Ý{���c��u�X��hIO��a2�;+�(��bc�V�2� �S���ݖUX,��ˏGҡ�dhm\�v��۩����~gT���F�+�v6����*붵���R��F��xm���� ڈ�����i���������l ����+��K�Ey-^W~Q;y�d���N��xe�y�D�O%����ܩo��x]������{~[��mG�       �%D���S����|�~31;�ܜ���DE�����1ɢ2�>�y�>�u\�t�w�NA�q+���B��墳���:����y�c����Y}*J��@�u��e�tC}���H|
9*s9"�G[��@���|���5��;M�����/��[g �Ú�?Mg��i�����:����66��$�-~��Q�
���v�/��K���s����R���������}��c�$�ӷ�Rg���/�n|iU��?77W��������M\Z�l��!���\��'҃+�Љ�Y  �FC��x��s�TT�����Szz
����CYi̫�{Foqƛ_dFWIv�?̋N�����7=#�        �a��)��
ϥ�,���JQJ�!��O.���}DЏ�������z�Ҳh�7�Ek�!ݼD���~���L���)�u�\��;����CAI�[[Rw7'��U}R����~;@�:.���-�?�/�4}9+�rxc�c�h��kD5FS�Q]�����I.ˡM���Os�����
!����-Mn/	��8T���)4p��ַ��%*B�hj���� �j��7���v�`��Z���tvv��sr�7�ơ���2jM<^'��m+��L�} ���ʒ��;�&~��  �ƌ�����Ԭp��Rӓ�������3�Y��b���S�xe�f        䯽���p�P���C��8J��uy:�Q������RZQA�l;L+�M|?9��t�>s����_D��L�/�70p���\�+� kr��"�p{`;+Kq������cz?��W�N� ���m�9���yt�W�)��iHw�����9l�h��寴v�\�Nz΀����?n�g�q��g�4��l,�>$�;�&>��Ѣ�q�u��>%��q)�B����bn�5f�**_�R�S�h��b9 h?m����T}�E{��x���S�aF�p���ފ ����l�ɑ���}  ީ֜p����T���hDeB/o���掷�c�ɍW==\��a���C�%       t|j�>�]�+*��eto�������^�"�Żf��z�l2��W�dW~�b�����R�}��jW���G�]������*�ᾙ4�Ww���H��C��.��ߊX6���E*t+L5&25�f|���?r����aȥ̢{��H�sS�)k��p9�z�1?�ts���Oy������>�.^���]�[</�R����=0���p��U'�D���y��i��Ƕ���yq1m�Sq����eg��k��Ƌp�i@��M
�F� �#�}a�q�\وl�����RJMO2�P�J���x�Ye�ee������:�xM|~��I����U�t_y�"      @�V8�VP$���%1�zK�،��r�/��X����l��
�W�'bkia�nE�����РL����׫�t%��ֺ���绍��{o�[���ف6>z�h�{15�LAbM�`���_��s�'�r�Q�q���}�n;B �s�T^YI�h��Y����cĥ��;�;�-�K����HOMBONBc�h��K ���Bn*GG'q"BNNۄ��{����>�v�f/߇o  ��/_W�����i�%&�Ҙk��ǅ��/��v�����o[�P�� �[08Tێ      ��B<]iz���N�����Κ\�l�BcF�U��)�v�X�R2h��X�>�V�k(��[\���gH.-�@���kM�ۥ�Gg:�r��冼���]�5q]|���s���$s�ܰ��%�r������4w@Oўv�#��p߅��Hv��[?�suL�?�mB����|�+�d.uq�)��)�ݙd�_r����W��J��5�d��W���!n���֖TP�6� e��_ٰ���-�f(�އ���.���'.*~��@q����LI{��TNNN�kk��d/���Ra[��i�hG�3  0y=ܝ�Ρ��a��Y�����O]��|      ��.��_0�8m��qopYn�կ�V��HΠ7����������0�����֩�z�[�x��v*1M{}L�_����k�U�� �`��*_h�õ�S�_>�cH�ಊJ��C~|b(�w㣷Ӝ�ג�v\�׆P�֧I�>�-�o�|�[<�z{�����"R2��9P�������v!ٝNJ�>~>�yw�#����tcD��pxo΀���a7�]��9��I���Ϗ��ꡌ8���`��Ej���d	��8���Z�-����6��mwuv� @��;N4������ ����ԧ�?���ծ.>SswT-?I�E�Pi��     0���'XqX���B
JJ���\�����M�m��=7�6�������%�}�yK���$�Ԛִ\����Z��q�_�[�6�Q�޷�jwm�N+ϱA����3-Z߬�A����I6j�L�G��ۭ� cm�U���m��T�;<���mE%��6��̸���tѦujhw���J�қv�?-�P��]�x.���t���5��y@M���;����!��u���2��C���T�+Rևߗ��wJ\F��=�k�+nrP��{2�t����z2��?M	:Le�'|�hȬ��@������wɒ-ԧrttD/	!�  �� �Tj˅{�����kw���������c8�     `$X�ӿ'��@�^nden^��Jˤ��cE��s:U�dei�A��]���q��ݗ���+i"`��S BSj��\cF�����$B'{v���-a����Ь/~�I���bj��z?_�z�i�>^n��80��qZ^�!��V\VN�.�&���b4�&� �g+��j��9�pU{}Z� ��}���=�r�8������Ά>�7�dǡa|�>�G�����m�:��h��޴�Os���dÙ���t�/��_�:;t�n��Q]񵥯a>�Ԫ�ԑ�K�gW����O�����'���\�z�i �q���L��)VV�F]�U����� �'�     ��_��[��pw���|6&�`�ZSU�ĕ4��      ��+���ֱ4S�rWc8ĕ�����a��ޫ�Q�d�st=9i�6���^۸_��R���~7�	��f��c��У�ҧ�O��ִc��Z\un�2��c�RIF+O^4�z̕q�����zai�Amn�o���YY�p�g{N�j|��!=�f7��W�c�i�Vf�8&*������	�5g�Fێ7Q���$U�;z���g��*�3�N-�z�/�.4oP�hO�{e�_\jp��� ��3ɪ��&B�    �n��g^r>�ڼV�nށ��\�h��=2���v��      ��&��J���r���BFQY9��P^I��p�gk��`+Z���[��Pս��&e;O�� ���V��?[٬���{���d���B���$֋`_����M��s����l�y�B�W>,�s٘���n0RF�9��29�����RhS�\��~��<)��'�qظ����qC�K���}�I4�����foӢu�*��s�^#�_R��c��������-��UoSB�m���  �	�>    ����Oc��=���J�g���@L-;~�֝�,v@     ��uss���\�-W��H;.�Ӊ+���]}8���&�t'ky:ډ6�K�Ic��Y��P�]��ߥ��ϧ{N�����������jX~ʺ��嬆��q�9�W�2ʺ8�ǧ�B���Sj�h;ܺ�+�1n��\on9$�fsH����ߦ�hq1���AP�8\��B��   �}     5�@�ӻ���:E��g�B۳27��wot9n�YP$Z#s��e׹�g��=����e�����P���y4��m��(z�����҂�����-���\��e[���"?�7����)�>�u���V��.��09�
�n8M�~��     d��ͣ��>>��U;)��m���s�Ψqyk�!��m���Q���֚^�y�������A{�Pl�Q֩�_g{�: ��w�g+�3�ϵ~���E��z!N\���mGĥ��y~��Lu~���i��'��ِ����M3y�"���N'����  h+�    �!:#��\��÷��H�2_���m���Yc��]��_ۏ���1I�`����Ft����<���kl��h��U3���6��£��P���nr��C��C}     2�����}��V��*N��JV��-{�Y����uѭ��)e��[hʢ���	n�k������h*���L��>!�È �l�T�&�!�վ��)�s~��-�x�従��v�*�+^���}�Lb~��G��;�PO����kO_�/�����b   cA� :މUTVA�A��@s��V���c��9+�dg���++1l�N�f���y��Q�9�e�jZs����v8.���_ڈ��9�0m8�󠻿�(�b��k6����c|�0�Ӎ.�f6z�1�~z߇�����&B��z�Pw�C     �����������t��i�9��D���ڒ��9���V�s�ק�v��F��79���zJ�
A۰S^�o�C7��A����b2���.~xa�zb�`�^�e쬪�w�2��c~;[��=�w��M6���`zv�0zd� zq�^���y2zv�Y�H|
�O�֤�s����2���U� ��!� �F^q�� @��2J��4��-O1u���ʊ�t%�
��Դb�,��6�lW���S�kxG6)i%��W̯i��)V��$}�z��
l|���#���Y���HZ~,R����U�f~���m<_^���E�'�!ݮW��
�L����JV%d�R77'��� ���:��W�� ��n����A׃})9��(�e�v6������uuu�q�Տ�϶�U����!    ��<l��c�5?X�+�Z��ze�?W���)��?o���?O$N8:����}}��K3F���h؎���YPl��W��=��j��ǒ��
�޿,��6����m�I��ϱ�.�*B�*��dњ�kkeI���!�~�=O-��۸��?����ҍ>�7Y�?�u���`����˯_���5}~�����)��[%w!�G���fO���Ҋ
��S@9�%d��ǡ?og{�2�~¯����:��� }+m�1.{`�x���ȉ-o�:�d��}#fР���1��t,�* @�B�   �p���0W�f��*��Ǖ�L3�ǡ���\��������wL�b؍C}e�9d�*�oS�J?G�?(��O�#���z�(zy�H:���@�NFQ~	B�2��I|��+,�?{�>�c2�aD���K&�?ruB�\-O���]=��E����Sq����1�o�o�i���G��~����c�����ҫ�������sho����p�C�    ��]T��������)<o'���/,!�pe���Na�����s�l�*&q��OJ�
I6j�����gZ� 1'�e�Q�P:�X��g���F�����&�p��ȫר����|p�$��?����!N�k��o3Ǌߙ��Ͼ�o?*d������4�ϯ�M�9�B����� ?֏�M���2�|�dc8��[�ѽ������mGh�Q���M�N��G�/7���r�(�Ә���ڽ$���)z�_ޯ6�OZ�b�����[�����a~e�f7��7��q������:y�N%�QI���7����[�+��0qR8{i�H:��F�\���ȋӇ�P㪪��(��'9?�t3z��4��3S�ҝ��H  к�   ����T��kj�O��KLny�����P_5u�Uʵ$oK$e��G��ӧ{N��n����a��+�F���[��ӆ�Ѩ�'>���_w�e�B���m�u�2��uZD�N�7�;�+�7���yC�{k��b�)�Gyn�N1���;:�yp7om�?�a;C�N��D��Ά�+�7FD7x~,����c�IC    @v\����Zh4"4�۹hji�$>i�q� !���Z��U��{��^�Ÿ?H\.�g���񙹔�[ ?�w��"+y:�S7WG�ՋB=����v.�~<r��}���}O�Ioo=,�14�2?7����(��l��2Q1�����\c&��~�zG�'�O�[���P<2���\J=�|;�NJ#Yk~��l��h�2�/�)N�����{G���������E�e�IJ'Y�޹��뗫�u��忙�.�"���t�w�"��a1��Ý��;��}v�.�T8��塞@��.��0�}��b�����빚#��<M�����  ��   @H�(mf�O��K�'�57ԧ���'�?���T<^�_3�5����/.�Z0��;���t?�
o�����ف�������g���u��KԻϘ@��}�S�y|��/\��wtr��^^�t��z�ۆ���>����x$�0m����a���V����Y\窒<n�    �pž��	-x��I���}T�Hu������h��x�y��U]����m�Gu?c{��KSq�!>٩J�lA�RU3\A�chF���/ۛT�����I��'nqŤ�㴩6���J��O_,�F!��b�	��&e���?W��[M�:5����|�Izs�!��շc����Ub~��_~lol
�M�b~���m��jfU~�UU���s�Aq]V�������5�����������b�A����W��e#|������'m��je|�,e�;��@�ϥq���}8Wz�r!�d�'�s%F����-^�Y�`og��$  h=�   �����}���.��Q%�����l�M�P!�
��r���g]�0���;v��+_�-Ţ�������r�Ν@OL,ڧ.=r�(�:�y�%g�}��;]\��wܩgL�N8�R��t���״�=�|�`�ܿ�`���:��܄�ˎ]��;J��Se,�E�.��>����\���2    0on9$*Aq�7����p~T>_q��tbz�a�2�'c��{��i�q|�n>D��v�y�8��'�p�q݊ߍ��.������t$>����~o'{z����J���t�������Vnw�s!W����t15�dv,�*���gQݍ�C����Õ�տ8�[{|\�����D�,���̯O'�_~��>XF/N���Q�/?/�uq���c�O]�]�_�����~�u�U6M���t�ZlJ�O��B�Z����p��=q[�`ߐn^�+�$�'�����}��7n`W/�  Z�}   @e����J�EiYY�oi�߶y��8C��-�hV� Ѫ���hjNO�����+i��D�hQPԌ
�|%��Y[�����rH���%�Į���`��h5�w�u�������N�a:m|�`���:���$Q��n�B_��o�[[�������@     ��Tb=�z7}p�$���~0�W�涴�y��-��A��p�#g{������U�L"l���)n��U�{y�Q��+��ۈj;vVT�|�/()���q2Fݧ|F�	=r���G�����8�j�t��硭�usX�8�u2 Wq{�V�3����v�mM��M���jVj��?���..z��>�����7S�������:~��_�9��ˁ��L�n���Jn�2�����������1�\}��S}��%^��3>6"�W|�m��:x4�+0@�zuP�t����5ʶ�u�}��S;�  @�A�    ��x����gZ88���Wo�Ơ����ҕ�����T�
n�p�쳶���|c�\>08��`�mΕ5��c��D��������y����nSq@otM��;���7�7�O�c�5�@     S���J�ɣ��L� � �}㠟_����p��5{hgT�>��B���i;�r��|�=>~�r�(q�ֈ ����7����'W�Ⰴ�p\
-Y����L�# ���O�N�/�P��T1�OK�+lr�T����P����ch��Ӏ���������;���N�����T_���L���|\���W���{9ډ�dq�n�ǥV8t��&  h]�    AJN�8���Q�a��CE�h�CU��:v�֮�7&Я�`�lj�yW��(!3W\�3�O^Ig���Pw�:�6���пkn����	�95�ϓz{���[����c��tN�    ����v�����>�oM�&���UX,�|�m��&UA:�����_�Y��EӨ������������	����s����v����t�'��s�������|��;�����T��ru�/�{~?��詽OG�_����%��R�a���t�_�!����=�V���M�߯;��r�>S|��kT�r<�j��Ǖ�U!^n���9̬-��X�����Qe ��!�    `D���['�嵍����!�hho2�]x�gbϮzDخ:�j�dd�P&W\d�x*��ã����V[mp;޺�}c��?-���Қ��3��T����S���1]\-rT�����ˎG    �)�v�kO_��h'Z��W���ճK+*D{ڌ�"���EWs��e8�.�n5�����#iɄ����(����%���;�U��)��l2uSB��'�'�U�䊔|��~W>4�~8A��a�^{mS�U�;��r����O!ߚ�*L�_e~����P��i?�u��������g~��ӊ����rº^���r����hZ��l{��\JN˷Ru�;�l�`�v1�v�'c�t��Yw1 @�B�    ���i�y�33�6�dcE��G/N�=�q���� ��D����C���\5@�n0o�j{�<T\�O_�;��s�����=Y{��`W���o�z�G��G�\�vGjeA    ���O�I��NKqŧ��c��N�l����t�W�	��U���NG�R��g�}v埽�a?���i���Ο��6k,�7���s*�'��V��?�d��x��{�ӿ���Ő)3d~�9p�䫸�5�9E%��2�������tsX��2��w����K��ו���;�������w̔����J{=������羊w�I��_��9Qw�����\��;����< �օ`    @�B�>�	��Bk�ջ�w�z8�ROOW��h�~�g���vO����z���6��[��T��y���;s9\�gj���Ew� /������ކW�����v��I!�h{d����w�]�C�      �O�O��I�������ߢuq����'&��,l��������BA�?����U'/Rf��VA��U�jU��q1�����j�N�-��\E�?����,Q��~�<~��u����J�xb���rH���/�j�`Y��=���~�B���_�����zD���mu��`mI���@/L.�s���n����4�e{/'  �.�   LX��|[CU�N�
s��vks�Ҽsl�Uh:�8�x��Pn�k��lz���E�������ⶻ��>�`�������<�9��N�=�c���A��Ҵ?S��o�M��������"��A�m/     \7�����J2� š��Ր��{sp�ӏ�O�~. �����;s'hO.c�Bz��+t��Q���ޓ�3Ʈ��ڸ��_g��T����tr���'=ru���Z�w��@?����)��Vq��}k�8��O�Μ	�pH�����M�:#����X��������	V'l������E:�k
�_M+�V�Hض��H�s����h#������	���/YTVN��� hm8�
  `�)�+�<S;pxC� 4J\��@ιW�9;�:�J�9E�#��%��l�*)�����F���.\�F?>G�+��Ҳ����MWs���L���^'�����P9��>66�O?ا�>މv1��Ĳc������a�b��h�6��ug.7:n     Y}�h�c�!J4R{7�� ����$���|�t���y�EKC���Cp㟷�����j������~�@<�<��gO��.u�:r�>[0ET��e�?x��~���ݢ���$��ߦ7>����ʝ�j���;�s銨r�noK^��ۜ.?I/��K�Pݭ�����9�l�T�5����I+���Qm����@��le~/�*B`�)���8�:��G/�K���1���wL�%U[�1q�պ�W�^g*��ߏ_��o���*���=���6��U_����_��&0�]YE%}���y�8������C��������̯]���7�v��:���*e[��nk�l�5�  ��$�~�k��)��{��<�.ڛb�FR���s�:�]�3����w V��.��J�#�w�p����������4��l�	�۸nnq	������&�4�I�;����|��ܜJ+*������z���$�c�������='�un<���6� li[�k9t06I�������Bh��(��_�v��Gц    L�Đn4{@Ozg�a�d�	Q�����G5-A�4����k��r��y�^����O��[�]|��Ǖ�ߨU��0�o
כ�]Q	�z��g�ի^ǟ��]�[���a>��P=^ݰ�~8a�g�5�/����|�%,P��U��b���m��	rV�4t~w_�B�Ly~}ݵ�/>����{E�P�����/�Ǳ����ɡ����m��W�HF͙��F��V��OϬ�%���tћ�W����3��<���E_u~��Ĥ�������ɼNv�=p��0"�zy�Q���?s��:�G�����ʆ���yjhwzw�D���,nK�+��w' c������b*)�3�A7;;;2oQQ�����T����	�!�_   hT����S���p�ڡ>��4܇P�DjnA�[S��N���҂u���q)7�£���M+xG�7ט��� r���F<�mxuqˌ�5��;��"�ajw"�g��    �)��rSL��UT���մP����5{��= �mt�����i��b�4
�⢭�7�oP���j�X\^Aoo9D��9!�X;��k�D��P�[�6�q�������)�:Ws�����_ �J�2��;����]��(~o\͵����n�R��_�L�D�ߝ5�Ԍ���ɢo7�0��&]��W]Uy~�T氮*�uͯ�������~S��o]�;��7���@y��W�]����m����_�9]lKl����W�RBf�8q��!x;�Oy��E�{P��m���\��|����GIII҅�8ԗ��g�`W�������D��}TXX�`�dp$  ���P�B}���/ԧ�y��Z�(�A�䲿V`ol�����xttFv���*�b����8 �-jN\I�����h��֞�L�Ι Z`��%/���?=�⪀     �������)��	3\���3w��mܯ�nX�/��zݖ�����%�l'��c������1�x� q�W�;��=z���j	y4�*�y�v�sI&�f����Y�=��}~�Zy�b���/�ܚ�������_Ϯ�E�$���WRF�u�x���3)���(��OL-�et[����=����˭K�0��-.�'W�lR�����{����x��/�~�o��{����_�G6z_���<�s'ҼA���ܚ�b��QC����m�:����,��vV	��t뗿��s�+�1_>4�=D�Z�Z�Y�1��q�O����k-����P�GS  :��3 ԧ���B}��:H��>�UTZ��1�Ys�oL��������M�>6V�?�t��;�/\�f�Ǜ_R*ڸ,�[�S�`���_8�      �����b��E�)�ӕk��-ҋ�e;��s�M]-���[�L�"��vm���V|R��q����L�b<��o>H_�;E��'>K����˯���Vn��O�i��hz�����W����П~�bP��-m��6���J�o։���$���|>V���:�)󻡎�]�l�A��ďӘ�����YK��G%e$��/�zx)��ee~'���<�}��K6�#�?�w(����~T����MBV^�,�;)XQiY4�_�#����{YC�]��S�ĉMy- 4�,a7nG[P�O�M��"�'7qDu���]lmm��De{��I'�WRUQ�o0f����F��%4�Ñ����M���3J).������<L:�ׄP�ʔ�}����˛x��>��/�A�Ft�!Ks�^Ž���q0&Y�f��|�I���WY�K�q;^����Hq�r    ��q����L/�IK&��F���g�w��Ov��۾��%&W���/��Rz���4⽟�o��j������[�b�8Hr�-.ի��>	W>�}8o2��$ns���΀_�-�ݵ6c��wLU��y;���8K�2��r�E�ߤ?������A9��/��i_^�����(�*���M�vd�шex�2
��TbT~W�NE�� m���nm�S��xꓟ8�jkk;����;0�>����u�i�����=Z���s�t�3R7�g�/q8��L2�׌P�J��. ��T2M�i�g��>�������-iHW/�`^#�����K���;�^�Yk�6�*5�PS��q�    ��(.��76��jg_,�FA]\���BT�ѧ����լ��!�=�ޯ�J_���P�����yҠ��z?[�l�?��ߔ��ѝMN����h��F��Et�w���]��O����/���W�2��M�i����{�W�wH/zg��ld�߳�F�߅�_�W�z�iqQq��\���b�&���
��u�O�^㭪�D����*  @eR���T1=G�L����>��M,܇P��}��w����q��ƪ|����k9�-���=��_W���}�sm�g+�Zfp�    ���+Ӎ�p�m�XQ%�̌D���YDe��jg�]v��DZ�rG��d=�Wwт���Ʈ/����W6쓲�%p�+����@��KW�׹sW�
R�LF;/&п�O�LZe~�G��=�ߥs����>������B�t��Υ~����N8��"㤮���� Y�uح���]B}*oRR����ɿǡ����/GW  :0��!ԧ2�p_KC}���H��>0%S�QF~��u��"�q5?C�R�v�=j*�ݦS1$���Uv
s�    �3���3�wц��鳅S���Q�P�**+��E�)r����g���T\U�[BN�.*�s��[���?��ѩ[
ʪ��;�� ��8qQt�1^���%+5Ч����@�i���S:����/u~9�%�^��ބ�m���˭� ����}���o�������$܇P�i�V  �N�p�C}*��}�
�i�'y���."�&����M��4|�������&�]�z�p��1I�Y     -gomE���7����9p�䷻�����M&��l<�'W�a�����9g.���O$w{[
��B����?��}���)�F�Cq)>�Wn��VL�ʣҊ���@ߋ�GД��$���&�� 1��B����yh��0����}A���&0��e�l� �o������Ӂ�d�VPD���2��>b�|�_|"�l Ж8�v��e**j�ך��e�U�3���/]�t���[�fee���cS���   ����V��d�U9ԧR�}��n#�Ry*wq�/��t*G�LLxt�^�>�~�vC�μ��G�    ��ۻs'�C������Muվ���ipW/Z�b;�t�L���5�u�Q�O�STB�o
��E�-���%q`��;&�̾A��}��6�{Lp�б�	���с~di��q��LR:���(m���[>��E<������Fy�o>K �q�����__��T�oE�:�G�s1zˇx����9,P�v����Q�ݤ26ȟ��6\��W_��oOe~g��[�_~�n��"cs�9��{z9�����\~���~����Q���o�2�<��c��k� 73ec7''G��ZCHHYX��,��r��5������<���H+  @'!U��C}*��}�l�P���}���I�C�Lپ:*�q{ދi��?&#��������}�e�     ����}4o��v6�۞Y��u��O�O:���s�ϞZ��d8��?��5w���s2���E]��
���6��oϞ@N6V��͉��i.���D�>h&^��U��U��?��������C�c�5lky}?Rye%�:E�+�\J�"������O�Z�K�3�~�������wT��!��������<qQ,s9=�@���������_�M~7<r��r��1,��)��]��ICD8�.���{X��ۅf~���KZ�]hsqu_]�xG���.\��O)�}����3�z����w�  	��  t"�+�wk���y�^Th������<2�HS޾.�����ʎZ���H�Q���������`T�C���~�A���;�t�-��kJ7���n&��|DJ���?������_%c�3��j&)���    �[zo�D�3���6�>f�.Zw������4�_K�����#{��_~�E�ת,$#�P_nq)��q�U�������b�Vp ����O3z�0��`�8���'�����h�x��箺8����x$}���^�!�K?zw�Djdz�՛Fі�4����$���J_<��r���!��66��(��-��hhw/���:��<Nq��~��lhT�����b|��>n1̕�tq�-);_�P`ge)n��I��4�^Z��d�U�y��m��k0�7R����߿_�1�^^���xx{��ƚJ����Q\Vn����������(%��
Kq��)�W  �N&�Տ:��.�Yp�/�3� :n��7L��
�nYu>ݵ�xw\Dk    0���[[�m�U�㖵|;����W��˲f�mk�e��x����;));�I���ǝ��@���K��u�8h��?Q~���� ��ӓ��UMk7�����h]Z^A=���C����A�"`��m�hhwom(���ϭ�#*ნ��2Lۚ���me~�&���۟�
s����4<�G;��n��5��|uf�L��_־��v~�������5{�~}~��̯�r�����^y"��e_�i�v��zZ٦�E��̕
�L$�ʼ̃���;��B���N�J{lE�˕�^�K�G��K�GV�WyN��������՛�z�M}i��7���F�3n{|.%�V��(N��+nZ����{�ʚ�B���N�Y~��Wֽ3*���w�$�`           H�?w��յ�"z~���TT���r!��}�3}8o2��$n� �~r�Nڪ�\Fy%���C���&U���ヾ|���SE{A��ā�[j^w6���
Jש���WH�b�)-���0H��d|��k����ȋ!\�%��+�R�7�x~9������46��=����ջ�ۃg	���{sX���"�w�^�����_H���7����Ӛ�~�+����i}������O�:���׃q\M�ۊ���ң��E�=r�B��7p�ݕ���K���*�*�ێ����<���*���0��f��%�[%�Ø<w|�Ә��O��H|�A��uv���N���t���с~����X  y!�           ��=��)"ZT��vd�� �=�m��Cz�;s&��>����D�����f�g+�-���K��^C��ж&h���Eȃ}���^�O�;��Cc�k��o��/̧����g{N��t���=8���r�?7B����q�>��뷾�I\��Q���r(��B}���N|M��m��爛ݴ�����"�_��v�+bq�Zق}����i��WuS�y��x�\��}����:�E��y�Z�n+�W���TJ�-P~��ݛ��
�g�ļv����t8��p��6>z�����++it��*N&��̼�� ?� @~�          �T�����E���
3���y��U�f�	�gV�t��Sq�/���5�/���9����h���Y���$���3I��.�[\Jq����]��j�>�q)"T#���餴z�������ÕJ�+�������ߐ�?��������o�g��rOS��&��[��r�}��ם�\oU]�hȡ��..�"�.����x{\��F�����c��ה$e�p�G�չ=ȡ��%�)�YY������~a��pp�����r,�*=�|E�eݰ��̌F*s��� ��}            ���cE��h��w}���Fo�6�:���u}��T�`�����:W�lHBV��%g�S^q)�:c�/�6�-��ds}~�(���9���(��[���{~~���9ؗd���jg#�V��R�歽έ���g�s��"�p�bV��x�_��ƛ�/�cN5놦{�Qzty�2/U�.�-r����?s�����B��띟�cҠ������t����z_�|"ȁ�$ �!�           �xj�N������p��t�^�>�:�.u��ޢ�!@[�*A�Ҋ��#\��]+(&0��-�hpY������ḫ�o���k����r���ű�e<l���E�gQCr��[ܪm�eRd�xݯ��rzv��T[�Z�k�碁}����R"M��]|?�ϣ�`�^2a���ۿKV젎� �           @"]]�\����2Qu���أ˷QG��LOM"�r5%��p�J�6�a\	�a���'�^�Oj^uE[n!��M�������w��t��U]m�� �JX�4�f[��š���/?G�Us�k�T9��]rJhw�9]�V�P\2�J��m: ��     @j�����!��dO     о��Jh��h:�p����mK��nɻ������VN9��~/�M&�0�������v(��S�}Eu��C�C7,s[�`����Ҳ ��jw��"o����ab�������o� �uC��E��vD=��<UZ='����^��\���,�5�`mE��%�� 9!�     ��k�/�&v>     ���8���z���v���u�T>������hmE�����M+�_�#�)7,��_�i�W>;�Rd'��@{xht?�-���YpM ���NRí�QyH���`{G5����`���J�3I�r�����@65����Lu~?C%���^�e4OH����� ����`ߚӗ\�������H۫����)�[=�7f*�r�"�3�?��	2�9��x��9I=ގ��_�����4�mH����b�Տ�F!�n��n���N��\����F�^ !�}����*-/�rM�<àgV  @�noK͛�P    �d8?�������X���|�;}��x�@��ϣI!��Q�����u{���z����3ǐ�����[/��{ۏ��� ����CZ��ő�P�Íya��$���a-�o��敔�}�xf�q�7��L����/U��4f�h)�����b��P���hëV�����h�[���e|��6�?9'B�<ޝO.�a�����s�J�뻥O��Sxonu�w�(��O�o�[��_Ee%�zr��q�[�������<8����F:��9���������� ���K� _�J�Rr��  Ӹ`���$     ���' �>#yz�0zd��zο��cPbv}��}x�d�d_��9�����"�  4쯿����"��-jo�	��8H�⺽��.]0$T|-�����rV�}c��G����=����ZR^�m�V6g@OQə����ջ����q���^�b�4���Je���T��J�����CTy���UU�=2�&~���� ��x           ډ��=?m���+Yy���%J��#;�س+���+~�d�`�ZM7�Ǖ�^ݰ�Υd@{9�}��x�����w>��������֜_Y����ѭ_��OLѫ����Ϯ��h��	���ݼ�u��������ق�u�����skv����*�z��;/�Sa��������j+9s����/yk+����*,���^{��P~��[<���:���5}<o2��z���     )�(v�j    �|�ZȖ�q-7oP��-���7Qqy���oo=,ڥ}p�$|e�(q;��\��V��"���a�:.� `�qq��t'l�y������F���.B�^��X�pv9=K�=�)*it\��M�����D�� ^��Q�oB3���+�x�^�{��,̧���9����:N�<[��]^VY!�1�^^����혌lz�ʹ���E ���<	-y�`     H�w�=�j'}�pY�k     ����zmx�dd���Z\VN���M/ԧ⃹7�Ҵ^��AXn��UX�ħ   4_��k����Ǌ�)����B'��	�r���璛�����g������aeW��j}�N^�wY�~<�Dc����S��K� �`     Hkŉ���������=    @��.*��g��X��V��,4�"�X*��(���d��*��T>�p5��l�'�}���I����rdm�͗UP����2u_�h5
 m$���h���`+�_v�=�f�8��1���Z��/����0��zy� ��>     �ZTZ�h=     �W���b��/1;����$g[+�56#����r�������Pըc㶕|��i�2�[1� І��9цG�jOn_u2���b�81�������~�����S�
��]mm �`           @;�4�n��S\��r\�E��[@    `��\i�#���lݙ��Ȳ�TQiX��q;���uK�F�����^/*+' ��}            &�)z   @N\�o�#s�����~SD4=�t3�WVRSl���''׃=\]>��]{��Z���           �l��6���Vf     ������-�KA]\������?n���������$J�+$/G;
�t�P/7���Y��V4�o�����	 �`           H�+�趟��l�(�ݹޟ�8��]ohYV^Q�
,    r��P��"��v\���~��J+*��>�������Μ	dfF���o��䟽�����Z|���K�#�Hv����*붳����>s�����x����            �������!�{�M�.�j���   �\>_8��Դ�����E"�ט3I�����u��o_4�7��I{v�UϦ��~�N&��#̧=?u8��?X,�Ŭ�_��Y�R^^������PNN� ??�ƛ��7��4 �     zv/t&My�������pڒq�**+�?�7��܊����ҁڃF��^�;�?��7>��r+����           Z�������̌�e��6���7���E߮�M�ͣ`�г��p��/:�ɹ2�k����2�[YY��wr������>1��x��JyNp��`     ��4G�믬��J�ÿ6��7�2�.�;$�ܩ����i����     ���d�Qa���%��    t�y�4��e��M#�a}D�]�O���I�-{w_J�n>D'����8�WZZ�f���̔�Svv�T�k�P��ٹ:̈p���     ��]���(r�*�Jss*Qn� ���m�L!v^doaM      P�)��B    �y��le���Oyy�>zc�і��ف��5��WH��(���d�֡>�������ᾶ�LX�}��>    �66�����~��r"E�e���H�O��B���^|_EfTa��J�9���Z�)����m           жJ+*�p\
���
��8�Ǎ�rr�&����E�O~�    ��[��)ô�/Y�ä�}̬���u�"��
�
�B�TV�O�daiC2����WE            �������+��v�O��"�'7�     ����2Ң��JCs+��s%Gw�h4���
rc	     �7��d�|~(*m�vT     ��d	��Z;�'�x��}     `Ts�8{SEy���QYQ
�姒��/�;���c*ȉ���p     �]��#     �


�
��8�gff�uVUUI�Sq���4���     �2#Y�vQ>�V ,/ͧ��t*�O&3�9��9��c*.L�i�           2��[Y������mD�X���Q�-�`     4���3Yڸ��ƒ4+Ҙ�WK�z���\oY+q�X�PAnYZX���          @��قdU�A �     M��H�M����UU�Svf<�{�FcN             p#�     ���:�See,]K�&w� ��             �`     4YsKś����S UU^���K���I��dV�wp�             tf�    @�23Ӑ�K0ir� �
U��������i���}vvv            �� �     m��}��=��:��s�[*��ы��D?+�\ii)            t6�    @�1�r kW��s%+�kʕӜ�#߮D�            �3B�     �L�]nK��[�K�q����,�˨�����8�            0E�    �,��H�� sM%搽�            tF�    �$��ͳ/�e�QvFYZ�Rn�G            �|p�     �anaM�n�TQA�����=�ll            �3A�     �������m�1'W��D���EN�����    @�f����n^49�;�z�Q{[r�����*�*,���<:��J��)25������%M��;���ő<l�m�E��WHg�3h��X:����u{;����7�~�J*%d�6y}�8�l��n��[@�b���-a�dea�w��@LR������{���"b��������/�̕�d9E%�+*�����`rS�_���ٻ�6���?I�{��މ3�	$� a�U�
��-��P
t���.�-�B[F��a��Cv���޲���s$d��Z����Нtz�;�9�������z��vƈu�3�g��<�j��ŏwΨ��v�>�<���׋q8t��A���~�1����=j���t�q^�X�m������t _�a���O^Mm�q���J��Q0|�}���X��q1:ճ�^;�
�bׁV�i��3=�hλ��e'%��9r�Ku�s�/����n��5�O�d�ֹ���W�@���x��2�[*��   �}    ��|��t:�Ŧ���l[�ּ����Y�	   @ג��M�O��&׽l��҄��t��,�`�xZ"�3���8N�?Jq��o�f��;Κ����o|�7�nm�'�>��]�^ߝ�ZÄ�^��kV̟	)�~ln���ۥ���*��s��Z(���ӭ�W}��������3]��	@�x_�}������{���	��}��������Ԓ/Z�x�\v�4����O_Y��zI�c���LH�V��bct�I��zj��f}�9֗��g�/.���cݫ_F����y����^������l������4�[����������z�&�ٗ��u��[<�9�~u�4�<�o���Rm ���0��m�����?���2�+��ooa����oUTר%Lx����[��Ǵ�`   � �    ���gWR�PE�Ta�N�޾\Y=r���    �L���.=ݪ�������8F7>����;�����y�Ӕ�L�ʟ�V��5�h�����SoY����k��/��*�Zj���G���*%.Ƴ��Z|���IV����gL֋�7�8|
��⃳O���	8��;����9�j���j�+&���3F��1���jO��E�ݦߜw�n�6�mk�Y�,��?m� �����������{y΋kO��,   �^�    D�؄,e�$��h�宗#*Qݲ+:�
Ng��ˊT�TMM�䮑ۚ\r�j�h�    "õSG��N��:^�;;����vi��|.���Մid�h��A��U51P:mX�&�}��ֽ�R�qLH�5[�Ά�V�ߒJ���tl�n:��:�tM��/�E�|E�mh�i�Jm_;v��_�����j��� ך`�e���g�i���F�oV(|g���k���OSEn���VpԴw=\Zn�z�y���T�u�@�7�o�Nڷ��>3�>���<B�^n8�g�/��jrlӶ���_�h6mn�i�۔�v�c��(�U�k�s�������MVu�=%�~6����oz��y�b�uOIԏ_^��
�^�Θ�����   4�`   ���JPJ�0�%䫴x�r������ԞJHJ���H��e��(�|R�%w�M4�   :�ӿ=������O�V����k�@�m�N�c�6[��T�{��u�3�_�����׹~cn�nݭ���j?{��~}�jA��ًמ��|A���gBR�{dZ�f�[�߷��~�}���R�LUkm�lSNv���N�O=R��Z�
�`��vt�͘��|�E��WWO>�jo�ϴS6���&Bz��������c��ZZ����!}�V�^&�:�g���q�t��\j�X���7�۴@�t׵�e�&�<�`������
��z�S���ժq���#o{��o�-�-��׏N��Gmn*6��_���M��T]������   ڃ`   �#&.]ѱiJL)Te��mSa��?ϻ�+d}�ɭk[    �랡������R�f^�B6_�;�o?=O�`���zf��*����?���Ea�w7�Й��7n����;�j���?TK� �gM�*�M�Ǫ$g*6�?T���/54;Mm�+�ت�f�<�K'�_>X������jEl���+��� طt�~M��Ú7��M�߿�Y؞��>��uC}����9��{P�<���|���j��&���o>�o�Y�w�,k9=!�j����(f�f�c�J+���_�jѶ�Mޯ���j��~����YV�>���p�}�ig��������c��OV�`��0   ��    t(6�M1�i֔�R%gU�*���������X   �8��d%�D�����������s@'?�r�3��W�N�L^/��ت
[&�7�����+U[��F��e�lgn���WT�7�ԩ��[�.?L�������Ǻx�0��K��s�����M�ϸ���>�`��5[U\�1Z���V��ڷ�7�4N��t�Q�C�T}����:S�-A��ru��X�oCݔ��X�7j�o��e�`�.�+,Q��$�:��(�>��P���w��l����k������[��|��%�j�=�V��բ1~�֧�{Å2�M{��N������   ��"�   �ò;b�Mnw��K��}ll�Z�H
   @���c���-o;\h�mڪ��J������Z��~-;M�͟�!���@�����q��u�?y���7[<ƳK�[�>�Tk.�w���J������+��&����� �i�;�o�V�:���&Du����N���RGaZ��{���W3&��s��&����{��=}�[�n�sk+s�4Pz���	����7Z�j�x.p��zӚٜ'��t�{����ie���-��х�tѸM�W[u�oz���ۄ~[���7��j��6�5�X�m�
�nAN  �H���84�9�   ���xEǤ��r��\�j   �x��6���#��*��5Ǐ��4LKܶ��4a�[gL�Bb�	�������ڭV(�TQ��N�BE����k7j��	d���Jw�_k��&�h2����C�W�����iWڑ�}f��	_M��?Z���'�=��h�*��y/{夯��.޾W;���>_����̦2�i�����=�`y��q��z`�2=}�9��s����߼�Hg�d��(�~v�q�ޜ�  ���rUUEfhtKHH�x���.W����A�   ��=3u�������m�T�A�[tl�5y�ݮ#?�����N   ��wJN?�|eu�\o+V/hj+��+7���c-�@���cVx�����SFY˦�Xc�>�&�=������3K���}����-TUMM����6�0TG�y�}�+����g��^]��A9yh_߲	���y�`�2N��ݷ<��ۘ�gU���n~����T��#�J���6yՆMw�y�y�)��Lݓk?�7,M�քo[b�g�}�mWm���p��o @����ݻwG\���r���$��>S/r��Ƴ���"�>    �n<q�5�։�=�5{
G���9be�L�p��8   �lC��}aü�ii��5L��}�
6WTi�����Z�y�/�gLԫUaA��7�w�ء��܏�`c}�On�ь϶����
S�ʹ=�����x�>b�UI�>Ӛ��#�H�jO 2�6�?��o�B���|h�r+�
ûgZ��k��!���U��
f����z-k�_����-MS�֧_�Q�:n@/�w��d��v�].k{M^��ܴL~{���q�;�����w�9_q���z+�s �EZ��������P"�>    m�p8�o�E"��v�U*   @�]��kS�`�chv�U��˄��[unٮ�:ˣ[ٚvɎ}�t �jś���#��z�+��Iu���7���3���Hy��  ��IDAT��8��`�	�ُ��;�{��L��*|�3϶#D�1�����9��3�g��[���6�U�Y�����N���qդ��ի[��{��HS1��3���nU��T|b�Z}�Hk����}�ky��  ��H	�;��)�[SS��2B}��`   b�.w�-�Z#X�b�)֞��:՞�v׸��L^&D)�o�z_Br�Fׯ�2L�   ���`f�)(��d$ԭ�+ ��+��
�y��T[Z�����γ�Z�&@W?�g������i����
$�3-iMp��m8\Z��l��~mxM�ގlg^��\�V7	_}��!�دG�m�)���;H�z}���WsN���*����:�����1C��W���`k��;�w��|�;F��-����X��bc�sǜ۳}Y  �i&�g�UV�rwK�ݡ	�y�;�G�/��   B잷[S������W�K   �@JO���\T��R��?N�?4�q���Sr\��ܖ �s�6�3�X��N��jK�[\���I#}���6�&̴p�M�Ǫ�v����U�ۧ�m��5ʪ�ze�utzo���_�b�����q����o�k|�m���z�~���K����}O/�� gZ����Vz��C%�z�����铭哇��I�ɴ�  M�ݻwX�}&�WR�P�W��}��:�}         ���~dQQ]�ǉ��8U��n�;�}�>�-&(֚B��
K���:uXE��V�ؿ�����[�>�4pmx�=�t��3��4�N��ʉ_����ZÄ����*��I��)9����h��>nBL�c�2HǺ?S���|˦�ce#Ǿ	��웬��ʂWM>&b�}�8�+�u&��-X�kO���y�T��e��Ԁ �N%��p���B�#��q�        aW�JVrlLP�~%�Ę�<N�_�0�-m	�v�&�g����`�����B�& �`Kp�~��ޟ/��*؍퓭�=3�n�a+�d��׳���?\�oO=����sNЩn������c��e�[���,�����^Z�Q7�8�Z6m�s�ӵ�@�"�Q�s �eJ\�1
�+�4�yn���\�>w��<�_w�s�`���%�  @��}��y�*�G��c!�        ®�^ة~�܀=NYݐNj|��@�B_\�÷�_ֶ ��k�Z�/��{g阞��žCV��˴�5����b��ɵ��.?\w��U-01��j��eoga�W��\�:�߷��>f��b�*TǺ?�V��jɎ}M������`�a�����T��~�.���em����~앚d-��)zkݗA;� �lL�oӦM*//�������l�k�`0�`noLL���B���C�        �]nqY��A�҂�8J�~H�����1�w�;F�mi����o�f}s�(k������U:�H{\#Xmx��Y��`߄���[���I~�����Վrv��t��j�����?���z	_�1�x�b����18HǺ��~=��/,���~[���*5�R��~3oQ���ۗ��`{�Ygy_Q�+ژ��|w��xƑ�3���� �� �U��v�йi���A;''GQ~_Љ���ڲeKP�6,GGdm/�F�        ���������g���d�q�.С�ruK�����Ȱ*� N[����%ۛ������f��rg��Gv�g�q7n;����Z�f��GJ��q�(M�ۺ��|��k��J��k?�J�i��TIG�ŕ�oUf~��_�ȴ�}{��1Kw쯳<�op�u/oP��'�O���0ǂi����$��̭�<6 �7&��{>/�����xj����q�����8^�]�I��5 N���r�,E���� �D�        @ؙ�ݖC��U~������V��@2��w��̑�e��~z�/�<�٣�Y^�mo��2-R7ȷB@��	����ۂ4��������ߝ?����ڣ�����H�o���+(L봧������z���8�
_U�>|���D�=�q@f��l*ę
C��@3!���d�+'���`��]���(�H�i�{+!&�j+�	q:~`/�r��Z�vl�s4U��gz���ֲ�����G鑅� ���5�{�+1�K���QZ|�*=�������҉a*vONT���E�oenQ�U@�B�        D�w�m�Гj�}�J�׏���[��y{�6_�ϸz��6�Le�����-WTi��=�z~&Xw��S���#��̇��[�I�`��gg���Z��6�����K��iu�-31����kwA`���.�~7o�;�ꗑ�oM	^�����uô1ּ����c�T���b��@8똁��?\Z�Ha΋��춪	I�1�5fH�[�^>iD�c��;�|y�&���	�;�Z����z* � �����7^�lk{�>P9���j���֙#ir�JO���fB�_�;��oԓ�ת���;v��9~���K�~U�͘���K+6�_��i՘ `        ��,\�N�k�v�	��ا����4��3g�F�u�	J�����9P��i��m�_�7��*�h퇯y~��r�+�����/UT�`M�DN�>���:S�U[�=�ҝ�u�߸�1�x�����k,�޾6��^^�Y?�1A���_�vꤠ���x���:��3�~����-.��*{^&t:���٪j=���=ߚ7U�.�q���<o����i�����V��5L%�[O�X线-X��h*a���O}�҄S�7}��JSq �*o�ݖ��.{�5}y�@��W�N��'���K�:��7��"���~KKw�orLS��T����J�1G��fM�5��O���{�W�@��        ����r�f�f-���×��K�+g����M��]C�ҏ
��������!���%��_hUx�I#t���eS=,�'S��T��V�2L�+���ɪ:��l���.y���w�I#[��/�f�߸S��r���7�
_�V��=q����4��f�.3�Z6���}��x�u�z`kM��S�2��Ҋ��:��H�Z�z��fk�[�}�i�����$^9yd��LU��y~���iq|��'��//h��w���6LK�@G��<�O�ܣ��j&7�4^~�L ��ii�]o�ϼ���Z�7�g*�.�u@+v�Z�rv�&��Ӈ��x����7\�Y���%;�w���Ϩ�3m�o��y}]dU4_\���;>:J�Ӓ����t��������       ����W�A���9���7��7�z������M��/:E�{{q�����%:��A�0����u�t�^Uaye��q��!��%�ֹ��s?֞ ������+�L�L��`�.m:����ږ˦�eG��ϛo�jBp���2��2�p��>��᫛O���֬���?Ԕ�����3F��q����<+$��X�z�1��'��7>�s����_M��[�M�д����ڶ�&0�w�V�9�Ha��}�]�}�%�v�V�4��T(�ͼEV������_.>�NHׄX�7罀?׻���z��	�^wd� Z�#����k��>]��,�B��ӳ����VP�T�3_v1A��� 0�_���O<��m ����+�
�浇�R��=�s�x}� D.�}         b�U��ϼ�Wn�@qGU���ҟ\m��LE��BO&�s ����)V����1��<�;7_bU.1�}>��U��k���[�h>5mrM�S��i���lUDӼ-IMX��٧�Gr�՞���rq���iCg���	s�U/�(�j�<��U��
9�z���^w�b��&l���W����1�Ա~��>��YS4�o��n7�>�6����G[�j��}ƕ�Gh�ˑ�3��ʵ����s���O�d'��G��<~@O�~�I�'�w�9Fo��Ai�h�}�[��WQ�T� �Ng����R��|�j\��Ͽ�wH���U-��
�8��fU��������i��h#�u7�?�_��X�]5�Z>�s?�}@d#�        "��m{u�#���ל�k�'-Y_z��h��lߧ��u��\&[g�g�j&�����:c5�y���=����?=���|-8Mp�_W�ԟ.��>85�TL���D����
��WA3�_�A7���^���hB|�9��6�n�Y��2A�|�G����R�	��-ͪ�g�2�3!�6������W�d*�z�eϱ~�U9�0-����5�y.[��pi�u�g%%�f�H3�{���JәJ�f��Wnj2<���oG^�u����;^[��V���>X��>��s,y�Qs�|t��V�ȥ���SPbU�땚d���&/���/������aK���EVu���G  ���>ccn^��3�~}�y�/�g����''��W��mr�~A��D6�}         ��V3���0�$�5r��:���7}Hkj��@�����_��jr��w������/������]��g�~m�	�����pY��>Q���~��E��㬩V��0�ܿjCL�ʴ�{b�ڠ>�P��m��9��XǺ��T*4Ǥ�qِ�*����R=���}r��u�yiŦ6??sl��b�U�0?'SY��U�i�p��,��ϟ�~~�=������1&<a*���s}���y�?L ���,����[X�On������Ws�]�o7��D6�}         "��/�O��q}�u��tJN?_�Ƭ�X�}�ު�w���E���p�U5��a����&4��G(�=뿾v�U!�PI��z&,f��k��fLЬ�C����τ(_\�Q�p����-��+Sτ&��n�&�׭�c}ݾ�z�s��Y��j��������^�k�����`�a��Fb��x�/����֔cu���;[�eLC�o�]�^O/Y�j�K�`*N��i� h^KC}�,�g�L��7��ִ���+���L�z�O��+ ��`        �h+v��Ͼm�sF��f}������8U���/���Q+v�*�3�V&d&�;n@O�]�	W%�D�pi���b�!m>�ߦ��Y�]i?�����o���G��oVXS[�}��9���kL�,�iU�K��QaE��J+� ��}[�J� ۳��1g��2�^{��v���g�Y��1=�)'��X7mz�5.�c�k�aϱ���u�7���R=~���f[�m&t����!7�]c�6��x�5e''hb�֥�\n�r��<�s��ֻ��3~��|kjslf��! �וC}}Ғ���^��oCL��T�3�]����=���zm�֣�3��u�Tk޼�0U����60���Qp���.�`        �L�7SI�L�d>�L
w�R�	��	���ڽ��	�c��&�  �xZ�����~��)r�k��.ٱOk�lp=�~��'_�s�<O=R��7α�Pb��b*`�/M���+&���,PQ]��}���xl��ݶ��n@]%�G�            ����f����[������o��p=���X�oO9Vg�`M��)���Z���Uu��J��           @D�꡾q}����V[�O?{�#��sP��-U'�~)�e�kFNm؟���T�j")D�.�#�           ���꡾czv������hk�/,���4{��'��/>�
�U9�ؒ5Z��7��J��q}�u��4 3U��?]����UO����R	��           @Xu�P���Wn�@	q��>]��{�f�7e`/=p�9�6.-���Ws��cB~�.\�'�>K3G����y���:�.�#�           ���꡾A����(+)�Z~�������nA��;Κb�����[|T�ϫܳ���;Z��k��맍�CVXU�������            ,�z��_F�g�/P��Dk���t���ՂT_bl���˷��_6�~Ay��߸C��Q�á�C���th�8�G�            !��C}�R�4���'-�Z~u���^����<2�}��L0����{�J|��0!��u�p�>            �TW��P�k7^�����k���g���j���N߼�&%�ƨ�����d&���+�^�P:a��`            B���������hp�4ky޺m��S��iy���/�P�g�H��Mܧ�v���~�卹�:�N�#�           ����>�{�������;�������V��r�����t�pk�3���WY����r�d�LM���i�}�t���6lXP�NHHPee�"Iff�GP�NLLPEEdmoPt�p�>            ]W�_v�F�̴�M0�`I��0�f�z�A=�h�Q��?�s]0v�U��4���u�;��M;���������N�Yc�����y�Z]!0�JJJ�`������P�������JKK��`)**�lo�:�N�#�           ��"�W+�H�\�n��#����ښ��6���9��KO��}�{d��_?ۺ���FqQGW�ۂ��g_(��P_UUU�'%%U6�ϡ� �a7��N�S����b]���       ��둒���i`f�l6  ��q���P��,۠å�-����za�F��wH?<u��5X�G�|�C}���*���~�"Y�B}^�ɵa�p��B����:�}         �&�練�;_)q1  @�sی�:�ї�žCͮK���3z1(��wX�zz��ٳ���'{^oǪ��i�0M+���
E�P�ܼ�����p���Zwz8�G�        �������O'�  ЁuK�׃�OՌ��iv�W	���i��|W�5u4�
�y�p���Jv�����T�p_�"�        B&';C���	   ���ݭj|��eM�7 #���	��(--k��+Tmj���"���            ���0����JE�`��"%��e�}��za!�HC�        �̦y�z���}   �i��\���|���	�uq�r���-R*֗��j�!�:P��`        �aэϽ���;_)q1  @�s��\7��~��ٕ_,t]N�Ӛ"U\\���K��n&���>�����noD� �>�}         ���ا�|J�����4��   "_��mU_��l���h�.";��mo�� �>�}         ����.     a��>�}             ��'��}�              ]S����             ����             tm�#�             @���             `DH��`              ^�#�             ��0���             P_�}�              hH��}�              hL�}�              hJ��}�              hN�}�              h����             �R!��             �5��#�             ]����fZ)��>�}             B*&&F��媪�R$2A���������r�(11Ih� ���            �>}�h���v3������L5�H�^�+--%��A��            �vs�\*--	�������>@��}�             �M��݂���%�p��            V���*����%�4
��            v�
��:����%�T��            BvW�ϫ�mo���p�>             #Ta7�;2Bn��^B}aЎp�>             ń�6mڤ������JE�޽{k˖-*++��111������R��#�             �i���A;''GQQE
�ͦ��+�Æ��ሜ��r��#�             @0�2�G�            ��(�2����*���kbl��''Z�(NkW Ђq.D�V���            !2{�0���]c�dkx��'�չ���R���㟮��M;[<n\t�n:i�.�0BC��|�WT鍵[��˴!7O@�ƹ�{��Ա��it�l�ꙩ���U{��+�Z�#�            ��#��!�����i�:w�`kzq�F�4�=UV�49��T���y�=�ے�bt���56G��4_�}�^@$��eg�aܹ��5����p4x{i�S��>�}            @�m>���{Z�r�dڐ�MOִ�}�?#�Z�qìෟ���8��z��_SNv��|��\�/Z�M�yJK��Ecs4uPo�y�p���_T�ZQ	�-�jz=�A�߹p��5�U�%���FC}��p�>             D��m-ܺ�
�5�T0��)u�YS�e����U�l��׿m�D_�o��B�������w�c���]gOխ����v��)��ǧUU�t@ �̹�ɗM���<Awz�_Ü����9�yEV`v��Z���U���sNP�j"�G�            ��Vlj���[���T��f�Q����>fP��>Ӫ��ic|˷��~�P�ׯ�Z�������ݪ�vŤzr�Z��ߕ͟���\��u���g{.�����*wV׹.=!N��p�>             ¼�n�/��+-��uN�_�ѵ�{�-�\��v둏W�W�i-��g��Q���6_��WjR����u(���            ����?TR��:���7A����~���l�:��R�cUX^) �U��υ2uZ��}�            �s�����{6������e;�79�	�m:����3��4�s����
�t��XW�=�N�/�G�            ���ލ����19��μ"��j�Q�yVӐ�4���Å͎��3�	�#zd�CD3���'��ZG���������p�� �            ���#�gj�5oZ��IK��!}4�H���.}l�ʝ�G�71&F	1Ѿ彅%�>�>�u�''
��υ�iI:iH_߹`����s��"�            ��w���IC�u���r���E��lC�A�Ę�����ʪ�����h��FϹpr#��o�-��o�R�>�`            A2�u�9'�GJ��}��5��։���W�r7�N}�5�yS��t���4��dc�BgE�            �+�|CQv�5o�z2Rt�ȁ���c�v�?=�8���M_���r��u�[��sxư�lG�S_����)�|�u��Y�\H���΅c=������>             J*�|���WX�E����Ek4��4 3U���O�G��s_���Fl���V�q�_E�J*�D��ʯ�g�s�OW��\h��sa�=��Ju�            ��3�Hߝ����E���'�?*�WR�T�˥�#Uβ���5%+)�7�WV! ���/�s.|�s.<�p��B�>�}            @����=�_T�)�Ꝗ�>�iwA��v��~�HC�Ҭes{s�>3�צy:�s�Wj�u���_gG�            �@�K˭0��#Խ݄���ѽ�� TcLe�czf����;,���s.��z�K�            @�9�6�:�����Y�y��>f�5Ґ>z�㕍�7�%�D[�������Q�Bi���}            @��9r���yӂ�@I�Q��ŗ�����l:m� ���iYڐ�'��Ϳ�j�����\��9r�K��            Bࢱ9zo��W6��������3|��.]/����v���U��q�v�q�I��So��tلּy�~�ZAzz�����UYY�H�����M�lo�"E�υ�74x.tF�            ��~�=8�T��~�>ٺG��TTQ%�SꙒhUܛ>���9Ъ�gl���,kt�߼�H����X}m�=y����ۋ��@��cct�a���Ӭv����)�,r^�)..��}f
���B*���}{Ͷ�m��5p.W:�r�=6����?ot�ѽ���)�ֹnHV�o~�g�?$h�
���3E"�}          ���w����q��}�֖�R��\��������6�M5.��j\���P�ʣ���ƭY�U��) �b�u����Ԝ�w�וO������m;\����M=��s���=Ě�=�S���:�J}�Z�	�9���e���j]�;�gB�������퍔p_k΅e;su��5y.��H�5Ǐj�v�����	�          '.Jr����Y��8��F����
�����<�K��ױɽ����3���T���E{V��m��꟟��*��0���%5�;w��\=�x��Y�N5����6�҉�=�ߝ?ݪ�g������*��]�9�6(ҙP_UU�B%��P���"%��υ���9�z΅�f΅/�BO/��E�BgB�          :�g����B{q���h5�Qx�#F���7.�n�/LZZY :��Vl�&�+w@F��''(3)A	q*����N��Vaye��6�K�k���핥�Dk�y�Z��:�P���L���;XPP��Ue��"!��ߕ��)���kk�*�UgA�          :��+4 ���{X��j�Tcs�e��e�R\T�2<�91 ���1��f
��%嚿i�:�p�����S��P��½�&�gBu�nC�s��#�          �T�#ں4��L;hw�����Jng��cR#2��r� �u�;��e�}&hVX�p_�lo���i�  @��yEm�	}Yj��&ב?4      2��wp�d������t%%g�f���i�6���| ��H	�y���V�V�/�p_�"�  :���B�[:W�\\Q1�r�eBx͈�L���rٴ�̡�8�b[�n{u�l�w�C���Vay�2�\J�ru{eu�>�]��j     t96�M��r��U�,Ue�>��WbR�RR���UE����.*�@WPZZQ!7/o�/��nwą��L��T*Dd!�   �rӄ4�K���mvG����R�|�C�%r��wg����^��7�-a��d��~����*)���z�ڴ�/�    �.*:.]�1�2���U%�*?���\�lJN�
���SuU�  ��	�9��ۡ+..�
�J�oo|||@��G�   @�\5��T��ڪwnվ�3��l���0]���$tW���      �d��X�=�=ZG�ui7�g�\��޿�ج��sH%E����U\Bx��	 ��Z��Mp���l   �z�$j�ȁA���R/��l͟1b�z�&�n[�c���;��1��5��k��}ڰ���E���J����U9�2����<�f��zŦiHB��b    @�x�n�6z�Gnrɶ��r�ɮ"��^쮩v�mQ��(w��J����-�p��96���}�@��'�Vb��V�'6���n�J�v�=X����   ��  �����.���7����}��j��_u�yE�z�3*�ly��I�{�kΕ�^;���R���*�J�-J��q�n��mw(����4E�    ᖶ{�5����ƩJ������������\�Sl�͐�}��v� E\B��š��ved��-   ��>    >޲[�/Z�oO=�Z�;Ϛ�����E���r��٧�B}��/����J�R����n�\ժ��Va�~%��� [��a䪩     4�nw���\���)����K���+�ӭ=fzD7�%6-Fgx���<�C����>r�����-JJ��9��б1�;��   Xx�  �.��Y���]�a��oz�o��ʩ�e��ooaI����D��~)��u'���5[���=͎�˙S4�{�o�٥����(6��]%*��R5.��UbR���3jo���<���     �Lu>��T������fE���>xKe���g>�#�]s��I�h�)Y �|q3!e�l�]*+ީ��2���[�%$�QTt�o�������'  @GG�   ]��;�k�=�nv���	�x׵����v�'�h��TV�{/���7\h��{���7ے״����q�eӂ��s?R84�����V���Y*ge�*J���䐲����jΪ"����ܮ    ��K��uwai�s��N�Aٟo���Iʭ��Ar���6�lI�nV�/��b�2��"�ۥ��ed���m6�����4;  �� �   ��i����5�֔��䍔�ͱۣe�L��DEǤX�u'�QuU�ʊw+��6ef���]5�r��    �Sn�=���y��?*U(���<��]�?z��Ꚛ�{ވ^- ����~����[�mPUe��zSll�   X�   ���kuJN?�L���j�{�Yu[�>�t]X[��^BRo+�gwx&{�5�P`�\���x�oQA�.�g�    ��s����5����BE���y����)���Y����-*oH� ��>�Ȝ[�)���_H  @��   B��ʩ��~�-yM�O�ۂ�s?V8�of�&d��>vG����(o��
r���]    ����[,���zqv�"\����K�ɣ�k�+��H Ħ��D�\%*-)Rjz�   X�   �0h�%oC-xM0�Z����*�ۮ�"��SZ    D ���l�����|u ������/I���J�{$�C �-%}��K��h���c�$   �>    L�j��P�w�oWGf�����UQ�.,/����Q��$!)C���_�%��.    @dp����r�,���M�l��{�������ٞ�I��.Q�	JN�jg��mQbJ_%&e   �A�   ��Z����ׂ7P�cS���Pi�N�]�;j+��t��|^��     r��Z宙�w����+��ֹi��?��͵�l��N6�e�\nTq�U;+���S   h?�}   @5Ԓ��k��iZ�6Īܗ1B%�U]]�ظT��&���P�iY�����r�    /�[+�q'�Y�l;��{o�(�����{�M�h1�7��$���w�J�����H�=rd��  ��#�   �Y���Q~��:Cކ�?��%f)**N���:��^��"E9����    D �{k�=ꬢN��*���e����gv��]j� �HS_�LLh}���`�vo_�n݇(>�   mE�   3Ӓ�֗��.�s��������mHBR�7�m�*�j�'    @p����:�쾛���*���Sn���mn='���n�	Y��IRl�n��(�#�
�EG�7��F��������ҳ\-��:��v�,�'   �   "��nG{��ͻT؉Z�6%.!S.�Sy���go��    a�)�uU��}�N���[^H���ђ���x%�Ul|�J��(w�j��JM뭄�4UW���h�l6�6�l�_:��Zw�K�   �>    ��e����N;��K'�>�B���Ug���K1��:|p���٠n�    n��{oy_]DaR��)��Sl6����tEǦ)1�Pe�*.ت�<�l�(�8Ke�K	��)�	  ��}   @�N��>MI�1ֲ���H{Zs���i�=�
g�:3�ͮ��d��P��mV�/�G��U/     D������~����]Q����[�J�R7󷝘�4kJJ����HUy��v5���e��   �   �����1�>��o���TfR�.�0�Z�����q��z�u�ٞ��Tph���Z��G��     ��R���������������[�' (�X�&d����-�g��  �n��K �j���   ��)�󬩾�yE��;�e�[a�^�I��7�4^��ޢ�rՙ8���wD�*%c�J
�k��U������g�>��(ϵ�߳U}e�]r����fll����	)�BBL�!'��IrR �G	�w0����p��r�-���J��팬�E��J��Ǡ�ݙww�^����y�    hc���»oި.��/7�+m��S�͸�<�dE�!��*�V�8ư� t>�O��媨��YA����V�:߲�2�B!9Q$Qrr���   �`�ٽ���J�WW��^��g�QIEu������S�=�^w�=p�tM��IUT��x����׷E{ש ?A��F��r7�xӌ��2���"    �Ԛ���V�f�.��������=4�����J�s`�T$\�H�Rftq�U�� tYYYھ}���}V�/,n�`�U/;;[�����E"a����s.J   �����jҐ����,���Ŷ�X�IO}�:֒wx��tڱ��[���p��JI"�?_%E�ھ�%$uSf�A���u���w��3�p���)\Y     @�LEf��۝��b(��O���<���%�w�r���b�x<*+�' @��p_M���8-�W���   ���̀~1���vnA�~���#���KҒ��i�iZ�=O]�!b�|	�J,٣��]v���MRJjO%%�ʭ��-ZjڴT��W	    Р�E۲�l�;�{#����7Љ�\.�R���<'�>? @�pJ��*$�}�X����9�>   �Y-x���I>o춟<���G^��UҒ��r鯗M�i��Ve8���0�JL飄�^
��SE�>�oQQ��pU���81�/��q�z    _1d�V�^l��iM`��磫�p8�/Q����S����>d-'�"��s��տ��盘\�9�]VU?S �Υ��}�����>B}�G�   hG�O����ƶ���J��zK��ޒ��=��)�t�{��+2���=�%%R�b�ʂ;j�������	    P��SL|B8DD����"�����s��?�W^5Oa��Cn��rJ��*�q�W!=�a*�S���v�_N� :��
��w��FG���@}i)�>�#�   �������3�j����D�x�������i�{[t+�zw��2+���w�;����    �n����R8D�_n�4p��524\���/��. �Si�p_G��j�w��P_� �   ��������W/�oy�}�5|QZT:�%���ֽ�Nӌ�>�p�k:�py���W�H(�T�W�_�    �0Cƿ�Z�2�~�   �]{��::�W���}����>   ��x�M��+��ܗk5g��FxK����5'��-QWf��MH�u��i�PD�e�T��\    �#�Ҋ�;o�R�U�������>  �b��֮]����6������9�o�p_[����S(Ծ-��2�   �66�W�~:������2���M�𖼳Ι�7Wm֦}�¡\.�<��j�_    �:�zC�S�_n��y�j�!   t���"�[��M���ɑ�㖓j���m2���9r��u���>   �U������.���6��V���M�zt�%����� ��;�Z~�aȉ�����    Nb�{B�L�]"�   ���   ���T��Ӭc�"�6��V{.VK��>����������*���-8�6��#��A�ʪH�{�m���JJR���pDr�Fת    ]��*o���P?CV��:  �!�8@��$%�<���w�4�����{��(-���P��KU^Zs.X�"�Ғ�q�x{��!��   `�����E    �.�����{c�P�J�=�k�F8  h]�O���zilV�읩@����� Ҽ�zd�2��zK����Q�t�Q�5.��R|��*�-�ݣ'��W��s!�3k-#�s!�s��q���_�7�W7��}�쳯�L�ݦ�?^�O6���        �b�\%4�����J�9����  �J�|�\Fݝp�j{g5�^�_�V�=�U��{���x\N�cy�.7���|�1���^�����ௗM���:s�[R����z/39ў/����>^�����"-)	���        t1��5B�2�F�}�   Zٚ��Z�#�n��;�XmC��S4yH�e�}� �{��ߨu�>iɱ���*}�y��n�Ӟ`�x'��ԡ���VE�׮�H3�{N���p
k.,۱W{�K�=jXA��;�i�ν���[V��R5uX?�	�����Ǩ*�/^�'�"�        �嘫�F2�F�E�  ������߸��ƪ�w�4�������yu�]�g��x���|���CG�?qP_=��s�=%ѮX6���t����hW?��\�����9��m{.D�?ٴ�}�+B����������:�����N�Nko_7e���L��ʉ�        t1.�{��8��M���  h�����~���]�.҄��t��!�mg5��`���Ӛ=�����M;������.���*~9=�ف@�#5f.����ѹ�[�]=�����J**�����
�u�+�}��e�9P��DND�        ��1�p��(�a�  ���b����)��zw~�Ʋ���ڵO#{g��c�{�C�x}��X��o E-a�`߈�g�Zc��D�        ��1�"��hf�{E�  ���Ae���hU����`_��' ^D"ͅ`��B������xm�`        @�A�Q\R�) ~Y�Ss��_�Te&'�2���-߹Wo�ޢ`E��c7���}����{������FD�C��${ݪ,���D ��M1 �n��m�A������3��6b`l}َ��7}�W�-o���V�        t1��C	�Ɗ��\|�_������̘��=��ܯ�*�'�����@{����4է{l���W�O���q7�2^W;�^��S��S�V	 P7W��uS���19����"��d]��<�o�^�����g�wp:k.�p�X]4���������ۥ_�u�&�ko/�ݣ���ʩ�        t1�pE��(��F���j���o��Ӈ8������]T�D�W}����{ܺj�h}}�0]��}�a{�����u���k��} 4ϙ#F/W�4�HJPVz���ְ���6�+�e����ʪf?�����I��W��W^#�@{�m.�<4[9=���7a.|}�0��z��D{�i#(;��bU��s젫S�        �b��`_c�J�>�	���Wp����ao[�S�{�
=4o�!m������/gL��@O���5蛏α��6�UEǪzc�� h�2��a����ju~��z���*oA���1&ɲ��*�W�	p�FNO�e.䗖������\hJ���3O�����X���^Y�^�ሜ�`        @c�T�Q��{��q�%��B}V��|�֠^�"d��}m�F={��:~@%x�z�gj�_�Ў�`��eC�@��Q��vv6�� ZSfr�~s�d�MOџ������#�s&��V��j��[P, ^X��~�Yѹ�̅V�?\0U=S����rp�>�}         ]M$�l�qL3��_8܅cst�1Cc��{�����U�҇_ч7]��i����}�s|���}�Yg�d��:g�f���  Mw壯��~����h`����隓�QZ�O?�~�F��Է�9��-C�6��}������>�+7	p�+�#��e�<�>0n��B���ft�4f.�~��rx���jh�t�;z��s�h�5��6EC������r*�}      hS�[�+s�R �c�t����~"9B�. �p��������u�Uy�/����w��}֨�vۺ�{��{ܛ�6�̑u⠾:q`�u�`��b�  McUQ���N�UT�O6��#���^�A��3z��?y��hq�ǵ~7?u�yv@�r���z��%�����:������F������_�-���� >Z��~�\/_{��B�Fo{e�z9�>      �)�L�* �fFZ�Jh*��Z�E_��P�N7&���f��m���M:��U��fw���ʰT~�����9�<�������.��u�D��j�����8b�����ok�u��?�:Nkd��	�{�٫��d�����;u绋ģ#��)�[�Bw��}�����3�Ǜ:�`         ��4��B��n���a��8���}c��hq�&�������'��'�j�16��[�6댑5�w�.?BO.Z% @똿q�]��wZ���S�H�CN�9&������&����>�B�y}��xv�\�HQvt>l�_��zu�U�#�]߯�|n�Bᰜ�`        @c�с�J/�}S�P'��, 7�wl}і]���c�V(��q����7���ȴ�2;h�n�q ���WRf��,i�>��WoV����_��D����%�ūW`��!s!��o~��z�b�� �˰�[�J����`        @�c�#nY��9B=�Ӣ�+N�+5)��qo������֭�5�ɉ�Ql�e;���u�hl��uK��N:F���  -g��J}5����7�g7�|����ߖ��_f�:�#�BI�Z"-���� �U����BND�        �2�*�}9]@�HJ��7���Ï�*�4&�g�������ځ�����>[���  -s֨���{V��=��Z��=]���B�<��ק+tˋ��4t
������wű#�jÖ/sw+���B�        �2d��2S�U`�=�$3G@���Ԩ�4�i�Z��|W��ݰ�@�/\��:q�])��S��wo~" ��.7\o�٢�����7�/�}�i��'��5�7 #M������~?y��N��֭���&c'%%���Y��222��|
9�|/��w�lm�\X]���7�����Wi�����Yg�t�x��T�         ������'���υ#�2�E^ċ����&��5FM��%���~�?���.�0B�^���:N��T��K 8�Փ��=����Vm���۵%�H��J�#���WZ����#�*��ޝ���]T�x�}�X��򪰪���yѩ>�����k�d�`��YK[0MSEEEѥPNP\\ܥ���Ict�Ӛ4�D��,�u���y�~���r�n�iW��Ƴ͊�g�_��h�Yc��v�K�"�   �����a���71�[�VB�!�6��ZU ��S��!e&D��qEUX�U^%    �L�[�/�ja���H�!N\馦bSS�	z\~iӂ}��J���K��S�+���-ӎ�O_|_ �#Y!�3�^�p�.]���U������z�ǭoT���tr��
��Bm���0�kaa�:�ꫬ�T[��3--�^wJ��)sa���\�G�s�H���	#�!�Y�EW=���^�S�   `�~B@cSw�z���׀�W�ӂ��[�و���G�R���?M��@u��[���~�`��Z��~����    ]�a�Wh֬[u��m��i�I�安2�6=Ѐ6�8w�f�d����٬1�e���o�[����Z��IY�x������?�R��9#8  N�м%�YԤ!�ꑒX�>V��/��֣�,��V::x��#�w�갛���V{��jԄ-��®V�yg��1PgQ���u��M����ezi�:9�>    ��+T*R�Y]��T���U��8�z��럘���^��     G3����oJ�1Fĸ�j}�'�n��Ú��R�Ԥ&���>r`l�jK�V���>�B��y��n�~>�D]��� |���k���������;;39Ѯ4V�Ԟ��ܵOE�X���?ԙ�w��FZZu徂����g�o{���p�U1��j䀌4��pK��?,��m�̀zD�V��x��,�:0^i�����Żl   �֋����ջO(�_�[�\�+_�Jʚ�8��d��}b�;
�zk��&�sT��:n@�����b�lx[ٽ�]%'�R�7I!�K�e��Tx���#D_��&�T��/    @�0�Y����o��r�]#
�#�7n��|V8��r�Ǎ���5V��4�>�l��T��뇋u��1v坋����� �HV%���
��:*�W#5��Q{��:�|��gْ_d/�!�\��K�#�   0�_/�}�iM:ƺ(x���zd�2�6.䷳�D�}�	�'�,U��θ�Y��xc%��z�s�O0Y�? ���jK��|u3<
x�ǐ�r���+1!]^B}    _cHZ���E�S���ϣ_\�HEUX�D�3c��=��c��k��6�/�j-�w��;k����`EHw��P����bά�OR^�i� ]OG��jX�>�=��¶�9�|��Ñ�   -0�{�~~扺v�]��;z}����_Z���OO^u��m����˦i��O��m�;Ι�Y��T�6䪭%�j��0eD�W�0�K��|�$�d�SD�q    Nf���f��%�~U������c*r��Ë8��GKtű#5�{�R�>=w�����^ԞZ��򬉚1j��n����-a}�GS�);=U�F��NP1 �v�r���V��K[���v�����`   P�܂b��;����2�-)A9=3�u�����D=���u�c���e�
 Z��.�0���;S?;��1w~��N���N<:�m����܏���?��
�7*�\n��S2�����|C$T����    �khZq�O��ߨ�2�5���5�[@�*�]���������qkd�L}x�������u���`s�������:w���m�}���_����������T�]:�޶  ��i!�V����������}.E���`   P+�w���z_�ףK��[�tOI�o�*��s���h}�
�*�����a�b-yo8e��D����V�{/����>=mU
,��T{h�
_rjo;�WUY�ʊ��lWIp�z�� l��E*CEڱi��H�*!   @�f�~r��w��p9�N(p�=ߋ~NǬ�+���z��s�#%�������L���S�ٖ]�S\"�ǭ�=3tt���zw��x���6֓�V�S&(�g7 P+�VY�>�o4�ߟ`��Z����ߪ狖#�   4Cye��l�>޸]��x�����V5��8Z�����1�Ӓ��Z�6���ʈ.no���4�2d�d�*T���\��mRf�!�ޞ7���    �a�+�D��zX�<3]�^ڥ>!�q���p��Z�3�l�NM��I�v�	��q#�9��>b@���ٝ�Y�}�7Vnj������7��>[  ԥ��L�sh�}   @l�[�{��\�:���[$mL��Ҕ�������ڞ��^RJ��s����g��سn��J�$�x�z�oS���    8�!�Դ~;~Q$ݮ�b�,OUPOF�c3t;����w���|�3F����7=E�ɉ��
+/X�e;��֪͚�a��"5ƿ?[�^�O싎ѐW������DI>o�U;�	   #�   ��ܕ�	��Ѥ�Ӓ������-���ȟԳIǸ�>�t����**ح��^    8�!�W�[�����7��. -������:�܂b=�`����>Zܤ���aY�B   4�>   ����/:d;39��5��zcZ�:�oc��	JM����*.2��ִp     �r)y<��wO.��O֩K���+E~J^    NC�   h�ϡ/��F��j�ג���Z�n�/ү�o��`U�KK梨�m�+���Rnw��.)%C~�W�F��.�K    �b=���f�O�Tz��;�	f�s���b��   �9�   -4�w�!ۛ�����}o�V�wX�=��J*ڷok��
d�UR�U�H�\������a���    ���1��r��xש��o*P'�6���LE^6d�    D�   h�o�p�!���֬qjk����/��ֈ����+�e�Tp�UU�ɟ�ߟ���B�{�0\�۫�D    �X�����5/���3��xc|_��y�)����H    8�>   ��>�]2nxl�2���/m�x���=8Էy_�f�-xkc��{��I�?����^�ʊ"y�RJZ/    �Ð��
�ԟ�5��O7�Q�r������   ���   ꐖ������'��::���q�HM�}�}w��Hk��o��Z-yO�鯞�I��"���yG���l�[����v��b�!E�U��x_    �(z�6Ј���2�ʢ?����ͬY�����ѓq	    �`   P�+�e/�a��}�?��i�739A�	�Cn�Y��-;�Y%$e*�T����    �����F���-&ޢ����O���xvw��O:K    '�   -��ڭ�����r۞��v��eӕ�=��zVz�f�~�~��'ꌒR���h_�*�ھZ�{    ��C�nHK)�����a�,���7=}�}    q�`   �B��di��~��n�8�0������jo:�X��l���ث��0\��S�6P�6���sb�z    ��^;٭����w?�+��O���� ����u�)]"    �C�   �:<��b���m��^��d�Х��	#��q��v���L�xw���ُ7�W��g����ʝ�t�_�˧��^�K�l�N����"uF��=��6T�w�vn[�^Y#�v{    p"�kU�H��Z�����0������PG>���������º��^f
    ��>   ���S;
�����z��ez����\�>�/Κ�/s�حy���r��˦�AA�ܻ����Ŷ�:g�`�;��5혬����	��;�*++k���(-c�����c�e����t    ��0�2��҂��̻�������ۯ-m�����?�ޙ2C�D�P��   �;�}   @3-ۑ��{]/_{����Vž�/��	���JC�j�N�	�{Ŷ����v��r�����Y�HJ��o�~��,ߠ5���Yy����׷E{ש ?A��F��r7�xӌ��2���"    �G�Ҹ_�������9{Nt����}���K�m���(.</zQ�툩����A�   @�@�   h������W��cG��})vH�o}��1����qBl{}^�~��{�Ku����+g��~��n�{�}��U;+�˫��!���UR���[�PBR7e��E"a���f�L3\�D���"rR��@    ��u��%�+�K�����ͳ�c��>���}���l�n�o�i�O�H�*Xx�#��A   �3!�   ��/���YGV �oo[����_��`Y��Z-x�v���Ӵ[�WV��s_��c��Z�ۿ��?i��h�:7C��L�ҕX�G%Ż쀟Ǜ��ԞJJN�[�����y砢~F�J    ��cFv��UѯWUE"J�9{s��m�Ls�)cu�����"��(0�U�n���e&+�gf2D�ˉ���=*b�� 9>    ��>   ��� ���-�[�Z�|^]?u�f��q���<�X����~(:�'�j/^����	��GJ�����Oқ�6k���_��0�JL飄�^
��SE�>�oQQ��pU��{W�I~y<�k�    ��4P�bgV��L��mʈ��U����{�o    �*�   ����wݔ�J����k&��>��ު}��v��i�Ŷ���7o,�s��ѱn{��XK�D�G�\r��{�+��%�K����)T�_e�ڃ�.�G.�O        ��"����0{iM]�|�2�   �V���\�~�ܮ�gi�j�Ղ��K��箮0g�n|�]�TT��8VK����joO���N<Z�,X���
���������        ��������^��4M%%%��x>�O���=�H$����9�   �������'�o������Ym{n�k��[��Q�s��i��XK��ϙ��VmVnA����Qbr���f(�T�W�_�        8�U.++K۷ow\��
��ŭ�s��Z�KJJ�9�>   ���..տ���}������C7�vll{WQ�~=���~�9�%oj�O�]6M_��.Ӓ��՚7!���[܆"*/ۥ���        �䴰�iF�l|�|sss
��ա��;_4�>   �������	G�Z�^���q���ϐ��s��並�i����=eX?]>a��\�J�\.�<�B~        gsJ���C}5����#��l�   �V���X�~�FW7��>�j���8A��d��j�*��bc����w�T��n�v�����K�;������        @�::��^���#��|�   ��_��^Z�GO�m/��c�|{iVK�a��j-�B>y#�ߧү���Cn�{<r����G�K8�mV�*9mH�������֑        ���}���Q�p8������   ������"        �c���3��Q����#�?�            p��
�ut��F{�/���B�            ��Xa��kת���M���}���>V����׫���M���|
��s�h�>             �STT�u�ֵ��999�x�r
�0TPP`������9r��s�h�>              �`            �A<nuOIR�ϣ��v��4t9̅C�            ��eFh\vO��.#{g*��?��²
�ې�G,�;k���~0y�.?vdl�����L�<FD�Bz��?�}�d�5��oy�}-ںKNE�            h'\>].è�~+�w��!���⵺����*������M�>w�]���{8���M���zsaD��.�������            ���=��t{���UT�D�GY�)�<$[�2�>�͑{���h��Vp�KN?$�8պ��Z�ۺsa��=��-.���            ���������� Sm�Pލ�NЬ�O��/����-�'�w6�1N:F'�k���r�.?\��\�D�s�S����L�����R}�iG�cO��Y��M�t�$�            �v�����1M���"M��K�b�v�Q����-U�:{����Z�i�>8Rc����}��u���s�lk.4"���            ���b����)�>NS�ߧ�ť�ū�c ����c�����υxg����|�8V��O~wD]QU��+�+          @�����W\ڨc.?v���`�����*(��"���B�qs�3��}%%%�p��е��
v�`_8�*�}          йL?г,۱���{�&�w�l��Y�A//]/�3�6b`l}َ�F�2�'�U^Vi�R�V�            �CXa�릌Ӆcr���Eziɺ���S����²
�����5~8e�.��\xqq�s�����k�����vIE�>ݲS�,]�����~NG�            � g��>�{�
�e��jʰl��;mK~�.��+*���w�sF�c��뿜3O��Jē����C��ӳis���a��N�{uZN{�y�q�޿��g[v���            ���wx ɲ��Lw�]�g�X�`�)���_.<�^�p}��l��x���\8����_Z������3Mi��<m�+��Ve�>i�vH���`�n�z�����-��T�             �LN�oΛ���)��۟�2�s��F�띖l��~�ܻv�	�,��}�9w���Ssᡏ�荕��������.C�8v���)v���[�r����c�ph[^�}            @�����q�z�ף���%��'���~6�x�o�s�"�$��j�<�({��o~��{ģ+�#��e�>R�s�Vk.��oF�L������/�s�pĴ�Yn�/�K����럑�KǏpl�K�}            @V���(��[�~�i�Y�L���B���C���c��G�96����O�aH�s����W%�_m�1�>j���΅>j���G�s���u��#����            аm���������.��<u�����kW5�Z�^��۪��ݢ�WG̅S���y�[�r��eb��Q}�˩�            3�v�jY�de��*;�����=���2���Eu��s�b뗌�s�b�o�_���|R��<�R�`����y��� �"�            8о�2;�dIK�IG��vJO�7j<��m/�²�8�!s!���m~�/�獭��*�T�             ��{V����e�ܿp�.��F����e�o�/җ�v��y��8�s��e?�'�[�V���`[#�         �aL��3��-��Z���w1͖�rE��P)
 �s֨��J|V��=��C���/u#ƹ�QYu��������ē�����f�������cb���&�"�         �q�p�	-��)��5s�Z�_�>V�I-�,l��
 ��K��VoVAYE��M��Kw_|Zl����Z%Wo�u��Ç��؉�	
�Br����6<����V�).���Woi�\xr��Z�cs�Κ-*�g��)�z�g�O ��.�
�_���S�         �0����V�y�;��Z<�����i-���YA
 h/WO:F�/9Mo�ڬ�vحq��
G"�HQ��dM��3F�˨n��fw��zw���`0h���-�������R('(..�R�{��1���[m.|w�h������}h�g�w��X��d���#�v���߼>߮ �T�            �v����1��!��ҕ��QYe��+������P ��+,�ذ�ꫬ�l�ǰ�7-�:��p_S�¢�ѹ��9*��}J�{u����R��HD��֧��_���            ��yK��0�IC��#%���>ߺ[�~�\O,Z�p�k��m�P�����׎
�Y��֡�5aFKG������s�m�s���υ9�7*#)Q9����rպOye��߽��%�����`���Z]��

���ϋ�� ]�ɪ���KG�r��޴��-�\�;M["auE�#-oC           h{�/^k/V���NMRfJ���
V����T�v�SaYE�=����x�ޡ�V��
����v��:!��BtX�e`f��-����[iꞒh/)~�=����V�ګ�pD���]���_f	h�3�`*�`�w�(�kt��О=�:�D��S�&��           ��)m�Wh/��Q!���i�����	�u��R��Қs!k]�~{�w��  q)��Ɠ�!t.��V)y         t|ȭFZZuq���9�|�p�U���h�}   >E_`Fܼ�         �SBn5�p��*����:�|�6��_᮳��p             ���Q!�V[��f���B}5RSS��g!�            �]Y���J9���o��su��&$$�s�}             �]W
�����D�              p�}              8�>              �`              B�              !�        �
Ҋ�h��E2d
�����Q����    t�         Z(P�G��},Chon�tԲ��b�4Uy    ��>        ��C}k	�u$W�RG-�p   �N�`        @3�s�}   }q1��*"n�"U��*LW��o���        4�>�!�׹�����_ZO��Hy���S\a L�ߢ ��D��̰�
#�r��A�        ���9��#bF��|��Sh=���3���8-  �3#�        �����p_�`����h�f0[[��j��..�}   �!�        �H���ᾎuͰLe��+��J�<Ʈ��C���nuK�6y��^�q�D���U�7i�*CUG�����7��=n��������n{g�   :#�}         �@�/���8~�2=a{�G�W�IB��=�g/���v����V�  �Y�        h ���e��F-[+	�   �#�         �A�/��	�   �3�         �@��� �    ��        �Ejq��N�&ܷ|��x|   �b����\t���         j�=o��N�
���� �[   �8>�Oeee
�Br"ӌ())���s��F"a�|	�9�>             �.;;[۷oWEE���
�����j��b�onn���}�pX����h�}@2M           tYYYY�
�Մ�ڊ��}��Z�>8�>��h�            �8���j*׵5���"�H���2���+�           @W����
����6�ա���\���bz�$A       ��!gh_�|�Py�-��~�>���r9Yΐt�|� y}���n�.��Q�   йuT��
�uD;ڎ<_B}�G�� �a���       �"�}*--V�>�� ܷ~S��*��t)���U�wz��>_��Y�!7z��A  ��h�[G�ܺ��������ria$U���       �ZUj�΂f���o.�޼]с�#�a���=���6lܦ��J  �����nN	�u��E���Q�7As�	�jy�       @|��}�
շw�Imy�Pߞ]�75ι}2��y}����K�  ����nk׮Uiiۼ&LH�{��t��E���S{co��\/bJ��d�(si_�@       @2̐vX��z���n�oǛ��g����۱so�|3��4��Ԧ�;��   iݺum2vNNN���[NRXX���׷��N<_ԏ`:���a9�       ��*�mڲOUU%�[RQ�3�6mޥ�F�JI��:B    �U�            :���V��$%z�
VTjWQ��hÐzF�M���3:fi�R����\�W�            �vrل��Sc�ˈ^ꖔp���e��!W�,X�w�li��V��k�����85����Qw�νzw�V=��+B:�5�F���V��}�	�1jP��CyUX3�{VND�            h'\>].+�W�@�_�b/�}�V?z�?��
78n�@���M�]����qO�e/��ؤ;�
�H�_6]nW�̅~�R�`S��ɩ�            �l��Z�=Oy�R�).���e��j�,���\<.Ǯ����Q�XV�o�/�����vU$�y�kі]*�)39����wZ� 'Y�W=�yP�\�2�߭c.l�_�Ź{�x�<IK���/-]'�"�            ���S�7n׮��Z�*��x�����������[�O6�s�����X�o��]�������Y�OԷ����5O�?���O��Y�ѹ���K�ɦG����>�����n���wcۏ/\)�"�            ������p�ԝ�.҄�������\g����c5�_u�e;�t��^R�"T�Ӵ�T�44��׻̅s̅���PK����=خ`i��Q��qU�:�>            �a^_�)�뛞R�>V��Og�����gީ3�ī�Wl�����-��G�����s��Y�            S�����j������@���;�8׹�ǀ檊<J�=Nvz�N��o���a=��9�>        �R����lp?ӌ�P��U������o�[   ]���c�K��պ��C�c�sWl<�>�ۥ�OE�v{_ ^M10��tG�����F�eT_Y��bS��Y� �        �
���U��obB�z�H�ˈ(^kŚ���7��V���%�  �+x��)cu�{{k~�^Z���}���[_�e�����x��s�Qʉ���Z�Z-z�����g�>�#+{�����ٮ-,K3u���t�.q��q��\'�'�&!�7	��8v�q��`���bvav�e�����F]i��y��[�U�9#�������>B+>��y~��>}w�6��E�0�/\�V��qx.�u�艭{5Ƽ�������&ko�k �        H0#�۾sbQ�!8Ы�V�l�gD}�w����a5��� �9G����{U���uK+TY�c����[��S
���񢼬��p$�W�r�V��s�G�VZ`�>�4}������-{a-Gυl�'62bs�\ˋrͷ�7�sɲ
���i�7u��=��:�>        ��l�wlܧ�1٨/n$�+ȓ-��  0_\������o�٠G��}Ґ)��9�ΝWiYA����rk�ޮmV$՚��~�r�\N�f��W�ެK��sU�X�bs��1��}�n�#o�r�g����W�{x�.G��S�}         	2ը/.��+L5�3���v�g	  `>�K��]���4��K��X�x�/?�{�#ύ���@7����z����������oVEN��ڿ�v�n���Θs�E�j~���[�΅�����a���ؚ��MS�o�D"�        H��Cut��nϙ�}CRu��WW�9ԭ��������FU]�)  ����F�#�1{]N-��2�$��k��u�Ϯ��N+������ь�C��܎�����֟��u�3?}N����fh�xzY![��2����r����hs��W���%y�΅��q�ry���ɛ5���ڡT@�        � ���/���!   �D��[q�A5u�i��=�a����-���W/�=��w_�v�����?,��=�eϘ뭚F�q�^.)3�_�ba,��Zq��p����������?p���O�ڡTA�            XH]G�����o5��ѥg��u������J}�mS�~����oEq� �;~.|96���VMtѾ��:�$�<7��'��U� �            ,�X]�X��83Me�*��:�]����\������=}#�9>��Tp�\(�J7�B�WC�������w��2���            ��1�!��:�}}wS@׬\h�{]�q��s�F΃C�R�1s�����a����mk��<�I
m�k �            ,�a��+��z�'\���}岳��9���Ԓ����W��ꄹ��D�x�2ez�����Nm�nP*!�            ,�U�����F�����5֫��_E~-/���\�in�~��>�z�����;$ ?��R�d>~Ϊ�󟽵SѨR
a            � ���ԋ�k�<�ugV�[�]>���M�F������M���.��&�������c�3^�f�xU���sT��rrr�bŊY���������$77wތw�s��ͻ'�-������sc�<��n��>        �Q����c�p��  @2|�����ۯ���Ɓ�vt�{ �H4���4ǎuK�uͪE�5^����/o�nخ;�Z����tY��썺���r�ټ�%���+�Շ�,5�7��?}��?����1�>�-��]������Ϋ�~v����>w����^��UcW�Ra        �(�*���ߩ�ހ0w�W�7m�~X
  0�ۥ�N_f��\ۤ�~�C�c^czw>��~��۴� [�,�0#�2��>r�p$��?����yPVfD}CCC��q23�d����٩d2��P(4����*q�d��۵���~����_���G�^9���o�P*"�        C��uZ��5�������Re�
   Y��65u����e�O��y�1������M;�mD���ӯu�?����<}�U斻�*g�Ό{���V��F�S�,+KT����i�b�Օ��/QQ_�Ub�^ߦ��\0��-8�\0�^�q�s�p���@_P��v�:�>        ��ػ��g�����  X�c[������f�(ï�t�����@oWS@]��I��X��ϟZ����涼%Y�r;�j��s�uNញ��/.33�|Ltܗ��1�!�q��[��Øbs�x炱"e�׾�TG�        0��E�  ��X!�`��<fZ(֛ՍJ5��uɈ���%+�K�J�qƟ�:6����J�         &��/��  ��DoG;�D�}Ɏ�⒵R!&��        `���R��o��V	H�H$���A�����^]��njVOc�zm�j8������b�x����x��z����QP���2e�>rO9E.�O  �%V������v���M�ʄ�#�.�>        �I �>�>$K4U0TOw�Z��Ss�v�Vہ2�6#�k6��v�ܱ���%��)�ࠢ�슪?vq�����c��.����5�˖���T;JV����  ��jQ_��M�l��x�q���        `�������000���.5TU�i��oޤ���p��i�)�i����&3���z��+�<?��k�F���H�#�C�ӎ�U�߽[�G�/-MK����_~�JO[��M  �
c�:+�\w<��3����x�^��K
��>        �) �3�+Y��ҕf���nGG����԰y����Nݍ�
G��8��s�͕��6��9��|�o��q��h���+�y��`hHU��������B�v�u:���خ ��[D%��$�        Lq�u�!Q�A_kS���nվ�Wo칱2_��%��a�����|�an�{d%>��x��E�u�o�ޮ?��6?��V_w���r�<��  @j"�        ���q�������`�s���jkmU�;��7O����\����6;w��i�~�7��F��t�̯��H����؟ahxX۞xB۟}F�������ew8  ��B�        0M{W�#�K�>$B�����YHUO>��}�d��T�����������.9�U�B�����6��G���Zw��U~��  @� �        �Fܗ�^/�"B����I�0�mw�������W����56���r:��G�ɵ���s�m9�.�4���+���J]������   �G�        0C:s�@z�`�������-��5�333����T
�t��!�ڴ��G�TU%�áB�׌�\
��g~�؟q85Ͻv�����w����'�]�@��a|�].�|w[���y�y�  �\E�        0
Z��n��
�q8�wť
z3��9�+h��^�W������z���J����o�˩��\�ϺI߱�큍(n0������F����u�ޫ�K/S*��>�`8��;  0��        LS~���n���/�j���e	��@ ����n٢��B�HD��Ҝ�^�o,Ɵ�X�ψ����b�y���V{m����'   k"�        �#� �K*[4��]��aZ�Ѩ�����ޮ�ohׯ-cm�R�G>�Cv�6#����1+;���WOjh ��>�9��>:  ����        `�������aD}��5��������v��������x�|��ph 6��ؠ�?�[���ʯ�1q  ���        LQ��q߲]�h��ˈ�0)MMM���V��^3�>�ݦB����v�1"E#V�H�g�7h����u_��   `�}         �D�g]�h�����Ң��N�nݪ�瞓�X����>�W�3�E#�Ǝ�^�?'[g��Q  ��         &!�e�*�������ѡ@ �Ϊ*�x��4?��8c�F�g���_�Bi�yZy��  @��        LQ_���V\�~����A577+�ե����ш�=>��I�g��g�=��Л�@K�(�   ��         &��/�q_���T���>#����A�pX;����U�v��_Q_��aW0UzTz��ԭ�z��~�   �<�}         � �K]�h��'0��P(���W��Z�N�2\.�4?��:���ޮ���;��M   H�>        �� �K}�}8Zww�zzz��Р�����nS�ۥ��V�����v��#j޸A�o����+   $a        �����>�-x����=V��q�#a��|r���Z}�r�>n�Mv�Co<��*[�F.�W   H<�>        �Q�jTN�7��㾝��R��柶�6�i�&u��+���>���;�;������Җ�׹w�%  f��[��f3��4�Ƌ�!�        EfW�����c�}�`7a�<
���ޮ���<�����r1Ϗc|>��q�X��_i�UW)��P  �4�ۭ���˃����H$�����_*���O#��>          s��Z_4U�
��v����ːlJ�E�嗿Ժ{�  ����L�����݌ȭ��oF�>���k�}��>          s��А����=֮_/�ͮ�C��n�@$��W_V��+-/O  ���n��m��=t萹����x1u�}          �@ px��M�4�ק|�KvV�;)��ci��۶�~���� `�X%v�����ȭ����%�6�>          sV$QWW���n���۔��Ǥ��4�������]rz< `�$;vKT�7�Ƌ��;V        ��\Z���[$�k���=�K�m��-_V�>�H�y2^XWOO��u��h��K�N���7!�W5��������� �lJV얬�m���C�        � i>��}��*Ζ�=��h��.���eu~�K��fOs�{c��CGL��Z_L��-
�3�ӏM���&GԦ=/�H� H�D�nɎ���x1q�}         	bӐ��:U<��͈��M�y�
�;�}���?15CCC���S$R�֭��mr����9m6�w�Tg���� `�%*v3V��B䖨����>        ��j�6�����׈��Rp�����^󱫶ƌ��\.�	���c��t�M��7kŕW
 �D0b���*����j��G�Р����L{��7����         ̌ݚ;UX�-�s���jj;hK��m�㭮�P{�Y�t�0�u��"Ѩ�نwJ�U�"��\��6�> @Buww���l�����B��b�vuui߾}�r���#�        H[tH5u��V__D�nr��	�6���={��就^�T��p$��w�U45�   �.�>          s�����ᰆ����ب4��mx���\v�RNy�  3��t(?�/�ˡ��!5u���'��T���4�K��߅ͱ����������|��9����gH���         ��c�}�����X�&�4�f���k��e�^�> ��;�\��E:��P+�r����zWpP��҃ol��U���N[�O��Z�-,U��5��p$�]M=�e��'v�T��0w��\�z�B�{��`q��Gm?\�ޭǷV�ۯ���ؽ���         ��
������G���o:�6��v54
 0=���ձ����l�ϣV/1�ǶT�yA�'Yq��v����յ���������|��܅k��<�w�[$��y���9����˩���Jݶ�r���f�/?[;{�>��g�������         �s��lm�-��N�7F��};j� �{[;������<�mC˳3tђ2-��2�1%���O��>�����D}��2W7���6W@;��@����܎�,v�'�I������7(�
��vj[}�Zc��$s�h ?=�\0���y�n>}��<�m�~�c���y���wq�>w��J��U���G>�a]�iwS@VE�         `Ή�����"��.�0���X����  �s�C��������7���
f_��,���/0��zF�x}ۨ���}J��o�ן|Mߋ]{��ߪ'�����|�r������ɘ�?0�\0~��+����{d.�����w��`�	�޴f�H�7��?~F��8p�5���-��ǯ���.6W����t�>&�"�         0�����6�ld}3��,vv 0=Ɩ�'�D��/o�Y�郫G{ם�x԰��F�7�4���Uɾ��z}��k��W�ޏ����֓�c����̅��#�-���K֎�w���>����==�Mz�J��u��R]Vy�^����         �S"�����k1C��|l�;#l6��CC��>�6>� 0��yp$�+�N�������-��Oz���Ս�g�H��88�������̊���n�>�zC������לg>7��%�         ��G}�cxpP6�L��>��`P��4 f�p82r��������ng�ڣ_7�& UG���'��0/k�뻽@]'���+�]�j��w=���        $�@(���~�d�2M�9ށ�3b,6N�t����'����rv�C�>c^?4"����j��w�[G���b7nui�I�gl;�Ɓ��G��m8q.dx�#����q�g�qyi>�fe���GVC�        �]���]�&t���WI��
E�~��ϛ�����x#�"�b_�H�gg��al�k�ICA f�Qa����J�ym{��ܶw�k��q@�o���I�[X���D�޾���
3����_`��#���o�:c%�/\�V��qx.�u�艭'΅�����t�[���y�y��(��         �#��;'���آ���&;��@��[E܇)�ي�v$��Xr&���o ��# �̸f�B�d���9~�ʲӵni�*s̷մw�#�J���Q��x�]?|Z���T����|�z~W�^�ScFP�=�h�c�4W&���V�5�	����B�����P�屯_�����G�������}�\h���c�YQt��L����         �&���)eLu�G�}4Y���
}v�K�Y�hT.�W ����ukuɲ����g7葷w���m�k����33���������hÑ�~��{���ێپ��/��¥S�-=���ڡe��؏��R���y�k]�>�S�y[�V�K�>        ��j�����
�;^#�kl���0_�d�l�k���v�ugN$*���\� �cu����"s�yi��}��,��ҥ�N�)�������xy��nj�ޖv�#��
4��\0V����s.����/v��kW��W�j��P�1��0�w�x$ ���� �}         	p��M��ɖ=�����]�����
�w��x�v����/���):l��B�7]v��������� 0S���o�<�������L]�j���^�׭?��:�4_��3檩��������.3��А���v����܊4#v�����y��0/K�p�:]Vy��}�P8,�*�-�]G��m.|��s��$o̹��7��sV�[O�y\z�o�w�o5���iIA�� 6��Cgp������+�;.        ����5��b����t:5<<,_N���n�A(L�=�9udd 0sz��b8���z��`�ܰ]O}�f3����%���5����Nx����[�].��fnYz�wמ��c�1"������N׮Zdn���?_���XE���q��s��o��_�{��s���`�xF���<�G?�a--Ȗ���W/?�<��ﯾ�U%y�b����gE�}          ���c�}��"u�es8ee�i��lJ+- `�նw닏��g�x����.=s԰�/�;ߌ��������а�}�ym��O)��1��xm���`eu=�̅/����^ߪ��<�֩������K�4W�,���z}g��酷�m{���w����E!��         ���v����'a����#{f���05���s(R�) H�7ԛ�]qf�ʲ3T;u���nl7����#ϟ�q��3V%{iO�n9�Rn�C떖��w�����BiV�9��o4=!��o7��ߨe9��n�Ü;����m|���*�r��Ñ��j��         �s������WxxXQ�K �*�ק��N���	 �8���F�d����n�|���4��j}��e�=㯾w��d�������������s����<�w�29�v�����c�Ķ�>          s���5}�����.�0U�K�pDy
 �F�g���=6P�9�٤�[�'��Ҽ#�=����0��������󟽵KVE�         `�1�>��.ON�<�����'L��aW�nS��e $�u�+��1ύmD[z��y��@�#�8ֻhI�I��5�߽���{�;����B}l.Lduʱ\��B7�^b�s��o�         @�Q���S__��Pw�ex�&�X�/<4���r8�3 L�mk+���uOzݙE��m��<h�.skѣEboxaW�>r�
��7�=O��ShH�����$+�<o��צ�FY]nn��/_>+�NK�k�B�Dc�<��xo=�R/�Q�d����'̅8c�ަ�uK���O\o�pi�Ư׏��e2�]        �(��es�ͦAO�0?��~3��Y�XM[ޑ��D �,of��:;Tv�U L��.<]߾�
�vW��8P���3,2"���43L2�kV-��H}���]�z��Q�w�˛u�����N-���_�C����z��ּ��a���"}q�����W]���6h(�����*;;�<fKOO�:;;e��,99�1[������%+��E����Bϛs�A���΅���k~,�����7���{�z��u9�(?K׮Z��W,��~�y��l����}         �h*])�PP9�ղ����Ws�Z3���������Ve-^�h8�a�K�<�ߧ��FU�]+ ����.�|�2����&�����\�ows���ȋ���\i�}+����O\o�60���8�}��-��;deF�
��Jj���o]]ɍ�5���,�m�3s�No��\x��Y���ǜqk�
�c,�?�lܮ?y��1W��
�>        �1�,8�|$��������؊����˖���S~�B����8c���PH��B�-\( ��<��m�V�..S~�o��ީk�7���mکp���ѣ���{�m���胫��s$�;>��x��\��X-����eff��Ɋ�=^�Č��Mͱ�pAl.�3~�q�~�iǸs����+��UQ���׆#���^��ŷ���c* �        8	3�J9m�}���o�2~Xo��W|�Y���c*����&̗����v-��f ��-U�a|[�07�������{�32C��Mu'uߝ�}��ϙ1ߪ�|U�d(��Q_hH���ޭoUG����Ot����o���h�o�2����=��<�m|�f�4;C������+v�T�G#�        G��#+���$���-++��r��P46�vٝNE�����9ry�����%_, ��1VL;�2��dl�k�pf�&Y�[����'j�Z+�א��fc.�b�ԨTF�        0�}���.�Kiii2~�[r��jݽKr��ߒz�C���檿�G9kNWZ^�  �-===J��ܦ�0�q_���8��}a        ����>���端�Oe]�����Pq���"�0:��._V�����e_��  �-V���f;�J���
1q�}         �@ܗ��p4��o��k�T]����mfվ��s���١��J-_!  f�բ��x�7���x1=�}         �D�gmD}��j_mm�*.�T��ܯPQ��^���c9���r�g�.]rϽ `6��Y1r�s�=3z��6^La        �����i�!��>�%--�<�眣ƽ����H=�5±2KJ��P�U*9�T 0[�Ѩ��6^La        ��,<�|$��>����X�«�Ѧ��Sw$*_v�:;�ü��rx����֍��   9�         ������0n�[���
Zr�u���ߨr�29�Aj��;��,-U}M�N��6e	   �A�        0M�}�Eԇ����WOO�
�X��͛��PyY�����D4o��ݕSQ���}>�~�M  @��        � #�k,]%E�q��K�������*//Wuu�V~�N�����t������ؠ�*��P��|:p࠮������   ���         ����xTPP��HD+���v���/�TZ^��m�o|YY�ث��t�g>��E�  ��"�        ���QN[5[�&A͢�Ԟ{������U0��.Uم�Ж-Z�p�|�C
vui��dd(��\��)�̳��+  ��#�        �&���Zp�m��URR���a-��J���u��N���*�h��Gs���WvE�Z[[���%_��   `�}         �@�gf���=�������Puu���x�v��'�ki�)ee�76���<��f���ѩ���������   ���        `����eA�;�#q&#����h�G?�w����j~v�S}���_v��J���ݭ�`P����'-M   ��>        �) �&�>L����U[[�5���v=���[URX���k=��R4�� ��P��jkoW��n������   ���        `������S�t:͸���N��[{Lu*-)U�߯�C��������+�NOWCK�B���Ͽ!wll   ��>        �I0�1�>�#��Tķ�mhh��;>���U�Ν*,-U���ml�@w�R�'=]Yee�é}�5�\V����9\.  ���         &Ȍ�Z��Rq��������.��T`�"��i���L��u76(<4$��;��(*�/;G���:x`�N��6�vÇ   k#�        � ���Dܗ�2_��y^Z����l�܈�REnn��~�\.�ҊK���G4��{{�r�-UK��mR4*ˉ�{*-��O/,T�fW}[@]A]���P�eJ5�pX�`�<_���sw_j����KϾ-  ����        `D}���/����G>Wl�8���cI�׫E��5=]�{>��M�T����+,Tn^�
cGG��E�a%]��Q��,���r�s0�C�Zx��ꮻ������GJ�ît��-�3<l%  ���         A����>L���`QQ���������b�>��j��]X�̜\��?P��3)[�[�������]����ɗ����ꯕSQ!   ��>        �1��-�}��ǣ(''G��jۻWu�����VeŞg��)��HC��f�7��3����y32��ʖ;-MQ��;RC]�\YY:�>���+   �&�>        �Q7�"ꛃ�nQ0=WAo������4���._����{����)=7Wi~��KJ�YZ�ၠB}}���~E#�)\��nn�kD|�����ͭw"a5����-���b���{Uq�  D��w�l3�;`��[`���C�        0
�@?ؚ��Qy��0m�QRR��իh�W��ղ�B!����u��-r3���]�ᐆcG��p�F�#�/ˈ��)��v�v��9b��4�[v�;�Q��]6�=Tgg����)?����{��h�  H���q�EbO������Ra�~�d!�}          0E������
~K����պo��v������������������n����m��ُ��X�'j�D�
��B���HD����ѫ��~���py�N=�,����\� �TTVV���z��n�pX��}3��:^#����3�>Xa          L���Mzz�yk�y穿�_�]]�ؿ_���iiQo{�B��2�>#ȳ��
}�j}F�g��g�p�ض7�*-/W���/����t�jy3Xq 0wX-v�G}��j�G}��>          �aN�S����QZQ{˥�F�V$�P_�B��B�}
���t���ʝ�.��k|�� ����v�g��СC
�BJ&�{�>�"�         �0V�s�\湱�/  x_��DE}q���I��G}��u�        $�������r�Ӿמ}mz��2c��b�u��x��+   �mɊ���%+�#�K�}         	�����ݭ��yܶ)�g��.X�,c�]30�}����#  �|��mj���%:�#�K�}         	bװ�:��Q_��)v�[xNw�F�זB�  ��HT��/n��C�        �@F���ԩ�ly\����D}�e��}?�  �|d�nUUU���{�^�*f{��G�Pb�8���        $�MCjj�TAa��N�����u�d�7��V�v���Y   �ߺ���w��Y�weee�{S�����K��훕{[q�89�>        �$0b�ں�����
��/�T7��    �a            0��y\*�HS�`H-=���+��E�            X�-gT�˗�9�|SM���W'��^�S_�d��<k��d���g �߼�_�z�m�nn�
n>}��r�Y#�7�6�k�|u��s9�ZQ����򵦬P�K��q��m�o�W~�Ra            �d�>��-�*��y[{����wa^��􇴼(���2�n�y�J�tF�����zx�.V�yi���uL`.��S�U+��p��z���R	a            �d�t�%�D}������|X��9���ޠܰ]U����{t���`q��N����+��ݧW�jX�?����Q�D--�3�KE�}            @]�bs^�/����k�O�}���G����.}�;����w��￱]������uN�]��z����O
�X�u��p�炡��[�ַƎmoh3W���^�TD�            $I�׭��2��XI�M�&3e�<���G��/�����]��BgV���~윕����X�9n��<uo�~���I�}�~��
�)��i�}            @�����T����А��c/kq~������s��kh�����H4��ߪ���5�scE4�>X�1J���8﫱�� 7sR�|ԗ��            �$X��\�8w�y���m4��\طp��ٝOz�owU����f��˔��+8(�
.Z��\0V�4���l�7��        $�`(���.�jN0����/  ��+����W�f�6�6�{�o��=V獜����_UK�V��a�ie�}7l�l�\��헛s����)ͅ���         	�{��vM�Z�7]E���&�Y�d�����8?��  0����|-��R(֗���v�A--xu��@׸�c�h�}��Ź�}��o\{��R�p$bnG=ٹ0W�        $XW��}��"7Cp�W�-�f�nK�rMv��^5�*�cF  ���uJ���������������v��v�<o0��G�Q�e�	H�3+��ך����fmoh#�        H��Fnq���jlё�O)c��5b�x�gK��  ���p�?��������6M�>i�c������z��t�K@29�v}��͹��u�sa�"�        H��ި���=����}Ņ�J�o|�¢/  �D��gkeq�"Ѩ��ȋO�>��V�3�.5�1��a����L_���)+0��=�Ҕ��\E�        � յ�
�{$[���3��v��fr�S`�   QY���^~�y�߿Wo�4N�^��"(c�3��fR'��G���_��-�\�_G������`�p,�>        ����5��b��  `<F|��;����P]G��{��iݯ?4t�s�G��7���T�wpH@2��R����Nc.lND�            ̲O~`��>��<���/�o�a����:���W��Wm{�Iߧ �7r��?  >yީ:oa�y���^�}-���            �lI~��h��?w];�uGo�{�rU��y�|(Ѳ�z`�5#�tki����gg���Ů��ji�Gυ&8.:j.���ң��\E�            $��&e�<��小\k�}�3�xط��@o��^��~���<���LS�F�:�            �l{c��ܶw��
3��`q�y���?녍�͎���:]�b���������c�����]������z$�{���sa            0�~�y�y���S��=�c������<;���8��q��6��\�Přij���ڏ��j�|"Q0[&:.]V�'?�y�c��0�            )���GOl۫[Ϩ4�*��M��?yF�/hv��R�y�J�+8�~��RANN��/_>+�NK�k``@V2����}Ra        �(�3��Q/�-Q�M��  ���]�|��|}x�R�������QU-���u�����_����[+hMOO���l���VWW�����W����1[���bc��\���@�>��c޶� {�|I��[�]~���
������"�>        �Q�����v�07Q��ʋ�	  `�8��'~�����w�t㚥�1��i�s��R_*��gD}CCC��q233�Q��ɍ���/
�����ʊ��f��q�-��ԧ�[=���V�ǿ��)@�        �jZ���}�/����	  `�ymo�.�ׇ��7�3W�3V�;:���֩o��y{��.QQ_\FF�����/QQ_�3ƾ;6W�        �q_���Z�N�i���  �Ly��V�_����ψ�>���T���i�*�LSWpP5�]��P*Ht�g�}Ѩ��]�ƛ�yx�d�T8�W��Mj.�z��)��"�        q_�2����ߟ-  ����7���j�j�����^�.qq_����dŌ�8�>        �	 �K=D}   �!��юň�l��ߖ7�Q_\�cFLa        ����>  ��`��/�X��0[q_�W&<q�u�        L��E�QUԽ+XQ  @j�Z���f�U�_��B�        0Im�K�G�>�!�  HF�f����v{f�~�m��>�>        �) �ͦ�D}   )�X	{>�o����        Lq�u�Q������    �:�>        �i �K>�>    sa        �4q�-QY�Nc-!q���*�)H�   `!�        ��E����p:���P(��v�]6�M�����9����y   FG�         �r����Pn��x���E���������#g,�����<3���H$���&  `t�}          f�{��Y�no�l��I���O^�L�{��������N%�5�+t�ى���w�58��U���,�eM���}Ca}��w&�~v�M�?{wW��}�N�h���]��+u�EZl�XX��wم?�-���,�Z�-5���K�j���)�62!�ə���:Wf&Ϝ3g�<gR�7���u=����j�   �D�         @����1p��ڭ�P����vᚸB�����v��K\��Z�T�.5-M�F�	   �F�              !�             ���             �B�             `!�              ��}              X�>              ,�`              B�              !�             ���            �r���bUf)H�m�?�             ��������KBB�XQjj��,X`���������D�"��}             \�Z�jr��9˅�4�S��>U�zu9{����}ꋉ�6�>X�>             �B�}V
��C}�b�p�=��!�            ��X%���P�]q�_�1�             ����:�V�����"������`            �BWXa�ª\WX�K��=�         `9~>>�����������c�O�n/�׷@��7U  Ȓ��n�r+n���            `�
����Z"���%��^�         ���a�$�7���.DŊ�\������JHp����%&1)��)�u  �6�9rD��✲~ILL��V��=z���/rG�         ���5�Wq7?�9n��l��5 ��DFF���34l�PJ�����𐈈			q�������>              ,�`            Pxx�T�`?�ML�KQ���"@q��]B*����(m����            ,`t���x�6�׷�� ��^��}j�+%��֑A��J��%��'�wI)����E���L�z����(�\x"�\�v��<=kU��}Kxɸ6���m�ҨR	���4�JL��<rF�\�[6��#�            ��A�֨^R6�/�����9����eL������S�תl������~X$�®
`e��7̅k�̅2�����r%��|� �g�w�?箑Դ4�*�}            @!�ψ���L��\2�r\R�l9*{�]��ѱ�i��դg��Eo���dᣣe�G?��K���?2�4�w ���,�m� ,*�T�U&Hz6�!UJ��0�[KINI����"�            �!���Ȗ�埶���6v��G.^�/��JT|�M��\���p�)�o*��?���d� V4�Y]ӆW�e.D%$��oʆ�粭����%/�*���2���Z�ܰWN^�+"�            �R�����^��#�eZ�L��R_�*9u�x����/�ˣ��u��װb�D��;�{��+msa궃υ��$Y��X�cSR���H�ZU�m�J���!�Ԗ���+"�            �W�u���%%61I��y��+_���
���8�bv��iR���ުzE�}��W�f�uʕ*�mhv��&ا��
�"�            ��jȄ����Wm��W#��ˋs�����@_��G��rw��s��ś�m.8#اRR/qy1:V��`            �b>����>��!����|�sہ�)�{H*,ʺa&?��%���}���g�v9u{���N����e�*�}            ��=?���.WJSR����3U+h�jVN����&[N��*���T�ӹ����o/OyaP�\������EYrV��`            �B��ح�����mr���mK���4�k��y{B�Rt� Vжf%�����p �`��Ȗ�����\!�_���~�kIu�O�����f�	�Z�>            �E|����q}���C]�b�L��h��ҵ^5s9<.A���N +й�Ѹ~��B�UywE�ͅ�$+����s�Q��2oo�$�����            \䩾�I�r�R��3�����ҿq-yyH7sY�M��TΆG	`��ӗKB��悝V�{cDO� ���%.�G�            p��Uʙ0��l�n�z�ӶթNU�����z~�ZY|�� V��>�\�|��r*�@�������������-�+�����ɽ���ּ��!�l�==k�X�>            ��<=<�1}L��3ע�����������K������/���;��j;j�\xeц�FT|b�emA-kC��w���܉�L���.-d��y{BĊ�            Nv��&p���y��$$9e;mkV������C}o/�*��&�U�۱���Y�\��L�ͅ��"���Z�?�\�g�}            @qU�\i�3-M�	����~�{��r��rRJ�4x��ѢZ���	��1�?Z�C^Y�ʀ�Q�|)�S�=`���s�[���l��s�9�����O�^�ҦF%S901%E��`            �""��}��#�X"�a�2������n�<?� V�G�Brj��GBr�D'$J� ?�X�[&��            �����e��� ]�V3�/F�ʆ����-o��-xd����j�^�n��}�W�6��#�2f#�Ċ�            N6m�A��wÚ2���a�}����8�n��2oҨ�P���٫$��'�i��Ԑ9G�������]��r�6;φI�E'�>            �U/$s!��K��S��ǧ/�lP)�ʔ)#�5rʺK����x��4�kV�l�b����Md���ML�q\�Ƶ�_���_��@����            �Д��JͲ��r|r�$���;�{�z�5!ge֮#be���&ا��DFFHDD�XALLL��߂������zȢ'd�P9s-J��D�U+h¯�ז����g������bU�             7T��_�e�^rw�f�OC�V�i�/11���	.%.�ɕ�+�!����R��W�h��,�Yv����"II�nuK�}             ,�U!7����+�������E-����rk��ҹn5)����m<qN�ܰW��>*VG�            ���GNK�?phl�W�����!7��
����K�o��3υo6�3�����)WJ*H�����#Q�r!2F\�"��I�.�            (TQQQ��Tx�+����.�VX�>;�]oC|M��Tۋx�r�Y��>             ���C}v��dg��

2?�Z��� �            �PX%�f��p����p�u�            �rڎ�J!7;{���Yu5ܗ�}�a)�             ��ܬr����+а[q�_��>             .U�Bdi��G�              ��}              X�>              ,�`              B�              !�             ���             �B�             `!�              ��}              X�>              ,�`              B�              !�      �J�-)q�*	  {��>     `G�      NU��Y        �!�             ���             �B�            @iii���!�Eq�_w@�@�Wc�\	�L�O\R���<F           �/������D����T	(Y`��������%�g� y1�O��2���'�c���$2,L           ((իW��g�Z.즡�����)��oJJ������"�(.^�(+V$��h�/,,LRSS       �?��-�Z5th�C'��K��=����ڛ۞��V&o=p�ؒ�޲�����w		������,   ��ja7{��Y����P��`�b�p_��      ��u��UYu�t�ۆ4�'I))����L��;������������&wwh�e�oD�R9����#   ��*a7mG����U��P���P��s�>       (x���m��μ:I����}?,��뎝����K�r��ĕ�L���ߎ3aR�|i  pG�vsuȭ��/�`�b�p_��      ����uD:Ԫ,��m,o,ݜ~���:֮*O�^)/�"   �n�r+n���!��X�p_�r����Cp�+W�HZZ�        �#2>Q8a�}�Y�Y��w|�����"3w!�  ܞ��n�r+n���Pl%''�����f��       ���m?$#Z6����擡���!��i$���  (
\v�Jȭ��/C�         p�:%�bM�>��mTS����[�  @Q�a�#G�Hll�S����'		�b��____IL� �`         �&�SSe��rG���kd|��r>"Zք�  ��&22R�=�u7l�PJ��+��������ۊ����         ��O�ʤn-��vMdP�����풒�&    ��}  ��\�O����O��[����       @Q���E9vU^����xyɔm   @�B� �0?O�,?O�?@     �"�rpI�]6Xj�	�r��R��.~R6�OJxyJ���xzx���rBr��OLB�$��J�����X	�������Q��������"(l���*[JV,#��Z�@�`�YU�c�ϻ����2��v�]$">A�c�ψ��O]��c���m9s-ʴ�-ʦo?$/�"뎝��W"  �[5��{�I����yf��?�>��{G�&���?.�Y�E �e�Od��N_��g���>��3���`������Z�>        ��JAҪzEiV��4�Z^�V.'�˗N[$c��)�î��K���e�t�	j��i��i��ҾVes,�b;��g��O�oKã���H?�b[v�	���d)*>\�C�޸ׄd�?%}��OÚR�t�\����OIx\B�c==E���\z֯)�)�2s�QYr�D��֊�=T�zʘu�>zFB#����AK�R�cKd|b��5`ݫA)�gB�������JK׺����K���$�O�JjZ�m��լ,�kT4��7�8//\�vl	ۓӽ~uiT��D&$ʚ�g�lx���<�|��_�����+�����t�r��[���SB��^���帯-�U4�4�z���';Z�V��y?�IL�5!g�cʎ����,,Wc�l�zZ��~f�����ۨ�m����o�m_c��_�L���_C�lϩV�\w�\��f=�v�]E�<=d��0�a;?洯�tlf��D۹u֮#�8�c^���z��ڶ�_���ٙ�s 3���F�4�<����x}l�?/����}����ӹ��s�s�q���ȶ8��)H�        @&<�ݠ�t�SE:֩j�����蒑a6�5!�UG�ȡ�%�=�z֯!=\_*d�`Ι�ҟ�8Ҽ��MC.{�]�-�BeM�YYq��[�4��S
�j;>���|xl��(��_'�nڗi���f?<R}��oצ�	���'Sy���_���j��n��.�-�tS�lL���Q����o�mZ��ٹkd��5(���婾�Lx����Hyx�s��H�e���}g�&�v��^��X$'n���ᬯl��k�j�n��'D�<�כ-�U��&4;�s���%/.�pS�,/ϻ�j=����݅�yd�2��ȷ��	�h�3��j�E���k��k`����]FK��IS�������I�*��o��R����������ג���3ϩ��{^Y�ф�n�`��Ґ�&�hw):N����T��H�3_�M��҄���]�?��X��f[����nV7��zN|h�b	���i;�'�0x�Ƶid��>�n^��^���<ҽ���j�p��2c�a�8u�䐫����)Ȕz�p\_�|p��F���\�}�b��=Q9|��
�       P�i�K�j2�I�ߤ�i�j5Z�jd�fQ�zt����x�q�p�<�{-D�tcZ72�U^�e8�`��.��4����e��7T\i�c�C5.��5g�Q9�{�ʅ�����}��߻���Vg�N��)\�aSmז1�4��ޘ>&|���C�6e�����VK[��]��/�o�y0�7U���?ݯ�	�i��n��ܫ᲌A4�A�On�oBo��K���~��[;��X4L;Ӷ]�qc�a.��3#��:o�(��Δ������<<BW.w���Z�7�i���?(���;q��2��ι?�lc{~=�sפߞ��]iɗ�v���k2�O�d��3d癋鷿o[GƖ�vZqvޤ���ݩ����c���y�F��^���ͬ_+*�`;��|�ό�u�@��
��<�vwN�h�����ۺK�m�~�ao����75��i(��{�m��6��^�C����z��}�����
�������ߨG���Ǎ����/���=G7����u�c��혷T��|�G���ꫬa��1�י+o���.�ʗ6aQ��qI��P|lZ'�\�����6�����ЩNUs����	��@炶�U���?����N$�       @1�ّ���ʨVdx�7��N[�i�C�h5{�Q�������Ӏ���eL�FYd�H��h�J�wF]�\6c�a���Pz��U&M[���5Е1ԕ�GZ&��m�k�{H�A3?�ӯ�BQ��vS�,#���y���QV�>�
�s�V��`�s�:�����>mM�7{���ۺ��ӛ�=��,�w̄3�z�S}�g�n������2�ۅ�z�ZU���i0����߂��th�e��N�y��M����C}=ܵ�|�n�yT^�� oyn`�l�j��!��Og��Z90�P���ğ��V^X��\�rN�,�n��v^8l���w��/'�o&�[�K�^�*���|����� .2��ޥ-�u��ώ�:_��2�5<�@�[�����'�u=L7�y�,C}v���}�f������e��N��'m��;+����L��Iuo����/�{����wܚ���p�K���v��`�{ƻ�{��ZE3��>��ߠ����[�v���t.��a.L+���;#�       @1��k+�{;5��2ѝi���:57��X����� �Ɩ�(xZF�����	��+N٫��8��,9pR~ܲ_~=|*�R܃�>��֛n�0�GȀg��l�L,'�~��L���U%�m�l� =�ׯQ��j�K��i`L[��v>�J|�*�5U��֭�k[ž���q�A�>�jJn��ڃ}}ג��������2^C|��V��y}�;֮�c@R��û�	��m��c�}���9����N��~}�u���P��#s��_jU6����[��65*���+1q����f������rv�������>7#Z60��ֶ���1��U+0iX�Z� Y���ڳk���Q����~���'����	k�Jm�]����ZU+������_+C����:��T�m.��6���`        �@�*���mLK#�\>|wg�yap����睇��;���+���ǏG������ܣ:_^h�J���h5�)��������uiհ�n���5�φ}:K�|s���*˩�]I��c5k�����|��@����ݔ_��1k[�`���>Ƒ�C�C�����L�x,��6���<�k^�������d{L��2��}p�������q��+���1�T�1���U;�瀎7��2��A]L�&{{h���^�����^Z��T8�O�O��c�>=k%s	n�[��rw����/�m.�        E����k�v�����"C�g��7���5��O�����ڐ��?N�S���Ǔ��-t?����{�6U��[�]�]m-جJ9S�e��0�MLJ��V3��K[���� ݹ�(���?.�jwG.^3�/��JM��?X�t-�~zY[����ū���k�����cxP+Gڏ���SNN]�0�>u�R��fX�^�K��L�m���>'�������������;<�H�1�:�ڤ���^
7�r�u�'�b�s��Ǉ8pn�NH���ѿ=���>����k*E���o����8b�����fus��Am�<wOH�۵m�V,<s-ʄ��@χ��k�N�v��|�aO�֧sD[���N����p:>�a.�/�ʭ�/��+񶿋2���.�       P5�R^���޴�+�L[�Ƶ̲�d������y����6����L;��HWZ=DâK���~�"�O�	\G[�j�ap�@�~8�֯[录�LL?�͍��ݳ�Q2u�A�S�[����I9�[�����-���Xm����ӯ�i�m|���]��ǯ����e��#rG�&َ��7$=ȴ��S��I�rَ�fӾ��sv�ȋ�����َ߸7�������=�0�~0�ϝ��kN���W#e��S��������T�tȡ�w��Ij������Wc��`Kv2��[��n�Lտ�$�����v���B9;�be�o-�5����W�l�o8~.=Lg��#�M���L�zЄ@ղC���T5��a��@����i�m�T�C}.�>Y�K���V�^|�}�Χ�ån��َ� �V۱�s����2�%�T���5���R�B�c���Jd�����l���������ܑo��ΟH�{�_g��]<?������;Ԍo��u�����$$�f������4��b�o_��2�}        !ڪH�t��~�������Y�����h�
�*Ȟ?�[5��cX�8�@���u��������u&��
����F�d���5��	���p�iז�@7,*�\���>mkVʲ�������ӯ�o�Nޢ�tʦ�ݧkv�����~�~�	�eU�L[">4e�	���c�ZiU��4�"�r)\���*������D�M�e�MO�ޙ~]��M��T��gp�����v����V�yu�F6��~����+2��~�r�TW��ō4�������<�j��e�s��,+�j0�e[2m��)Ke�}C�/���_oܛ�z����F^���L}����&S�Y��H/۾�ӱ�M��J���z�ٽ�d�t����r#m��ȴe�n{|�rY��S��F;΄�ˋ6�_�����X~~pxzK܌���O�`jkϧf������)Ȩ�H�C{�]J��S�q1�E�l�y=�w���~}��se�3�|��X��<��4�Z�2�֊'._��ڢt�C�3�\<�Imi��8���O�J��jW��	�w�o�C�H~��'�/�<g{_an�]�����>��o.���'����u�[���}T�@`e�        (�u�_z��'���^��ipch�z��V����L�5�PF��Sz�P9���c�����ƽ�RǑ�L��2��t��lc��i +��nӶ����:}�}<Ӝ;ǵi$5�˅�h������l�	�e4��奡]M�� _S��rT���p}�
vJp�[(ui!�vj.�msJ}�:)�/�l��e�����y�o;�Ӗ�ڶvΞ��[L奌��^��N���Ѵ��v��.]�������Tڎ�����[;H��5���>���%�d�.V���˷���s���t�کV��|2���{h�Yw�yn�qtB�m_O��}�1����]���ݩ���w�!��JT✲������T�~]�^�ڞ�i�L���e�n7���|i�����}�ʒf�����AV-����r�\؏K��<rZ�c������Β�l���H�r����}�m��Y.Egn'��y����3�;�m�ԓJA%M[��;�{+��0_F�8t��m�ڷQMX8t�|�a��`�i7;����}�_{�T��	�i��wWn3�׍��qpy�k�ߏy�c��?n=�i�I��l�ڷ��=��}��R���7�B/�}?,���/��dG�Ǻc�L���1}��2�aϗmsR�?���q�Ѹ�A[}�zwŶ|�/��G���\���[���υ~f.��h~���?}�����1�2_�{����n5D?�Q2�3MEY�"�       ���𕶨̪���a��:57�M���V~�yD ��c*�=Ե�i���y{yʤn-MU���;��A�i7'�A�V��p�ylگ��1��x�iu��~Y��6m�U�tqĿ�7�#4Ԥ�1]��(/���,��؟��*��{����v���<iGh���∼>�aQ��Y+��}����qԪ�g����L�1̙hHPGh��g�6�#�^�&N^,��0��/�:<�E�����Ǥ�N�>�9�qR�Өf�!\/>��2ӊ�u���V�f;?h(�ޢp���Ti����syB>[��v[�R*�̡'f�����RC����<�sA+�.>p���t#���vMM�y���?Pڿ�C���,�        pSZ���a����h��i��/�4��3��6�ŕV	{mx� �=�>�k��۱�L��4S�R�_V!�U�~�j�I+�i�a��3�z5(5m�!yc�f*+o*�6U�&thjZJkv������&��*�.��X&�ׄ
wѴJ9�k����g�v˦��k�U�Ʒoj.�{ɦ�*�V��>�����)���_m؛����F+�j��9�4A��e�e\���v+"�       �j[���.P�\)A��lPC6=3A^�e�|�nW��rR��W��Sno�X�?]�U�oZ<�ɱ�e�NÑ��T5�S��^�}�/��N�r�*���3�rφG�ĩKm��*��� ��6��Z�^^�e��𗘄DS�0�Ј�\ף!�k�	��5����������:$`%Z5���ZL�^]�1_���.a*w�|4��5�pz��p\�����"Ǫ���!geƎCrG�&�����	�       ����&vk%��f>�F��F�-S�F�L{��1R��k\K>�״nC�� �~`߫A��̕r-6^�==��l;����yݱ���r>"Z~�q�T#ʎw����w�� k� �V��ʞs����p��C;�y{���ὧc3�N^��JC�m�//.\o����߹yz�'^!1	��>ݯ��)WJ�RR�i�$95U w����լl.�uf��B^���=�״Jy�*�}        �	���mc�7�%p��{�.yx�Yq�E��>����m��#Z6�v�*˟~X\ mŊ�wF���8�V���d�i�;u�Aڼ�lZ�q
zf�j�pEP�m�?1c��~x���t#࿰`�����v��{m�;�[KiV����l�'XB�r׃����Մ�َ��v�n{O<��DsY|^�����|�J����|2|!hl�F2��z��k������Z���+��\��f'�\�a.$��B�s!��³]� ?�*�}        ���n��C�Q���+�/3!��./�������������KNW�t�	��e�r���� ��*Ȅ�هK�J�#�[ɛ˶���-��������4�Si5��m�_� E��c�d�'��͑=�U���6}O^z�<=k�	�i��go��:4rwǦ��FZ��:�
wi_��ju[�X�eEۚ:�>�^fQq��p�?:��.��~��m�	�       `q��������}p�����m�Y��2q��ZZ�j��wG�6m�������U�/-o,�$E(#�o��6�,�1uL�O�������R1��i�I�c�xЪ�Z��Z� ��/��Ff���n����wVF�lH���7����}4�q��K�j��ŨX�p����r�[O]�\�J��e��M�J�Ρ�g���K�q�}�W
t.�U��U�/��P��j�W        6�E}����U5�z��x�w��_͓CaW��َ�7F���:5�����޿�ԯPZ��L�SZ�%��ge2�SR�$4"Z ?�£�r�*�s�o�ҹ�\aڶ�f�M�5e����L�B/�}?,�r�'kv�'lw|���������!g����09:z5�!s&�4���0�"��Ǵj�[u�X�>        ,������Q���Ñ:p�Ze�eɟ�ʽ��"��Z����h��)����*

��VM{�1_Ε��D)�_	�u̱� 9q$�{>�@0�ʖ-+�5rʺK���xkU .n�[�F���^~��D�%d;�|��|=aPz(\�p����bU�        ��{;6�wF�2}֡��~h��}�j�j�^qͫ����&UKQ��*���L�q4��}s���KC���)��a�u?h`���wɱ��G������ҥK��yۈ���ܿl�
���R�L�8Kdd�DD�/N��ss�pl_Y���l>y^�\���$IKK���%�k�j2�Mc	���o�Wm����        �z��-�ߑ�	�Y����b��@���beC�ד/�U|��ҡV�����脢��\���۩�iE���z�|�q�\���ǧ/�/��2�3y���'D  ''�D��n��v���돝�60�5�1�Y]S��Zl�,9xRN_� ֣����$�o'((X��D""
7ܧ���D��]\���L˄ZI_oצ�Yr���j�;>^�S��`        2�u#ykd/�����IXd���%g�EJLB���%HrJ�	0%$�H�m\� ?)[�Oj�	�:�J��}Kx��x�_{���^e��j&uo%������8k��aW���p	��5�=~�8�IL�X�e;�*�6ZU�K�V�u˗�z�KI�RAn3w2V�+��go�h��z5�!�uj.�?�-�w5m4�9��t�[M�<=��k�5��M�Q@�{�׭r1*N��I*�ۮ�W�'�Z��84��Ѹ�R���m���Ty�vyu�F���9Pl�*�gl~V��U�>;3���[����h�ҰR�l���'%�q��!��]�#�       �E�k\K>���ۄ��GD��3a���E�S+���Ĕ�<�K�<�*��V�+J���{��Ұ��ZP����]B�񫤤Z#�ǎC���tm8q^6�����.\��s�:n�Z�G�hP�F� �*�M`���|�	�5��ս)�g�����0P~<C6���>�e�ޞ�&� y���}����ҠbY�����x��U'���ۻ��W标?�ַ��ΊmX��#�������
�.��ա>��
��:�gg�J��Yu��s�ӵ�����e�8�_�%��G"�̿U��I)��.�       `B����7}�l%���d���mݖ��r!2��֭a��W�2e�As[���ҿqmzK=�٠��Y���]훘0ك��D��x\?��]�*��P+c,�\~�B���T���`Ʀ��b�!{ԯ!�֖>k����>�R���?��L��T���{����l�X��	�)=������y�Ѕ+7ݮmzs����{L�X ���B}v����u���V����Y�_. �­U%-%Y����      �ڴe����H���X����2k�QY|���8�Ҷ��a�~�h���-����J�:U�J�qyy���_dZ��}r{��mc��CaW��-l��S�ѕ���.Z�I�حMj���e@�:ٶ�r�;l��a�s�n�ղZ�\�h��� g��M�ΉV�ժ~�� ���Cnv�
����C�@��,��q'�`      �L��hk�j���.T[���{���;+i�2����BL[�N���T��H�����ɗ�����-���0P��RO�D_�;���l��b��I2g�Q�hEȻ�5��;�b�v�/�"'�D�l�c+*�b���>�� �'_o/�ύ�`V	��i���v�wN�͊���Y�5�� p���?X�=S$҃     ���:�{�Ud\%,*V>\�C�l= Wc�Ū�\�&��R^]�Q��B��ZJ���Ò-HTB�<1c��ڞ��{�Ȁ&��*�e�W��g�v�5GZ�����;dt���d�Ҹr�B{<���Ƿ���K�ޢ��l<q^6����� 8���=��(f����Y-�f��Zu��>X�> ���<�(�e��     �������][�Ð�Q�������ƽ��,�BCco.�bd�ӥ�o�V۹�C3�IH�g�q�������L����H�����'�ϗp��ܴ�d���2�uCyap�^H4�Z��w��Lu�������U�6�e*�fE���
_n�+���߳����� ��7+���||
��CV�_???I�B�v�#�       @!Ъ1Z��#��pN�l��u�|�~�[��"��%���{���]���M
�y�Խ�����V�p�6t�>�7�jh���5��U��ݷ�FjZ�	���{L������P(��T(#��&O�Z%�N[0O��T>��7��\v�<>}� �+hE���*�/U��ĕyt�2�z�-D�FhyD�       �B���>R&��ж?g�QSUNۑ�/��-��6�=�}�I!�U}iH7S	Q+�9�˶��ٮ��Ĕ�x�Nyw�6��/:5ⓒM�A�&���n����1<й�,;xR��wѢZy�K3���em�Y�|����l8~NƵi$�*�5Ǌ�ۊ#� \%95U&|�P&th*��7�:�Jɕ�8Y��iɮ_�ꢝ�T��e���=|ݱsR�� ��>        \L?T�������Hyf�*Y�F����z��|w�<շ�Y|��\��W��'aQ����LO�j#�ۖ´��y���+�p�U)���ӰOg�C]Z�
z�%\w��������ۓM@���r��9��xy�^*S��uj.#��+�.\qjK p�Vf�~�~�ܨg���r�V��{v����  P�       �B��Kʿ�u/�m��{L�iY�����&����2gO�|=~�4����}Z��ۻI����K�
d�w�kb�=v��p�|�i��Nb�����-[O��ww��e�]��
���戞r���ʴ��[#{�g����
��"]�;��I �"=�Mඛ��J���w���k���	  \�`        .�Ґ�R��ץیON��]#_o�+ōV
���t�ψrw�f.߾��S�4Ԅ���_~�k\K>�W��O��V�{p�9%���3��{�LPS�:�ʈ���mޮ	9+V�H�VY����W(-��Ց��b X�+C��ʪ��7������IJj1H� ,�`        .ҡVצ�K���w��n��9wI����$y|�rӢW+�����jP��	���r�h���'����j��?\�C��x�$��Jqu-6^�~9O>���m7r�vߴ��ޞ"ɩ�|�[V����} �H�kW�qL�R�rK�
���E ���       �Z��Q=]Zmm��K2拹+�~�~9x��p��ٕz7�)/�*��`]��[�L��zh�����]�;�
v��s��-�'N]"��c���]��ƕ��}��˗��%;�L.ƁP ֦�>G�6+��j�  (�}        ����lY-��Ve��sr�7�%2>Q�;��������o�fUʻtۏ�jc*'��y���h�`ƃ�]DT�C/ێ�r�j��wii"���V�S��	�k�
��If�:b�Z���Q��9�!
���"cLe� ���.  ��>        ����C�1��˶�p�1y�����"�YhD��d�L��0�\�����c�ȁWLh.7�2������m��mS��̄��-\'����η8}[e������k�j>X�Cƶn$%}��h�ou� +J���4}�aS5;����3ע  W#�       ���޶�4�P�%�ZrV���b�A5�� #?�#S�*}�t�v�"��6U#l�!;�����K�z���>^�S�_��T�C���yz�*�\R5�����߹���|�\�Xվ��e�w��	�L�_��m9jZ9s,��-\/jU��U���;�2�3�  ��`        N��'z�uɶv��(w}��P��ⓒ厯��w�rI0ˮn���ٝ���*5��Ӌ��ʘ����[�]^\�^�}���D�<6V�Wunkg�>ܭ���t�X��#����˸6��E�
��$kC��/��g{��Uh�~��3�~̗1*�/ ��sT^[�I¢b ��@�        'ش�KZ��\
��_͕�D��SRLE1m����}�֑g����,�r���_z�&j���&O�\)�m�'ț��$������;�\I�nkb�����f�����6�}S�]6Xb�d����}�g�vP�x{yJIo)��+��%�[����JL<��n$*>Q^X��,>^^��;�^R�T�D��\��  \�`        N�x��N�Flb���v�\����?B+��f��~x�t�S�e����e�ً&e����[\I��˟3ע�i��?�f�t:�����C3���]RX��J^�MJxz��vg�&���YS�R�/�F�X�ս�BK�`?)����՘�|��mύ�XIT!�4�׬Jyi[����^I�W(-5�I��@���~�ke��1r�J�
�*/\�-'C��ūnѢ�f�`X�Ʌ�h�/b���>l�2���F��}=Z���y~�:�t�  �l�        p�&��I��՜��'^!�î
����d����1.���4,��]��{����z��C"M�%O�&�W4���ƽ�@�[����z�����6U]��Z���Y��[���Ѹ~r�����Դ�|9~���W=#�?�-���ؾ2�e��?;g�|��*���Y(-�s��=���U.ٖ_	/��vliV�TYՐW���]Bj�+e����j8qM�YY���,=t���A�2���w�:��k���;��	��E����U�e��]��2�(�������) ���       �$�tl��m|�y�L�qX�Z�k�W�d���JU�P��W&�7D��D��?L��]���?殖�6���lP�T�r�ꥃ�W���(ɭE�m-�0��Kפ(�^��yΆG�l�z�Њ�p���%��.-L[��Nz/ж���E��.�w̼�k�/�"���wh�ظvM�d����o
��i����֯g^?  ��`        N�[�Kno�ة��*}��ZPpN_����[(s'�4��+h{�5��\��e[�Uͫ��~�;��4�Z>���q&L����P��eE�n����`�h����ַ������U%�q�kW.��>��yg���֯[]��1��
rpmɬa�Gz�v�s��5�Z54�Ν�Wn������-�j�����[�����(ۦQ���Z*P�֭&+��  ��`        Npk��R6��i��Bu�i!�����y�������]�MW��~�yD^_�I�@}�u�V�+����ȡW�*�;'3wqjӡ��6��n���@Z�C\�J�0�Ѯ��w�VqUq���78�VC|wtoS��0i�Kmi����_6Ȍ���0
��mT3O����M�T�O�uU�sW�L�  �L�        pm��L?�:,kC�
�c�փҢj�Խ�5����G�-�t{o��U���tm(���[#���1���ϻ��h�@~ز_\E���g¤S휫�m?}A��z�KK�ZUd��P�o�q���P�Z�KC��Į-�Ze3�����w��m��/�|��ˋѭ��^|iK��/E�JŠ�ǅE�  �D�       ���]B4���G'$���_'p��毕��H�Ƶ�����ٻ����G:
���Q��{�ǖ��6[��l�n��MO6�W[,����;@Q�~��t��sg���=�<���)̽w���yS���ˑ�_ �N��|�� �گ�f�!�`-�n����\���)�&]EU1�}�E�}Sڱ�O5]���ܥa`�V��щɈM����H0\五�l8�U����
�J@������RaЊ
1���y�pŠ����x�:cX�F���Xz�$�����Y��?� ��n޼�jժF��j��0�GDDDDDDDDDDdf}C�k��%�[��4��h-��&�����^�u7�s1���H���֪��M{U(D��ܝ� Ε���Uѧ����xip�ە��7�l"��e���-C�¢-��p$���&��-:xg��Y�>e;37W,xlZ���g.��cɡXv���+���}v���`o��4:6ܫ�mB�d_�&Ui��L��7������*�y;i0}a�fd�䂈�233�����S	�U�^���[ W�����}DDDDDDDDDDDf�?\��7	e}���2����bݳ���[%!�'Y���+ ː}���{��Ю�ܾ]�j�դ�l��C�sZ,S;4U-d���Xs��C^A�l�<����;��Ʒ��a��c�ݷ4���j�qYʬ��1���FZu�>2�ܡ��/��~�����_N���#'��/�nT�h��z�OL-eofn�����p<���������||8��{�.�ߋ���F?"2��u������I�/=��Y�}B�Ϸ��|�U����>"""""""""""3��$H���|�6�Yر���>g-fL
[-��ߦ��i�,�۝���5��	�x�O�x/,ڌ�bvT,^�U�)o'�x��M.e����1�;���5�j�@���[��2����1cO4
$mF2�W0�������	mB�nc��2��L�E_Z�o��n��O�d�����=�,$�7����pC#�딒������Ha��V����`�5���kjr�2��mA�'Ko�ۃ�w���w.	���	���Y9��'������������+c6G�l�F']�����T��*�[$ܳ��yՐx;�.��]�cn�ش��e�	WT��*晞��ܲ�?w	�~^�x�>q9�g��Ǜ���fO#ۙ�L�`:H����L��ߡQ�1�WV�れa����a]w�ޘ�vDd>z	�Y*�V՞/�������������̨K�@�n[ڙ���Y�[kv�y�7�D4���1���R�C�u|��lk$  ��IDAT� ��R�A�����~^��X���9G��uK\?0<X��i%r��Q���m4�'-eҴ���(�ߧܮ����e?�>���Z���Ne��1.��_���<X�4���r�گ>����X����ol����S��9{cM���<�y���P��1�O}�az�V�vsUםJN��wa�~�7�UV��Y:�V՞/U�}DDTn���W��ȫf�Cײ@DDDDDDDdM�������Y���{|������Ն-���8k��)2M~���ǣoh}Mn�W㺚�^��P_!	����*����I�XV��X�I��5	�ɘ_c$H9o��{����	���X���H�F���E�#�l"~|`0|ܪ[�~�6k��&�ω�u�&��#S��߾i��I3�דb�m�ǆޞ�f� 5���M�@D�a����BnU��R�0�GDD�v�����)՜q�Z"����������C��&�+�0Q��֖���)?,Æ�&�艴*-<xd}�^��}-��B+��O�д�u���o��]�[!%�`���e�'�n	c�K��7ZmWG�a{kI�c��2vW��Z3�WHF;�l����b�)�M9s%��\T_˾.u��3�Ec�u�f5���޼����^�ˎ�R�jDd��Y;�f��[PP�7������l�SK�ۖ`�͛ 8q9�g�����=JL���/�҇��O�P����à����0?/5��4���㗯���m4�'��Ϝ��)&�����hP�ɸ�w.uy}�p\ON�O`2;/_�&Hcd�w� ����v2go��`_u'G�n�?�>��b|��R�;��aL�&xw]$��|,v�Kȭ�=_*�������������$̯�fA�_�yMOV=�7F�O}�A�d﵌,�>d��aM̙R����g5��ަ��G�;�t��(nym��x����w!!��m.K���u�gA�'���:��-�y�N_DU%AR{;�'0�?.(n��K�I�b��*��)�W�ӽ�u��*{"�8	����!3S�൓�rr�����8~�x�y�T6�������������Dڭ� �kU��ּ�r'���_�6#V�0VE����س��$��ķ�&$���%�s5#����\GƗ�_KCU1;*/�z�������,��7�����es�w^A�{ln�:F��\��o�ك�쾶a&����WR�~�c�ϐ.FF�K V������2�IJ+{"�;iii*즅��88�C/�U����T�8qB�����1�GDDDDDDDDDDd&aFZ��a��s �)�y��Z�M����kB�g��?˷Ö4����?|�2�nñ���J�V��ޚ�d�{�#����&����UjL��$}ip��f��75K�or;�!��Q1���������)�QUui�&>�L.�mb��}�_�:�l����/����)K����`�����6!""���#""""""""""2��]�N^����W�ۣ{����BSm�g���q�������Ӭ��ջTã��8���=�@�Bzv�Ю��=��W���-�WP�t٩���h3r�-�~&#T����m��n\J(�^}�e��P��lS"�(�qo��e2�SY���!.��4u�		B��5�i��>i�3f߹$�&^�_��`5ڸ4?�>��lj��&��h�Ň��Rӱ��95��	���rg�h���Im�ѵQ���_n;�#��&2y��u�7g'$ޟ2rrAD���>"""""""""""3�[�]���~�r��-c��bK�7��϶�Zx`��Kxg��sPgX�~��q�*�ݣI=L���*����n�m��z�}ǰ��EX���$M�}&ӊ4Q�{�6��c864Q�ߋ����@N\NAU432�h�O��&�	����֡&�h�,Gӿ�Q�2�^��UUgG��~#�˗>���l�˥��T�O�}C��:�l��_��v	�;�;��o
�[�hzv�[��m�"s�*��jS�}��D�u�r�����={b�0��:��bا��UH����vL�Wc����Q�x��M&�q@Gj� %A�A�̃1�GDDDDDDDDDDd&u=�����Ù+�����m��i�g�R�6�Š��6��j�����k�����
�e�4�=�1���a��Pt�u!`��S���Vu�;�Mn~O��)&���������O�-�Bg�VG�FU6�e��e�/{K�.9t��e�6d{��>!-g��ۀ���@S/��o^���ӈ�I�[�1�W����\5��W����4 =��OWg5�[.+�����M�>�}atOx�p-��Z�B�Z�hU׷�����	�b�������������$��V��{297+6b�,O�|��`6�q"��+��y��a��� };xA�f0i��R�@V���ai-^�]�
��ᱮ-�XV�����U\�@_40����IղD�\ۣD0Ƙ��ϡ*+m���W��'37K�����F��h o7W]&*JB%�OZ�I����G�*��e����=9�=��r~�Ͱ�F�M�����u�5
Դ���U2�W�]ǁ��;����˭`��CǡW���gugh��:YEG]ڢC.c�cj�%��/�ҿ��ڴoj���do����I�J�v^��g���*�v&�x����vM�*�7�D8J̊�ފj�S�r���>������':�\����r����7�d�O�!2^���PYHP�����6��O�X��yX!��Ր���IS�9��w//i���ఢP��,}j�Z�]�vǺ�G(� 1���H���^!�G����Wo�٭.e����.�~ƞh��}DDDDDDDDDDDf�����Jcَ����}m�`�Ҿ7��ABj:H��qM��<\�{���ZC�©����qG�O�����U�֪H�`d4������!��ҭ�ٯ����C�.��{c\<�b��{���b�u�e堪�ҡi��Us�Ɩ�v�-���4ԯ]���:DT�`_�`�~xx�1��f:�{+L�~v�b��=97xlo���gG�T(��D�V�1V�x��\����i��Jz%-z������}f�é������I�R�?k`���������������)t!��-[r�J*v���ZP,A���V9U��3��BZz\L~�7�j��C���\��`�섉�-EU53*��~��2Bq`�Xr�D�ok`�`��������d���B��r#'����֫�^��ī���QZ�����&$�붤�P���گ���~mU�Wס���z�m��B��|p(ڿ�s�;L���nj<n��X�������C��g{�V_�>����f=' �$i����2���y�M����#���i�Q��}DDDDDDDDDDDf �-���l��#'-�[|�D��.d}�ا;3�Dvi�F���{��������C�����e�ۅW(�7�}S��f�t��������f1�ƞ-������Χ\GU�'$H�&L�Y�mn�a}�o{��2��փ}S;4U�>S$�7�c3��>Dգq]���V��Օ;UfE�}}C����}zי�6��Q�խ����++v�?�2w�O��z6������Ǽ�Ǡg�����6�W3�9'.]��}K���S�J��������Ѿ�u��H�OF�UE��3�6��D4�cY����u��Z5�"�����>��8S*i�*MR9^�ʪ� �����@\�n�dr
��Ѿ~��Ƿſ�nCV�S�M�z~e��6��u�n��耏��U�Xُ��~�·Q<h����$|��섴�l]����/�Q��������ぎE�v_u���V�#""""""""""23�j
1�g{.[��!���H;Z��e��UTtr�SUC}�fF���{��6��t��2ocB�0��!mN���tq*uyrz��I��`#�l�u�g�*�8go��`_�}.<x��<Ǻ�~<���A��塚�d��݄�Z��-�:�l"���P���1!��U�I6�#	�U��[rT/���T)sG�EUN������c�����������������5l��oY�W�m�������̭�{�&`߹�R[�>�z U���Ӫ���~?�}�r�&�3z}Vn�� ��I�Oi2�ߪhB�P�1e��ػ�����ƈ&o[Zm9ط�Lƴ
)u�]�@T��`z�V����G!&��P�1�<���/(���&���W�u���y���<ܹ9&}�/pd/�4��ﮋ�዗5��^M�T�VH�}��x��}DDDDDDDDDDDf��x9Wg�m	�e��jU�d[���x��̭����ȌUX2}��r�c��;�`v��Uf��8<�ۇ�Ņ��B�@�`��i	NF�{]&�Jl�{.e�k9�o�{H��O;��拋��3iKÛ���Uѧ��vS۪]G�hlty�� z��B�uآ�1x�w[�{�]��v?�>��r������6�ؤ��`C�]�VM��������h�S����j�HSi���#i���s�a;^<}4z}8g���Țd_�dB?�/�]���a_(��~��>9��;������������� K��O�lΨ�M,v_Ú7���-*PA��U�`��,��;}%�ߟ��{����`��8�������9	�eƞh��>1�}S�����Njnr�,'�}-�U�W��$�c�������l���}2.\�)��������.�/W��.������,�6���s�v* .��?�]��K�����%�w-#��Z��K6�}�q/?1Z�����#�\"k*�/����d,��f����c#�Y��A�F�>6�ٖP��h]��"�4����F�m�bT������&P"���W�T2�hB�g�2���q�B��ې���2�t\k�=�]���'�C�dLޕY���ޗ4�98�n�t,eme5�C�R���{o!�����rz&|�\�.��.ﭏT������dtxg&�G��u �QiC��ٹ */	1I�I|������1β?��ֳB�X���P�8����xW?3^{6��޻8���E������}a��F���&.����:}Q��������������� ]����5`IYy��$�&�4/�s`'�A�%=Թ���kɱ��Fd�Z�q��x/��G렌����{��A� T�~7+2�h�����Ã��H�ᐈ��=��������^]�kb�@��񧺓�����U+�'�	��"��{		y?^����h�l��N��y�"l����qH]���^�'㯦��;��6e�t�~�&�����)���8u]�����g���B�\?��O������xm��DR<�>#2���>"""""""""""3H�������%������-	���>���k?��_Û7��ɇb��~�b��������}j�[E8�۩���#�*J嶝<����m2Rv�Yˆ!e��\��FǟBvj��\��%��ܽ����͚� �E���+ú��o7�]��`��1����1��,3'0�n.�C����*hjʜ��f	��
�����t�O~�m�����w߹$\�������vAu��Z��,m�r.T����2Ή�Λ
�}auj��d_�쯾���j�VZ��U���s��`��������������r�ԇ�P2&�ϲ�IH��*F�<����m}��ê�:5�Z���}iٶ���1�B���Aw}��g�Q�N[�QP����y���ҥ�u��7�}�
�t�jF���5Xm�G��3�; �V�*9�� ��{u�	2z[Ҥt�J*��H�>��t����6��2���1�蛻�t�WEH�(:�j�4ft�&xa�MZ��o��i���5!\0cO���lFf�m6ג�5��T�����R��~%޽Q]�y�	�������u�u�I������<c˓��(����������mV��o��o_�Vl_�?�i|۾`��"��^|�M�Og�������������L�n���y�}uj�P{�o��d��R�3��9�Ĵ�%�]������[Ѳ�/��U�O_����6���p��l�~032�h�O�)ǵ�[]7�]�
H��(��g	�7�2��r_��ܯ3�*����  �~k-҂�K��or�<�3f����,���ȣZ6V�8[!/����J\/��#��q�,�Χg���v���\�u�}�p]cm|��W00<X}��X��qW��KJ%k��}����.�[l��{�0�GDDDDDDDDDDd&��S�ħ��o�m��Ş�4G<۳������Ю������F�>9�haHDC8ٗ���}��?���u��2��.�D�o��1�9�Xr�$�ޕ�������������2�'�[a˜1��<�Y���3�����ھ�M�����+NB�Û76�'@T��	�XT�1�>���V:YF>K W�I��5s���V}ݸ��(��(�S��,��֑�+f��ղ	<~�LN��3�5��>"""""""""""39�����M���)�����KLX�}m����Xl���O��u5�]����4���t�"�1h�C�;��-}�	�hT�&Ƭ/:x��F��թ+)�.��{k�h"H*�r���yip�t<�dK�4������enr.�:�Qỷ�Q���	���o����;�y��uw�����j�{�om�s,��uݜ�0�Y��﷜8"k(�ЫI=,zb���h��1t�}��=�6׮�`��ę� �^�	��t���?O7W腌���~���,�o֙0�ڨ���m��ͱ�bj�c���SҬ�h��>!�i�\��ۛY͈��3�;|�r�˥�G��ʾK���L���M��I��;`�j��>�]C?�T������#�֨��\P�;���w��eo��2����u�g�w�j�Bhh�&�]�Fude��Y��[��+���QUH;o���7o�}�`k�#""""""""""2�Ce��Vx/x��+dC��Θ^hS�z�o�V���g��G�U�U���#�����*�c�<��TK�IW�7>I�P�݄�a����*��Ϟ���Z��<ޓ���Z)��]����lJ��"=�d�^_�S����ղ��\զ������yۆ�u=_�p6�ёxu�N�?��M���~0�Ec����h��?��~��
��E+iiiHMM�����v��ꢅ��^�oZZ�8fM�Qt �l0��`��Ș,��`gg��Ѽ��v��vi��;D@�&�	�ʣ����q�>�k-\�����3�8�,ي���6��|�~�}T���h��>i��`\o�g��lm<���ff���k����h\�R��;9bt�&�#	��		��سл_��S=Z��DJT����'I�%	�M�n	�?5�}<ѳI=u�P�\���D���¢�X}z&����\��f͚���I�/''G���f8�yxx��+{�O��I�F�ϴ�Vd������^Ƀ^9;f!���':DDDDDDDDe���Ct���1�m?б�}:ѡ�?��z�����y��
g�u��Z�;�i4���4 ]N���C������.=;��<�ڶ$@%��o�0�t8����z�`0���;[j�oHDC8��#'?�Ѩ�������Ҿ�M�_�������v2����Q����ڒ�g����A�0ٰ��]	��R�!s��x���.�;��m�R��B��Y"�W���$䗪��B-���:5k���`�d5��>""*7=� =?6"""""""�J����I������]���R�H��Oӆ� ��ծ������]����;�:� �-=|R]�z����#�\IEv^�B�CZV�=er�1[N�ǹk�7N��Ɯ���[�\^�p��R��UFS��so�!�«�+��Ȅ޽�vN\N�_��GX/u��A}$�����:6������*�s9��m���;�X^9wu��S��_BJf6��ҡ�B[J�5�ޯ5���{�o��sw�/H��n~No�#""""""""""2�m'/�"��ls��f�u�::`�CÊ�l���`<Թ�jW#�Q��:j��z�<,�|ʭ����:����^���!�J��'�B��Y6:N��=YBc3�Ѯ-+e��~��� z&!yS���4/8�.�.N��3	��4��>�}��ܤ��!�B���꿖
�Y+�W�V�}U�}DDDDDDDDDDDf$㭲��U�������ۃ�t�7�T62�����U]_ؚ7G�T�+�	������iAZ�,������[�x�w[t2BV�.Y��!�b6�8�����p+s]��I#"��[�D��鞭M��/�~�lĕ��ߦo%c�-�)Ǎ��㠝�#���`��#����N���<�i���hM�p�M���u��ڡ�B�j*��a������������Ȍnd�bS\<5m`�ۖ�/i|u�N�e�s`�
�o鉳�=~�6�>��ư��HՓ=ZC+�g���Ky{tO<ڥE��$�3�u(zyb��U����������m_��!ӂ�cU���#xʰ�
����놑_.De!��va&�����Yk,6��o-tn`t��*����E�+]����x�c���u���oُ�W�B^A��<��+�u����	og�B*?�������������l������][���q-#d�[6)W8GϤ5L�}�?���+z�Ks5S+[OXn��o�����A~��)_o?�eVd�ܧ}��ib��v�.]�R����M�ӳI=Lh�����2�����&�K[��B}b���j*�'�th�m��H8r��}�_X��K#������}u��5 �{��P_��p�����6��0�GDDDDDDDDDDdf+��Vm8��.����g{��++v��ס�?>�4��`�-��W�w�]x�^���:*z�:��;hzkc��R�6kT�~0�yc��9����g�ɰ�r�r
"�-7N�����!��������c{�1��IWa릴/u�<<�7G�P-��H��?˶���z1�y�;B}�Ml������@DwOZ���\w;��ݪ��{�`��I���SЫI=Mn����1;2�/sT����rǌ��v��bz��8p.	s��B/d��Ǜ��y�O�6�l"�]�g��Q���f�*9��'�R�k�����[��T5�mU���r	���s����ϻ��P�f&�qsv�Oӆb��lzl���3�4kdr���\�8z
�$�E�śl3�c����Xt�8�B���Y��>�{S�Bd7��O�`���i��}�x�����"�6j8;b�C���^�͇���0��s���7�Ҳm�Ld,�����/{c-;w-��u�\-{�����K�B�����T���M	�eO�Ũ/�bj:lѸ֡�җ9���<X���
��)��*��S���_%<G ""}a������������H���+ú����&��;$�Z6�Շ����]5|;e�x�2rqt��GGb�'��������>j;����q�$���A�L����	��v׳r��/k���ѥ�����Ixb����ks�ڡi������B�(m��7�oh=�q!�:��ܵ�G<��DD�1������������4 ^ό�Ɠ�[iv��]�/"1��|^޽�V!-l9q�<Jm�2'������d�M��ԣ�w1V�"��M���X�٫i����xsd��%����Ƥor���ҭ����:F>2�"c����'��x�{�@��VS�RG?'�gbc�9X��.=rۆ]nW��k��7DA��-5$Yp�a�$����`������������H#_m;�'��TVk����L��_.T�L��=ݳ5�k�4�X�U���rԯ]��WG�||#ABi��ůH��ݻ����\ﶚ���X�[�6��0���:	<}�e?>޼Ϣ��������'�Ң���[�]�[6�,�>������d��S�۳I=<ڵ%���:M�ھ���_�!�� ֲ`�1��>1���?���c��@��q�tint��k��hB2�����`�FN_IŚ�3���ukT��j���[6�Ec�:��E��jF&}�L�]���g��OE5m���f�_��_-DZV��թY_L�Y�����L̎���ۥ�O����푔vC5W	��B�Y�y�������k��؄o����{񷅛U ^��e�ѱ�um�.1�W�H��g��\��ˣVu���F� o�		B/���!n�=�MX��,����I[���|�c�x�cp�j#փ�nDl���O;x������5�1��ǉ���#""""""""""Ґ��i=���;a�$l>n��z�A����j�@�CY���`�O+p��HU	L}�1J�,�m�<6
c�^����iߚ��P�as�r�]璋�Ʒş��Cx/��዗��H,>tTyI������8-a�mƵ�,�пc��Բ�n�B~�BJ:�n =;�y�p��C'GT7\j�8���~�����F'\��r��V�[S�\I��@佒�����xWӁJi�K�O2�_o?�ov2��5��D���1�GDDDDDDDDDD������\�����>��0c�P�t>��݅N����!pv�����a�zl=q���_]���*�a)������G�&,i��@�4�����}���U�!�D����_��5����}J����G�H��\�[��d��͊�&>�4�6�c���S���6�UA��������������ղ1��h32rraiC�5³�ڠU]_�~�;�ƻ��`י�$""�4������������4$���l�?9V��qwq�/�G������
�P���I��%IXcvT��e�$���UX��	�m��$��O�Ø��bj:�|�3�+F�lb���~�a����<߷�����	�cN��E�I���ׇs�ߑ=0�B�ri$���x{�r��K#�4ϖf��cЃ�����at����
�͊4���tT�"��w�;$O�Y������#"����>"""""""""""�m?y돝E����R]Ow�}dF~�PW����ƧZ:Է��	��jW���H��X��}�ΰ	�~f<�~�q���J�|���c�����||�� �dR��RG��h�Ɇu��d+��Lt��_m;�׆wW#�---+3�ŗ��p�jZ�~���ap��3�\�c�&]��<H{���L��e�%�}���������6ùC�DDdi�Y���w����R0f�"�K����!9=d��������p�����/��kT+_Y�_���&sQj`����rǆ��ã3WcU�i�qӻ�Ŀu���}�i��B%�^5�\���V."=�ѫ}?�E��wo�F�ʸ{���Ė��@<��mߍ)�K�;Ogms�XZ��s�@4��ĩ��<��;F�Rvqt��6��p�^Y�}DDDDDDDDDDD m9�P#k�y��M�����g�Jz�ss�3��j�$i����2d���g6���_K���Q=aI2
q���ϥ[��V}������[�=,v	���`c��j9�A��@{�'e�)���y�f�����{��$^)���%5+[���u&A]�1u@X0�5o����^��o�|�ul=q��[i�|�!���5�`xI(el��艴Ή�A7�봪�k�`_#�Ze��[DDD��`����j'�5kh�ѯau����q���%8i���NZ�^�Otki�����S���i\�b�A��y���`I||sdti�g�Gj��a[ �w_�բ��+v�u���V=��K+�8���G	Y������Q_.����[�.U����?�.BF�˘�Fޞ�[����}ݪ���ܝ��:��*cue|��r%�-�u%()�ٕ�mӍ7ܶ�ہV��Y�H+���%��Ouj��������9��Q��`��ȇﯬܩ�R����럻O�s���LZ���:}C�[��e��s�c߹�����-ڄF�׳G㺰�-#"�[mG�.\FUu+���uma���<��_��B�dt�N�52�]Jي�'ATYH۞\�rY{K]gM�P��ا>�G}-����%1�GDDDDDDDDDDdA_m;��-��c��E������WW�����*j]��M�^V��w�G�=ݭ��L�iV==�~�(�Tk���Z'?۲�7Q�H0��)��?̲�м�꼩�_�4�M�n��[5�U�����"c�}�n;Q��v���������嫢OW�?� ""�`������������Ȃ$����u����pq���}JӘ�mS�Z���c �JBFOtm�W�w���e~׷[p �]��,�u-#c�^��ώ���,�ٰ��:�&�	�ӿ��2�}j���0�*�]���.A�d,��V��p۠:�i8�E�'�B�u�Nl�)�Ko�ddce�i|�yR8ڙ�tB�&��j!��<���+�^��Ҙ�gù�50�GDDDDDDDDDDdaq����5���!],z�2R�c� �a�:���#�z{�����F��z�<���V�9�EF@��z�j�6Fkh�����q�j����Ee5�]8��n�N�o	���>��ܵ��RȮZ5|3e ƴ
)����;�xc|���W�4%"��u��'��D����$�.m�rn6�˅h�Vu}�[��ݧp29DDD��`�|�iG4D��u,z�~����##0cO4^^��镫����O�l���G�}r��%L�~����~۱�Wp���Ոeg�4����<�1o�ٍ�v5k���j�8��1�U;�5HX�љ��f[5�{���₽<����YJ��:���Ԯ�Rt]����L��������K�BDD��YA^A�
gm��DԩY���?�CS�����=��&'��4K��F�J#�5����	�.Q#J�"m�SX��Z�Oȶ��>*!#��ƞ���0�#�[e�,���[m�%��-J]޵Q "��q4!DDZ���-�+�do�O����������͛7Q�Z5TU�������ܦ�;B�\� ˨戙�m�vQՒ�vO�^�_���Y����6�����܉%�N�d뚄�^�}C�[���bj:F���gh~_�����)����צ��=:{�����69�9ԯ6��=�8�Ỷ��������::�V��D�{1�GD1�MH��m	�?ѭ���F��899!3399��A̽�y� ի��=��|
���e�O?�#"�rk�n���-����Us���|�^[����j����'~�0�\I�[���G����k胧����6aV�		���W�{��E����!�'���Q��/_÷����h��΅�ի县�m�Z,e��5�9����o�����JZ��3#G��"�Z���N˺> "˫[�.Ο?�����������z}��q�ٟ/����¢�dy��ʱ��DDDDDDDDDz���(����f���8�a��Q=�����Ø�7֢!��qy1�{Ktkd�f��
C}��0>U�}5��񄾰�I�F�Zj[�ǠΘcؖb���%�Ix/<ٽ&����u}�|�uL�a9��l���K�oǩ������]g.����T�:�e�CD��[ح0ԧ�=��P��}DTa?��[RDDDDDDDDD�&�o��Y��O�T-t���^/��wTbs��b�㸚�e��Ժ�/&�Ǹ�!��
=�f�����hd����tR+$㞟��R]N~?�����q8�t�*����C#�.�ѥa �"#'��[f�Ζ�������X���G�!9=��{�V��/3�-~Dd~;O_�c][��Ύ�Y�^�nZ��
������##��>�b������������H�g�`�7����qj4�H�[�`uy{T/�p	���æ�x�9��,��j8;�g�z��O.n�#i4��"��A����n�䩱����ٮ_��A]�^M��cg�xl=qiY�}���ℾ��1�y#o��-=�0��3V���˨Lv��X�O&􃇫s��7o����5�Tä�>���Z�D��%�ջ�.�,���eɡ8���o�����z Dd]��Y*�W��ϗ�>�c������������H'��k���q�t����UC�z~���>�T�/&������m�������*�T^�����k���W�}���V��g1�W0���HH�܇eYy��Ӝ�����	z%��Ý�����.]þ�$�=��#�U���bmn�%���>��W��A�h���m)��&��^�UѧQ-=|�N^��f����Cg�ĜQ����K��Ķa%~F��y���s����GADT^�*#֧v�Pa�Ԭlu����]*P>񻥆���w���n��WT��T"[f����C}���|���ȅ�����|j,jUw�^�8ث�r)NBZ���|H�������� �p)((����j�����]UK���ʲ��yL�~��MswK�D%���^z'�ma~��er����R�e{����kY��)9��Ӱ-y�����2B�~m�=Z�0Է�@*3y�~�sg@oD��w��
I���Q=Uk�Eg�H�$�'�{��Z���<J�3��6���Uͨ=?���-�ී�=���������Mr^��9s���?���,v��ܸa�sK?_��l�}DDDDDDDDDDD:�xE��,xl��[׌��V��5ԥ�Z|�����"�W2δ��s1��������>��$���/k1o�1TU�څ�����cZ�����@DT�]<�W�����2]ߛ�������D��3���T��ڡ�B�|���������������th����W5�R���n��[�7V�R̈́z'c~2?O����!'?���N5DUe��k���W����;D��<L�h����AD�C�nqqq���fT���3rr�����8~�x�y�T6������������tj��K��|,||=�A�s#;W5�I[�-�q�c�^��F��C����+��z���rl9qUݕYfY��Hڂz{��^�Z�٠��4v�BHH��ǳ��T�8�Ϳ9��|�l��Xܥk���\�����)�1��8p�l�4��i��:s��WG~<d�i70��%8|�2X}
]�\.��+��R_{�:㙞m04�!j�pA��4̊���{����DT�I����u�(�����s�E�	}�.�F&��,��r#""""""""""�9	�X޹��@�z~ �Y}O�Y�������X�&^��ӆ �6G�Z���$�'�2���Ø�.��F����^��:5k`�Sc��۳h�\'#5G4���!7� DT�5����ڠ]��j���O�Ǜ��Ѕ[a鵱g1�u�ɟ����V��VJˏ�T*�ޮ��k�����#�$�9HV^>��g{x�pUܔt=��9�%�ـ��L�t>��S;4i++7/-ۆovR�a���z~8G5��l���9Q1���Mj�3�N���_.������^!	|�y?^_�K}����%B}�Ɵ����k���*�1�B�Ť�p��}|d/�j�D����?�7V�� �1������xs��Jҧ�a�a�� k�ȳ����\�<�7o�;5C�� �pv,�^nc�`�a�f�a�7Q�$��?�$���������0�{+ti�b��^MÂq�h�^��@�+�}DDDDDDDDDDD6BZ6����N]��c{Å#U5�t��X��	ɨ��eda�O+0�e��,ct!�	���x~�ud��'}�Lt��/�� {�$�oy{�wHP���H�xgݞJ�%��I��gK��
9�����!2>��S0��_���h�S�h9K��M{Ad|�\�Θ^�]ݥ��R�;9⻩�0�i�˥��Y���<ֵ�z�-l�$�#�/����
]+Ǿ �F�dB?�-���+��N5G?h�7�.ù���_�DDDDDDDDDDD6F��_����@Ow�yH�苭��ʝUbT٢�Ǳ�\��4 ���GB���q����v�J���.��W�?��^�5\q9=S}/c�$��<�ن�x���w��?"�@��MK����N������K���L��&�ബll9qWnd��^I�T�-�G:�=�d����|�x�O熸x����Z�ۓq��ۄ��I�����G��;3��?���Q%C}�Q�ڭ��цsA!�ˏ�Ī��H��EC/�~/m�uj��/����O�#6�
��>"""""""""""�7>I�T�6S�T~xn��*�\"���|� wn��br�!�����j�A����U"��̜�����y��A~�1m(�=܊�˨��.���V��@"җn��bh��*�t��4wo,N&�-o�_v��i������<�.D��W�څ�v/i�l����א��E�����aB��r�\��:jo�mƗ�ޱ�g[`��T�IS��/-�"�l�d��Ⱦ #������R����|�e?�����<\�������|��}DD��͛7�������#������.�$�NDDDDDDDD6OB*�[�ک�ӫd���5����}*�Uܼ�ov���'�úab�0P����¡�%��9�j���up#;W���?:R�ݮK�@�p:��w4�ɸ��>�j?8~�����'�u��<�(�Q�/}�ᥥ�������߂��)�:D!�0�Y#uNԫI���㯦iv�0zlo��Ƹx̎�)w��_X���#�&�	i%�璭�v� �}��1�Gz#����ۊM��aVdt����{�.�Z��o�	it~|�D�m�:��  �C��~�G�U2���HOO/
���333U����M����������r����H�ޘ�%�:�4	�̉��k�v�bj:H�����`��cxmxw����M�g��ޅ/�TMQd>׳r��H�&i��q�o���3=Z��p_���X{V}/#�1���ֲ(8����6D�M{9���ԯ]���������\��ԫû����ycD�޷��)l>~ckm2E�!�Wvժ�C��
�I���P�^�M5��y��oP�B��ϽF���ϗ��O����)�pK��� ���}!��R���hSϯ���v6�nzv��uD��q�C�#""�IS��P_q����5��HDDDDDDDD�������r���֨��s�2N�=�Y��	W@wZg��l�;�)���;���NRYx0ΰ-mǹk�A��`c�\���^mT�Pjf���w������˼-�)����n��;�����튺�����MFoC>�}�G4�F~A����w����3	w�+��'����#���S�Ğ�W�Ʃb�FI[���u��VM��Ĵ*������edݱ~���>�#6m g5�tƞ�jĜ��AU�B���޸�zlr���s�b�>W��ȘƖu} ���O_�;�"��8����Ǻ�������O-�a��cg��5�q,���9;�f�q�CQ���
Kk�4�^622Y~����������T��7n�2:��e��:~u7��Ύ��M���fD5��?�i�ֿ��'��Q�9�N��;5ã��+#:�s�UP�ջTs��\�G�m��&T�fҶ+B���Ʒ�����f��k�Z���?���U�)o^�Km}B��券KWU����U��v=����}ۣ}�?/�E���{���s�ܮ)�wo��'���r�<�4�N�_�c}iYZ<}4Z��+q��;���8�r�X���G�4�)r�/蠂}�:?e؏���+ۗ�9�-	�ʨ]9��)���?��c�a8.��!B}��ʝ8k��+�K���qӮ��mŗK��HO����ׯ�څ3������=�p��j8o�s���2��d8����v0�GDT���݂r�E���d]Q�"!�51g�l��x�W��[d4٫+w�P�N��~�}D�I���
��l�BGt�j�>��ʝ8|�2H[��++v���G10<>����ˏ�*vsv�/�o}4:$�Q��um��DQ�%�eX70,$Ḿ��UP�9k1w߱�f=4\�9,$���֡��� ��\�Z�
IXm����[��:	�N��J�}2O��
�����cT���~yhW�
	o� '�����ľ��z\�o㋉��.������s}q@Gu)N��|��ܼ�y�Ѣ��C��ƈ���swqRAs	̍3<i�-�{X��XD�{]'a6	���?��)��e%(���0X�^��I�m�K�b���iCKl��xB_t��g�/���&MYų0��عA ��d��WH�������.��:g;�6���X�c���J���k��u�Pe!o��x�c�z]:�D�3�vM�2<׀b-Zr�_��W��!�-P�B�z�}d�
� �;�{�т��\]"��P�f�ݷx��c��a[�l�!�����Q?S�\���k$��i?�T��B.������x�
��뫞W�wg� Q۠:%���H8S������4mH�&&!�A��c�N����:Ȱ�J;_��`N6&˰���>�9��ٷ��.��G���㋼�|�� *JF�j�S�rl(���E������"�ܣPZfv��_-v)�a�%�?��>"�J$77�%�2�GDDDDDDDT9IS�4<}���л�j�*O�2�<�4)I0C>����mI���K�d$�P�Ƕ�>���t�5���$���6�a���U��4�.�j36��vcZ5)�P[�P_qP����*4\��&��⡾����)���E��գD��8	��;��
0		�|=y`�P_q��U��ﭿҒ�?�ؿD��8	ԭ?_Ғ��4�#��w��2<�s�QJH{]�P_ql�z� �}�g��+�+N����������8���B�a�72U@AD��[��ۮ����j���Vm�[Q8A6�Gd�
a$��=���ⅻ�.�$w�K�z��=���w�[��������?L�����y��z�ð�۽�	�i�L��A]��w�~���<��	��������Q�+���9�e�ᓕ�fچ�liP�9�}�x�����C3�����0��/3�YR9ӝ~���N�5Q~�l��[:lC}�n�OV'��k�.U�Ӫ��w��j^��1޼6����_mC}����c��˕�?[ƅ��Iuia*�ixЯ�P��u9��7�o˴��d��=WZUQ+̖W�7�ӽ��̧�Gd��_�sYO�Y�;�T�,�	{�C3ǛJc��౶��+}�g�r�����p�~?�{��rZ����kHQ[���W��̞_m�_R�m����+'�U=ii@��}  �*+s����,     ��I�<��&S���3�ɼ�}�;��޳t�!yf�.9�$�F�i8���{�Q���)�Mʖ@�ku8}���S��W=�1���uZJ�ʕw��˝\h/ݩJ�J+��D�UF�����riyYi��u�O�p�~>�d��^�қ���0[m��]������cW�����`���j�䨡9m[��XUm�5.:�T6�p�Q	��N-�SMtY�i�K�΂qV����}a^Z��Mh�E�bpe���1kl[�!�����Cl4��\�=�=���]dYM4D�A���v�ڎ�&�� �|�Y�㴂_m���7�2ا�Ě��e����s�`��K��c��*W�Z�Q�}	�Ι�}M�����6���j+m����τ��1!f���؅,Y��
���:� ����;$Ѧ�^]he��^Z!o�3�|.�z�lN�*�'3r�k��5�,�g��������a�p�1�w��G��O��)R�-��	����n�Z�[U��!2T|�> hFZY~Upf      �8z!S���������Ć����4e�X�#Q^�v@.��K�$��I[+j�.�hU��&��Xް����e�÷iu�����T���Ҋbw��@�Rk8�ku&3��o��F[�*��^m][^�}�j��е>']����k#��uj O�YW{�v�/;c�\{m.-n�}��?�����c�	���`�ڸ��//�+���պ|lX�Ӫ�U���.W�W����i��,���}��c�j]�o��-��˕�HmC/�{�{�Ξ$�u��TC��g��=M0���N[?gɲ=�ek�S�ӛ����~<�zG�ַ��9���Mx���}��dKOV�}�oH�k�4&�-,�^�-����R�r�M(ܺ?�'!8ۮ�3�jX?��@� �?˗^i�k����
      hi���
KO��!�G��oM�R�_������	��O���9uN~�t�i���>��4�GgsP����_k�Nʲ���e�t�=���L�1�~��mťe�m�?�ز��@��?�,!�n^va��&�����9Eŵ����Z��om�
������������c�}�<�̂���ٖ�S[E@�c�.��su�h��ܯ�c��ۮ�.���U,�jɻY{NQ��2WSE@��]y�:���0n�\�2n��RC����=iSM�G�6�y�mhU�ްG^�~@��Җ�Z)s��x�v��.�u�V�|��]���\	�ۏ��6-���|���M��z�F�U}��p�#��N��]����s��j��ۃSG��N���,iض����������L#k�R�o[������+�V�z�� hF\��f�      ���5�N~�Vzs��1-���/O���7�#N_j�ơ���l��L����f<M�ݥI�~.)+���O� ��
�t1dߤ���}������1�~�s�:��M	�3��<miX[�T]��rM-g����#'�e��jj��
mI�.��x�	R�T�NەZ?WL��_;��Ǿ����3�ty��O�=㝷m����R�����Ԉ��.�!L��W[�S�gLT!���ױ��>�gM����gU�kM!O�����5�O��[[�j�r���2��q��$�[����2�6�,��t|��_
Uj�M�������Ǯ�[��֤��ʬ5/�jCC��t�q�g���������,�ߴ/n*�2��&��Jۙ��_n3�������u��Z��9٥1i�O�}�y��Ӷ�^���~r��&���?/l�k���g���G|Ui�G�(y��)ru�nr�KV����0��-�x�sYKlMnض��{�g�~W���ߙ/�n�c���{G+��c�t�+�﷞�Q�Ueg_C� ����`)))�5ܧ���     @�;s�L�t�9 ������A�b}��%4Т=7?#��2m��{4��Җ}fҪ�{v6��i@�Ɣ���g/�j=�����3�-���{_�T�ϔ&�l!���/�o���]�6�ۼ״l�jP���w�.����3uF|����Z��M��W�o�%��uX�M���[_��`�Wn��gMp��ܢby��/*�֐�ۻ9jhP+�Yi���㇘�G4Pf��m����6�q����#)�ٕ?�b��w��N�����ZX�Hi%��Y��_o����Ӫ�VZ�����M�őӖ�^���;ɴ�ӽ���X�s���p��_����#/n�k��R��
�-�#z�5��!�_��(�9i��?���ʿ�[�7�R����������/� �@�~�9�jE�7w$V��ہ�1��&���olO4aD+}��y��n<zZ����<}�zt���m��硆v4ȭ��t{��/�-x���~6�~^ח�o=5�Y�ż���w���t�e4����y��Lx[���f�x���F���g���$�߹a[�P�W��ߘk*q��˃SG��*��J���_
����=� ��	���\��>��&      @UZ1���m�'ˤ�=Fu� c{t���:��C��`�?�r�|�:�!I�igJ�l?�fR�i�k �I��p��N�2�s;S-r@�s0ϓ4ȣcI+�lIN�/�������NE��d��u�6�Ӿ�	������[.�]4C&�����a;C�x���5t5����E3�Z<j��o�o7a8[������򷛮����9��l�Z���q��Z�C4��k��U�;z!S��39b�����WI^Q��u� ��V����ڵ]�j�7>��<{�2���6��t�!yp��*�g�reγ���f�*TV�y��58nK��i�(�t��|�B+������U�-��к����	����� X�����Տ�Yky�JM`�6L�G}��6A^}�������rݠ^v�Ѱ�w�ZeתR?;�s�}��ko���7&؅�����?.�r@N×�|��ih뭝M0�9�M2+m9��%�W�d��6���ߞ2®B���r�mj}�n{i��c�4�:ݖV|`�g&<h�}���m�����C���!C���7X����Ig��V�[�����gx�~��>�b�|�;�s�j�u�z�5泹�~}���ϻ���Z��J��߲l�	�����4L�Y������n�ݲ-�c�}����X�w�H��U�����	���ǷU�?��+��` 43�,?�5�W\\\Y�O����IPP�	�      ��),6�IuR��e����6m�4|�)2���������V���4�v�d)+/7�TZ��Bn��e��ٜ<�8��+�ϥK��l��4m��ku<��4����m"MU��1��%:B�C�$"(Ќ'�DZƗ�����2�b^�	ꜷ��t�e�jEG�h�/�&�T��O�r���f���FVC]�|�	�9�-g���k2�WgS�O�kZ1鼓`�V3�V�W��f�.��g���)tkH�o�w�+��˕}��mF�|\�gYiXO�?�f�L�'��~�y�<�氕�V{���weh\;ѥ��\ޚ|�Z`��@�E���7䊞�M�W�iu8ga*�e�c�"],۾ޟ~�8�^�ݘ o�:$W��*mÂ�w�VH,*�������]gB��z�IH���?sQ���:|�Z���W�P�5`�=%ͮ�-}�~�-x�J?ť���ipD��O�b���g�~��<g��4h��th{s0�?|�ݰ-}_4L���d�s��,�{[r�	�U���=�~l*J�����4|�l�j��<��y]4�]PR&�,��>&G4<=�/�D������"Y��b�<M�Oj5�O-�3�>�f�W�Kao�D5$�L�MUS�|�����~��}�?��i�y\�Ε��X����=&�ix?sr�V�Ԫ������2�����\�&�l��m��Ͷ`K���Ă�?�"}۵1�7-�>��`Z����j~�:\�Ĭ�u���E� �����!>�       w�.^�i�������l3M��tr���Zk�Ք>�%�aKCb�T�pWm��R��M��U���$�`�N�������.?�i��Uz�^+v�J���N�|U�s��yU+�9��U]���
�U���DC�u	�$}U�����sur�~�۞ x���̤�1"����|��=i&:ĵc�z"�u٪�mm�n�֧۫�4S��d��S��P�m��mZ�	g�yZ���������_D� �'��f_yպU��۴          мi�:��z��>x�s��)�7���4��dw�,ޙh*�6���\
)k�P������54]V��mUW=T���k�V��O�r��l�Ʊϲ-�s[�+ml���D�U�  .K/iؗ�g��c         �n�Φ��Wʃ﬑�{��W6-�m�t�
��_5�L-�k���u�`�.�-��Sm���M��w)̴/��������j���:&�RXO[��ԎW��N�����Yתw���pU߮���7���k���J�:���\�mHC���`            �,m���=������#��mcJ�6v��#?�v��욱��D�	�9�Z{u_���W&&�ͣ��5�
�
;������w�XtTZ�l�	�Z�7�������ȺCBB���@|E���l۶��'��[�o�4g�^:-�yK�)}��+wΪ����V�lL�            �,9�)O|�U��j�L����f�i��Y�n�J����L%e�Ҕ=�z��8��y~�:����/��-�MR�	,���]:ȷ�7����d��?���\���6��dggIVV�������|=��o���2�p�Q���bn�i��36Jf�%��Q��`�;|�Z�"���*--?��7          @�PV^!�&&��mX�,�_n3Pw��[N�oV�������Ȓ݇�Uo}h{�ﾵJ��y�	���V^�s�����L������������4�W\��Jj��QҪU+��̔���竚s�oh\;39SQ!�▽���k�e_F�@����/'N�8֦M�z�          @Sw1�@�ݰ�L|�e� ��[.<(P~}�x3i���;��=Ir6'_|�ۻɾ��icd����U��j�o��3��}��BnV�&����8�>o?__	3z}G%:4X:D�V����\6=m�yn������h������222̿��          4'�.�#n��?�bBp������u3�ym���L�͙$k�N�;eٞ$�<Fm�����6R/��_�Ą�v���m"$28H�KL�����%#�P|��CnV�c���5���0���p���'�-<��f3u��1��9:²m���ʓD˶��[� �(��\��>M�GDD          ��\����K~q�˷-*-3A=�:G�ˢ1�ht�􊍶[οuk�>���k��k�������N�5SS�X!7+o����6v�BOJ��3�H�4e� ����.==��K�         ��y`�yx�s��=I��>��z�d��_Vm7�V�����`D	
xGNN������o��;�g�X�
��} Z���B}�D�         @K���9���������́=M���>]��+�>+�igfO����P��>�E�@��_R*���Ϗ�����ʖ���~          Z�Ry7ᰙ����k�{
���B}Vڦ�|��Z�}�-�4 4{��pAC�ޮ          xޑ�i���4��!7��� ���ןopp�TTT|�>             ^��Bd��PG�              �!�              �!�              �!�              �!�            Фu���y��zl���%�Yb� ���           @�6�G'3yJJz�M|I �[�             �C�          �Z����� �-*����8���$-;OJ��]�]�_k�mä��\���KyE�  ��        ���'􊳛��_(k���H[�u�
�����9I��%  ��� �ah�&��L��E:X����d��ۻɓ�wHVA��۷�%��P����=Q�ߔP�2#����ʼa}�mX��WV^!G�gȺ#'寫��ٜ|��}d�D�gy.��b�}��v��>�b��h��&�ʿ7�����K ��`        �i�;��Kw\g7/��9�����}�ʑ2gHo�y?\�Z^"� �1��&ӽ�ݼ��	
��Q��ëGɂ�dγ��؅�j�����]��z?k�Rj��ʾ]�;gITH��[��KxP���c�e�����o#g�	j��Cg�M��{L�|k�p�ڿ��xf�	��i;��#�& h.�       ���͟o���u��{_   o
�o-�E�|���-��Hai���w����FI\t�	�]�ԛ���3?zg��;	�%�Kwz��q���{�7-�5���Ǜe�ᓦo��`�9Vn�Wr��WS�o�Z^��z�;|>C�o��W]�a��f���S��]�|$  ��}        ��[F�˼a}^׷}�}  ��\�SVL6U�lie��}􅔖��Ϯ+�;�ʔ>]k���Ɂ�}o]h0�_7_cB}�N���g�KaIi��Zeo��Sfrd���&����}���P�Z{��������i2wHة�H�(  �
�}        ����tzݠN�2�s;�{�   xKmmM��y�	��aq�jm�[W��2�A��e��B}����~��M�N�jU����������M��Ɂ�� �� �       @#ӽ��S�2��(?w�   ����RZ^n*����v����7�~y���`^M�Z��ɽ���Շ���dӱ�r���rU����'�  ��`        ����k]��������L   |��nM�O9�Y�����m"$:$ȴ�ݙrV>I<^�ͯU�V"W��l.�HI3�j�y��H�p�.,��#MV�;&�����=&J�.E"��e�3�Φ�`_��5�d ���       ����o��q��UkK<��;^�P  h��H�oVA��>t��e�0wr�y�����֛��Uu�7!@u�b�����rۘ�'C��9�r�����'���U���9��麈�@s5- �7�       ��0��9�l+-;Ov�<+��������  _0D?�=������[L=g����Sg%%=��=�s�9a!&4X���Z		𗗶쳻���`u��a�%:�T�{m�~��u|s�0�*o�;Wf<�Dv��ܮWO���,(t����*/�� ��}        4�;��}{�!�|�L�`���%.:BNg�  @c߳�<�p������ݘ�p9m�;�W�؅�mz{�����1W��o#O̻RV<a��p9Π������?���
3OOvX�;IV}o����s���.��M��_���R����:�� ����r�U�Z�2�;��狆!�       @#���{�U����M7��
�U�V�����o�w  @c�P��{o�� ���۫�.[XR�0ԧ�/f����~�H�����O|���������"�Y��2�g��vQ�^�K~~�8�����ɌK����˷����l+�v�*��6h��~���y��\\滁)8(���RT䛕2���$,,�m�k
�744�p�!�       @#��U��h������wv�oOaw�m��<�f�9�  �M�P�V��t�����GRҀ0��Ȱ��Y۽�	���*����lN��,�Ⱥ�'M�O�k_�˲i,�ض����0|Sai���t�����ӧ}.�VVV&��yn�)_}�����3�>��}        4�֭d���j��<Xy���Ղ}�c�e\�β����Dp�����n�V�ْ�Zm�+zt�Y�{˘��O�6,�����˾3d��t��aX_��^��iy�r1�P�^Ȕ�����c��D�����YZ֠�O+�����n^~q�ˏ{P�Xib7�йI��u��W��*Ukh|q������6J��'S�t��b$�r��z_�-0�GNɧ�ɲ��)�Eۆ��ܡ�eB�8�f1��w��P�}}���
$%#G�[^����`�E ��+lB}��w��>0�u:����]���-�^�/.��� ��<��Oɸܾ7ڦ��q�J�U�m�mإ�Ҳ����>_�YC}��k����!�       @#�ֿ�t����PZ^n��Yi�>��74���r����`��޽�F�y�o��/W����Ξ(ë��.i%��\�^1�[Gyb��oU�^XCn:i��W�2�{~�l���������<Sҳe�^��:vl[m�Zqhܟ_s��ZUhΐ�v�~�t���e�K�_��y&j��o�k��J�7���`�j����12�L����w�i�xo��>yN�A� �s\0����9\F�N��rF|yh�x�jy�l��NJ �oխ�,��\�����yOr��S�����>��~�
c��mu����Sd[�/_���}���c�=Io?���,=YM��x2�W�W�K+:�﫶�p?_	�y:�g���ԩSR\ܸ�B�-�A	��.�}        4����6o��s��;��n�W��u�W䙪2��[��7L�oN��u=0y�<:g�Y��Fv� �}o���5�����]ݯ��x�uv�j���O��@�y��p����c�������gy��'o�:$���c� P7|{��Lܽg��M�y�m-k��J�YꀃʭZ�U�}z2��ҵ�^U��^>q�@�}8oeb�,/3���~�E��j��q_� ^y0Y��L��E�5�+��'�����y+�gեK�F�]
��V5��`        ^�-J�Գ�|�6�VKw�G��$~��q��ahyc{��[�V"���Y8���u��a& X���iRTZ&竄ᘆ^�{v�B�VZY�;���}O�>Y��d�D��գ��t�iU�y�/7m� �g���x�}�L /1�������_�����S�+���՟o�ʴ�U����̛;�g׌5��Lc*���}��^��I8}N��ϴ�^��j�O+�j����ؿ�(	��3a�W��]���v�Ϫ��}����}        x�B-J���G��U[V�MZAf֠^v��'�}L�0�w ��$��hZڅH\t�9H������tx]qY��:xB�9%�Y�&i%m��-��!F�}�4yx�FA�4���lC}�%����i���93�Z�n%q��yr�.�mm������2�/�׹���Pv�++��uGN����~XW��ѵ�\?��� U�i���d�3K��  4���\_����,�:ݙ]'�V����ݳ%��D��:d*��HdH��le�7u�5�-ۓ$_;]m��
�7�߾v��;a�����^F~��,V~ey<�,�m%e���w�W����&���%�/�a���IJ1�y����oOa������}��nS�X�>+o���5�        �2mWZջ	���^ߞX-�7�g�􊍖c2�]ڄ�C3������\^�b�<�n����qxm�[�����MW�`^U�8.?\��a+�o�cn�a��=�<����Wj����%$��a�>�z�<�1A����p�Ӗ׹G�(��]�D�w��?����}O�'���q<����%�ˉ�l���(`�y5X���~��ko���x 4�h˾�U�}����Ԁ1����D�-[��zm}�>"T~:}�ه����������8����^%Q!Ar̀��{���~�<�f��i�p�Q:�g�U�o��;�g�Ҟ/\C�        /� ��N�+�i�9gV&&�*2�n�JCs�F��c�lv�cӃ�V�E2�?�Ɏ��o��y��Ӽ+��e���>�����n~�}�����+GT{\pL+��Y����%�˨q�GNɬ�#����TK�uۘ���Uۥ�����ՊGO͟Z-���ۘ ?o�Դc�z�FSQ�;fU[�]����^ �'>�jB��8��gγ�et��%�V���z�-;1�r�e��s�Ξ$9�vѥ�����r�؁�R�V{�j��{y���
���w��ޓ9C��M��J��().-�#�3���VFӥ�<�����Ұ[RR����{d����RT�z{qO���

��b�8F��       ��44U�V3ے�ʌ�ֵKv'ɷ&���hL�<����ԝ�J�d�s�eϩsu���ԛ;�O���=j\�zh�S=�Ѻ�XNa�����.W�9��+�|��t�uv��D���d�q�c�j��ҷ]�j�������R������������7k��{W��;^�P  ���=��V���]��XN����u�7Q�}��M:hZ�������Yw�~�����deeɑ#�����狚�       �K��e��~��/�y�� ԛ������U}���N��a��8�	����\m�V���w׹�R��O�����u3UyP��?�T�Vtp8��#q_U��խ�K���&�6O[�{W^Q���󛾔[FǛ�N����T$<��#    �R�       �K��]���f���y���j������mL�[�}�������u[mշpd�j�_޲�T����9���{�g׌��|n����@�o�����&ڇF����-��/��G߻�<�G?�,�|�����[�q�Ǖ�   �	
�a�[Tl�_hz�       �%��Tm޶��E�+^�q@~?g�ݼY�{K��`��/t�cԐ��⭏�q����Iz<�j���
���%�:_m^�6���n\�N��iP�!��N���<�f7|�8  h.�r�U2�[G��׊ڟ8^�rZ!��W��[F�K�vѕ�s
���}G�5;���t|�'�� ��2�C[k~���V.U���~�d�4�        ���1�2�w�j��LtyKv��Ξh*�Yi�<m���M_��q�;|�޷���Ui%��'��Σ2%1��wl+pnkr�ms�IN�޾7ʅ��c�W? �AUG��+��}�����յ��nժ��}  |Q��h�*$[��u�m�䭯ϑ�b�]aٷ�et���O\�Z����o��ܽ-�~�l�&����9�>��D��}        x�mcJ�V��2��=�]^���Zu���سں���}�l�o;�A������Y��S�������z�V+�T��bU#�Vrj��r�=ݯ}*�   �څ�H\tD��g�r����Ε#�U��ɿ��_��A<EO���b�ż��ת�oc��_Rzr��6�$˾Sth�|mx?��+Μ���i�B�|�;��>��8�5E�        �0�4�hL|���B(���N���U�}Z�`P�X�k��29�� �+:G�U�� ������e��m�*,)�6/ȿ��a"B�����1h�q��::D��  ����dr�Kձ��e�_^wۺ�4L^�~@�zf���WH��,i�M]�;nY���cV/|�W�5A�,�տ����2�O����W,�l��-������������*�Z��)"�       ��]շ�t�� bU�X��/�6��v�o;P~��zi��bi�(U�2j�����_Gs�_���R�UƠ���ꂓ1�BA  ��L�ӥ2ԧ~�|����q��5����&t�tIÇV?X�]���я7˕��%ZuY���G/m�'@sr�S���ʉKm�ni*�       �a��J�j�:Q�uik��������_0��<�bS��n�50�(ؗ����V�h\��*$��a�l7�W�N�XF�4�r  �s�5yx��g���]�m�e���
aC�ڙ��3�{J��pIu�kl�t��/���돜r�\yE�<�a�<�h��[���CsS�ySF�  �h~�$6$���)+�p��e�����2)*s��~f|��6>�K�   ���� ���6?-;O�3eD��Pm^lx���C>�{Tꫢ�a�+4�UUIi�4-�|O��V�%nx�4��+� @ˢ����^��?����5w��:����͔�#��_�Vr��x����k��Qy���k\���ds�AÊzřs���T���  -��vQ���1RRRb&G���%;;[�w�|z2S od��vq|�7�<��   |��#�;$�k&w�m���J������ (�-y�ߣz����*2��:2
  �ֵ�=*������In]�3�v�`��ڿ�G�}R,)/����U�رm��)i5.�!��s2�C�ُ���v��3����c[h��       �A�9h��)چ�cd�����W�pT]��"�}+����ZZ:-��V������:�&  �٭c���I)n�����99��+���ex��`�,)kxEj[O/�&��u�Я��KJeGJ���wL^ݶ��pS�V"}�EW��\C[a���&ا�;����G���`        2,�����k��ߺ��<j��}�Ni��W]�D4x��c"�}�r�]̫fk�����Z4佺��(��  `kx��}�5I)��#�3M�/$�_������ܺ��}���l��I���������?�UO8�mX``eJi�6�6�t��WԶ-|۲-�t�-4W�        ����{�>�l�`_b�E�گ�ݼ���JCn@8R[�V��*���n���[϶�!<wY�8hQ���   lu�
��|2#�#�q.'��r{�~��T��[�o��ϐS�9�_\*��CeB����}�v�!�����m/��O�v��@��OAIi���_|��YxPëk��Ҷ�����E��BsE�        ���#�W���D�y�c��ǜ!}������k�F���$[��x��E;O��6���Z5��X�C۝i;���vp��A�dy�J�תmL�N�'ReF|�y�^i���������[Ց��_(   ��C�*/��jr޲���U���-�	˹�r���I��sx₶םk����׮��a!�׺�<w�2����؜�RV^�R��B�}`��4�ڶ���������i�����\�       �f�����[����貄$��)v�V�k�`_JZ�y�~~r�����yׇV �i��,�k]^QaY��Ѿ��Ⱦ3uo��A�+�v�l?Q��փ�W��Z�Yzp~ڀ���+9M   �

�{q���/�˾������~��o?��:�T�ޗGL���[`���,�H�M*\��n�b������>����$�u���Ee�;�p�ڶ��Ͷ�!����r[��0yⳭ��       �n;��<m��b�Q��G^Q�|������n���������r��ْp���ko7������g��=&�ʧE����	=���?�?�x����ܢbSі�g���f�n4Z���	  @Uy��x�O��Yoz�����O� �nL�Mm��9�W�`�m[]�U�k�l�̭gUm���^�o�#?�6��=s`O�}        �~���pX�����Lʝ��>T-ا�oo�G�<(������כ�}S�t���˪:���5ԃ6�aê������������+��A�e{˝��͟5��y��9U������N[m���˶s\   �J�/��u���}t����L/���je�`_|��ծ�-*1�
�����."TRҳk\g�p��big����/�V��;����`  �(���td���Z~X�z�J�+.����7�oʒ�9+Mn�_QQ.��[�{%�sϥJ���^{��n
s���>;>�7���g�3�   hY��m�W�%���~_�:!�
�U(ъ���[��<2k�	�z�kSe�3K�LV�K����,��Ǵ��IY0��ݼ��:�ʆ����`�o���>S�#��c�N3��Zۏ��|����R9����z�J߳�^kZ�V��{]n�  Z��92�S��<�w�����@�@��L��e��;����V���|1[���6w����ݟM:�.@S`�-heJ����|�>  �1�E�20q��W�KNN�T8&5��Lז�j�5�����WB��"��D��������_լ�筌O   ��[4:�����B����IkRRV.�&�oL�oY;�W��6J�/f�7e�c�l�?λ�n�V1\~�<���%�\F����!F^�k���;���'��	�����ir.7_6=]��� �o�!W��,��m���)A�5y��|}�>�֍���#�F�&mB��7O�kt�v��nc�*+ ��C+[+<k�h=Y���}'��:�'��~��'-�K����(t�fW�y�`�иv��1���Z�o�MPQ[�M��Z��m���&�O�>s***ڈ�+]�rlA��n_oI�nR* ��������P_s(������$	]L����ӗC}́��|�p   Z��}�H���j�5\�΃����>T-ا�5`��O����gӗ�`dSϖ���h��{�nyk�A9x־BȀ�m�Q���M+�J8��З����;��	C��k����I^۾_�؞(;RҤ��������d��^r��A�B����4Lp��>�l�&Wm��+6Z���ya�^y���jKd[Z�qް��ëGI�����_+�|����_\"   �hef���ar�A��/�t˺u��W_�>l8zJ�M�G�R�r+�Um�k0kP/s�J�o�g7�q����;V�쒘v��j�@c��򶐖��b*z�kB***~o�g��8��t�����כ5�k� �� ��}��\G����  �����h��S�&�1�ͪV��ut�<��VS������}�S���_�NQ�v�i@�����t!�@����"C��V[�S��Ɇ�ԣo���6|miٻ�6��L��1V��g��5;��	����ݭ/�p�~���oY^+�2�$-+WJ�˥]x�	�9jY��������� ���@��u���������I!��P���I�ep��ʿ����6������]5���6!F[�?&��0��WM����j�ɑ;l~���pX���ڶ�tRZ
�}  ���B��u��*:t���	���0	�CBB���XJJJ��yyyRPP`��N��Ȑr:�p_�B����S���6��I�   �XtH��ܻ�|mٵ���ݯ��^���	��Ҡߔ>]��$mU6��e�⁯U�Yņ��ə��3䎗VȐ���x�
��o|*��c��ɖf�bB�����M	��G����J����^&o�s����n:զ��L~�t�,ޑ(   5����?�"K����'��}�\��w�T����[�3���MGO���.��Kv��U���V��ǂ�����<�*�#z�������L �O󮔻^�H��߳��2*�\�}cg��5mڴ����{d�aa�RXX(�ē�744D����W趰˲-��a[��nO/�f�L+�-|� -�>  �6����;J�޽�K�.fҰTll�DEEI+'g��D������ٳg�ܹs���&�N���'O���~�s��B}���ϟ���T3>uJII��I�   ����%8���z_�;��U�8�)m#��>u�|�\����E3䊞uí<xB��SI�w�o��v���ȫw͖.��Ry��M�/�;v!S���m�ͬ����CĿu�:�ckr�<��j9�zQ   \����%&˵�=��}۵�M?^$�|�,�uH���\^W�p��+�p�����;���a}��;�������ӓْ]Xl�lx�i�{����ճ�ȞS眮�7����%*$H��#/�1K���I:�.A��wʣ�O2ժ��lv�~����F���)z�(++S|�r���1��deeY�s�+Z��<�X�n��:%=[r�JL኶_m�T���l�O:�4 ��El�i]y����S��]�.�ҽ/"������D8�RB �_�i��H||��~�ի�	I��h�J�I:����ʳf4,���/���&<u��q9v��߿�TO��S��B�����ٳ��k��+�S�C���   ���h�0D�x���vi�-��t�R/<(�T�������=Vg-�B+�\���2oh_����2�{'qv.Siy�9�������J:V}�G�������+r��ar����;6��9�Ų,!I��f�	�YeU{<�2\��?��D��K��u��뎜��¶����U��V{>������E���������}����uU��VUPRjƿ�u�i�  PW�����������p�����7�&��]�d�T�~�Y��[`�=��Oi5�>����.�ej�nr̀��7�_��^��Hs����3<�j����ŗ��7Ը����L���� ���^�t����Z��)T�����E�i~�df6n�OC}ڭ�Ӭ�%|%�X�m��_��nM��D��Wvz�V��z�����������IsR��4 ���X�>mYھ}{7n�<؄�����f�P[���q�c����*~����9t����+��K�S���   �w<���F�������e���疋7��m�S��Ps�cd�t�
3�A2�$�\��:yִ�J����j��g��2��ݭ�����))+�y���.�R�:��!ʆ<��4���wŝ�U��ǂ\փ�:i՜>��H����j._����~N��{Ϝ�<  ��x����孯ϑ�V��}��\9B�##*�������nk���&X�N��R��e�hP�Xs�#�o�'<<�n�l<zʥ��;|R&��M��SL�>(چ��^Ȕ?��fN�u�
�YEDD�+��P���-��L��ƴ�2f������ݻ-4'�  @�x;ԧa)�r6q�D9r�8д4�j����l�T���J۔)S��t��ٺu�	Qy
�)�����ܶm�<���O   ��:��/�&&��8��m&x��Hu  �$ݧ����M�ͅ#�;].���L5�O~�l�,����8�w$�I�L]�DJ���v�Mh�9�%5+O��9oNF�+�����椕!��I��0���Y�䔦�ۡ>+��aoW�k��y�r_cV*�Ķ��ޣ��HsA�  ԛ7C}!!!2t�P�:u�>\���|*$Uwi[`�g���ѣG��mǎ�z�j��Ӓ�S��5��g�m߾��	       h�K�7>���-L.F���Z�&�s�/��g7�1�>O�Jd�.d����yhe��F�K4F���R%;��+�g�Xaƪ<�-4u��d��]*�Om=�����Ew$�r�-۞�DDE5|}�Ŗmپ�F�U�,6Nд�y!ԧg��������eҤIҳg���iJ���4�ԡC�4,�!0�%&&�G}$���n������B�������P3>�z����Ǐ�����       �Q��s�7?��}�L��E&��,:����`i,A�~�UX$�y�r&+W��H�/����)gM�^x����:��V�<ߖ��C}V�3�nHG�ɨ(+�r�h�
ˇh�=X45�,�^EY��¥�^_y�e��I��|���y0ԧ�L;w�,�gϖ	&H۶m�}4尔#���6��X����HZZ�|�ᇒ����jI�)���P���?~��n�Ƨ�M�RSS�       �&AC{o�<h&�._	�Yi%;�p_cW&��p��"�  �ē�>�k����M�fE�10�Hxx�������p�=��˗/w[��%����Owb|^�JǧV�[�l�        ԛ������>w���k�T�B�  �̓�>��w�u�Ɍ3�M�6-&0U��=�ѣ�٩///�{��TH{��$%%���o��)Ƨ�9�Za��W_e|       �:р�/U��*00ȭ�ki�G�����EEEҜ��;n����gZ���� �C+T����)(��_�>�aq���wy*4�A��c��M7�$�{�6c�%����h}�����)((����g��~y�7L���h��)Ƨw1>       �;���.gB�kN�8!-ALL�	���� ���vQ���]�6x}yyy��hzz���h]\ �׸54�a�={�e	f���:���>{��y��x�	y���O>i�z�Sx���x�         �g�  5�����Ŀ��m����(���k�n���h�L��V��ܹ�	P�:uJfϞ-�G���{NΟ?_��6����9��?���;w���$�       �E��H��6�+�UXZ&[�� ��}  �)�ڿ�m�д
Z�^�L��'�ִ�����������{L�/_ޠ�hM9<��P�a���G}�E�O       ��}mx?yx���WJz���K �B�  8��P��Q�2e��r�-K[�z��VG���VG�;w���Ǜ�h��>�bx�ݡ>Ƨ{8�4�%[��         �`  ��ݡ����˼y�L�N�P���i߾}�ĉ'O<��������z��)������y��כ���e|6���Ԡ_K�         �;�  v445h�J�NB�C}�Z���={ʝw�)cǎ���2��H�޽���Ӓ��)���o���_��?��^�k
�K��U�_Q���q���o�!�V����	�       ��x��<��&��Wva� �7�  ���� 7�����ȑ#��_��t�֍Д�h8�K�.,���r뭷J�N�L��>�/���곎�{�G�w�������S[��|�ך��       x��if��`  0��������M��m۶R^^.���X	

����0a�i��OJIII����)w����g;>������⺟�H�         - �>  ��P_hh�L�6M��.S��!�B�DDD�ֲ��ɦJ�#�<"�=���y]��rg��:>��nHH�Ӌl�g\\�<�������^���뼮@�}         h�� �¹3�.�\s��q�&xCh��4�ֻwo9v옹�裏�o�[��֕/����ӟ��,T�����̔��]�u�        @3F� �̝����H�9s�,Z�H���M5"myګW/����7�)�ޗ��U�u5fx���<9����u^���y��Rq�O         h� �B��R��7�����4<��ю=Z��կ~%���u^Wc���9>����>���Ԫ�����        Uu��)}�H��hil�@�֒UX$�y�r6;O��H���礬��  |�>  Z w�����ԩS��;�4*��<����TFkժ�<������F


굮��?K��S��W_}��~��O��I�       ��{'���H�vm\�MNa��:tB�ߘ ��� hl��d�Aޢ�")..6 �(,,4Syyy��$V�۲��ǝ����`�<y�	���A����Ä��r�/�KS�������F������6����S�p       �\�G��?�x�Ą��v��r㰾f�`�Q����r1��'����C��A = O��.��4T�������O�URR"h�MiKӑ#G�Jh�!4廴j]�n��ĉ+>����/��{��p�e���$�       -�/g\!?�fl��3gHoѵ��}v�����' P�  h!��jݺ�:T��.���1�O����H�ر����ʀ��o�ŋ�k]��1>[����[n�7�|�^�"�       -�}�9��e�Ɇ��dǉ49��+YER\Z&ѡ�$C��ɸ�M��u�V���!��'W>��dZn �F� ����)իW/�?�t��U���MC�v�Lܴ�4�3g�����_|Q�u�3���`��g��S����������ܴiS��E�       Z���m��s'��������������1�l0a�d�h��]I����^iF�6;i�6MҤ	ً��3l���{/�:H��C�,Y�~�|��ҽ�}�Œ�:g���/��O��)�Uu������k��Vr�9����Ğ�뚜`��o) �k�  ݷ.���P����84���*��6����cǎ&�w����;�W=5������d۶m�z�'R1��F�G�3:,�V�����ק��>O�������O~��U~�Q�>?���       h�~7u����8��]�M�|�+))�py;�g�O��R>۲G^��|��7�_;<]��z��>��?O^�X,�Ԕ����3�  !�*�������d	2m�4BSJ��v��Uv��!����<`�~�]���7�>��S��9����4�����>�6��>��q�       ���qr~z7��g[�ʭo~&�}[l�w���b����KL�>�{��~�9��2�����= ��㏪�*%66��֧�W����?��aLL�>?B�  �D2�����}�{Ѽ�IC�N�d߾}&���P^x�	d�g�n�(�ݻ���'       �{n�OBCN���J������oh8�?�6ȏ�4���+�[&~�m-P鴩C��]�OC}���M�S�����.ܧ������ �  \ңG���K%99Y*++�-11QZ�j%���2v�XY�~�,^�XU����K.�>[����U�        �9�w��W�o4ᾦ�������g��`��X��.Y6�4=��S������C}�?�  @�4,5~�x:t(#N[�:HAA��ԭ��*7n���	4Z�:�wذa�g���O��>o��6ٴi�dgg        v:&��)��7Vnn�u�ΗŻ��^�����)���_�n�����E��  �
�~���ԩS���B�r��V�4�ٳ��4����K �ǐ��N}�@��ܽ{����ˏ�〫O       �w�Nm%������b�y�i,�{�)ؗ*o��"����:��܏W�`��g�  @��u�fBSqqq�8m����%))�tB4h��5JV�X!�"--��l����#y��9z�hY�|�        ��$'8ί;x����ή����\a���\�\��P_` �  ꔐ�`ƛ�^���\�#yu����륤�D���>�D}�\�۷7��#��>���       �������EM���_��������n�r����  ��X,ңG������J�r���Ijj�>|������
����'������믿.        $D��喔6��s�O7BH������n�ރ?��|�x	��}  �V�3f���V^^.h�Z�n-YYYr��q����/�����W���ر#���s�������u}       N�����UV���Ա�������^'�|O�n۷o��$���)+k�@hc��^;v��ǋ��  g		1�ЦL�� �۵k'{��'N��7�,�?���#�Ϟ={��ɓ�� H�	       �n��,ѵ���WVɎ���;,$�q޳�`�B-����噰�7���[��B�_��!����s�N����/F�  �A��;VbbbN���������1b�t��M���#��^�z_���(�	       �V���_,5sq�Y��d� �v�  @5���&03n�8�����m���ݻ͘�k��V}�Q�'ڭ��^ڵo׮]�>���:y�G       ��>ݼGn~}�����ңM�	��{���+MO���$!*B����x~��T�
�Stx��M����䕔�1��H�!`DGG�7����$<<\�}7[	[�՛WUU9.��ׯz�y] ���-**�nhA(..Μ�������HfR���;ʘ1c�� ����9h� ��O       @�>ٰӜ4dS\���vH�[Fh�u���o���dx�v�?��$��:Q���&S�w�!�R%>*��=y���1��j���r3!?����"�B媡}e�m�S���$.2��uN����%�e��#���!`���9�[�]���w�'c�W� �'f�W�?�!?�W �K��Ν;�ȑ#��ڴi#���)�_~����`��Q�FQ�A̹>g̘!�?��        ��B}�ܾ]�)h�B��ult��{���!���~xh����Μn7Pny}�l���4徠A�箚���u�1���s�z��ǋ�ʏ�*�0�C_���3����kdd�	i�O� |+55U�j�b����SBB�鈗��cBt:���ѣ�}�$%%E�B}9������'        ����	)m���v�K��X�yN~���l8t\���c�w��=;��}۵�9w̐�Ov���x�/�iPo���H�d�����"ӹ�k�x�ث��O�3����IEe��f�b�W� 4�:����v󋈈0'�i�O�,ҕ	�ëA.F�B��<xP���e�����K/5�]2cxG�M}<8�W�	       @c\��l�{"ףul?�-/-� 3Wo����3�?�[y��i�&.�t,{���r�����\g��x�/䗖���Α��IvQI�׉������'6�w�=D^Z����������v_�w`�N~��OC~�UC�=�5ޓ��(}��5]��ǟ#8%%%ɑ#G$++K�L�"���z�@��Q�p��p��a��O       @�q�GA w���4��>�/ێeI}o�/�sXnzm�̽c�Y�.~�S[�@ �R���cB}�*+嗟,�]�˰.m%�b���䟋׋?"��/i����"s�N~����E:�Rǜ�Ai�T��8q���رce����v�O8��lժ�dff�E}       ��ӂ=��5#˥�i3u�ޮ�Y�)U�!i��ͻM�OuH�E���� ��4�g��;�� ��hu�i�~�د�кuk�Ӯh�~���O�&99���>/���}        4�PN�#�!@���:���XA��+�} ���JJJ�)**��ЄRRRd��fvUU� J��z���7cp۶m+>��'jc�[�^�����ѣ       @ J�����*)(-��6��It�����0��/������7�E�@@r���Ę�~�Ӡ �ip����dqǫa���\?~�����>��'꒘�(��Ŏ�|��       �@��U���.m%:�d����R��?*�7��Vlj�p��.�G�$s��j�o���<�}!<4D~7u�����,�;xL��yP��> M�}eee��R�� �EDD�NW]�ve����}&L�y���D}j�'�>       @�ףc�娰P۽�9�;y��������m�b��q��O6��������������/|oP/I��4�S⢥cR��۷�t�}Uک��Wf����"� ��XƢ�"����5c�JKK���u�֒��.@m4X��U=�j��z�)���Ԭ����ˑ#G       �@�5#Kvϖ�9RTVn�G�w��:뵱-������W�ȼM���;��M���of-����/�ts_����wj�3.?��/���D>�n��W�w��`�C�����Idd�y�_G6j�@�����W�^�9E����͸���|>|�̞=�gۦ>ѐ��G}:T�̙#        ��w�l�?\(;�g��=�7}@yj�df
�]��5�����+�E%no뼾]�i��ymLv����`N� ���}aZ������^{�~�U�jľ`����|�DI����?n�G�@�b�qu<��k���3�y�{�՟��@3
		�V�Z�1�t�D]4�w��1�2d�ς}�'\���gdd��6l�>       �ߛ�jK��ӷ�g}�Kve�ȗw^%1�f��m�ɟ?_��v&��$��<MBC,f��-�O7��_4�/��xz_��������}aʳoK��d�G����)I&4{���#�c��-=l�����W� �H��)77Wbbb�y���)11Q�u�f�Y��u�cihh��Yg�%���&@�m�'\�\�	       �7m>rB���:�o��|Az7��}����[߿X��OF���T��d� �f�ѓ�����.��ھ�_r��EA}$�@��yP��b�||��&����e��O6�D�@�VTTdF������7���48���F74��b�Hll�鈦P{��-�6m��v�O�¹>�V���#7n        �v����o���ui+���R��L=��Jy��U*�����v������/?^(/]�Y�s�P�} �\�˓��̛�t}N���S�N�� HkpJ������$�G}�U5�`       �%8���8j�z���7��1E���ea��_�F�4o� ���!���~hP���J�CCdh�*e~8�`����}�?>>^����h^�:3�jp�cǎ�� 툦��)o�>�_�'�O��t���2�[�
 �y����m��x��q���k�����%,$D     ���3��������w���Z������k'�o�L��#����of- �ٻO*W����VT�``��(	������fc����Idd�����C���������n�O�b�MK�0�ڵ���p:Y�A���&lW\\���	w��>\��3p�L��E ���2\n���|�n��=�[�˜�̐.�	    h>���w�	�yB?llw8�@*��n^�;��||���ul�Y����̸Q�%���q��m_��1HBT�$�
�j���R�G� ��WPP`#�p���_TU�DW����,m��i�U�S�pEHH�#���֭[ˉ'��=��p�O��ۦM����)�h�@B} ����x������}��/,���\6�P    ���&5_	�5���s�P����n�6I���Kj|�Y~m�&������,h	̾0�y_8��:��n����3L@D�@б��bbb̛���F����2�.�c��������`�	wլO�}h*S�u h.:Nv\�N2g�.�ktt�y}�    ������é9�WX�u�5�篚":�1�:����^�kr�̺�{�.!�,�\�E�y���kժ�����+뎍��I�eHNN�����m_8�C�Yֺ�ג��|_7"]>Z�S������}���/�X�}�_�������>����
AG;Wjp�ڇ��x�4���իW{m[�'�U�>W�Z%       ��G�������o�*_n�+��<(��򤠴܌m-c�u�������h�m��h��?t����~�43�X�TT��<9���"۶?X�]��6��`���%//Wrss���t`�z��������ҫ�߬�uk�~u�hy쒳e��=�r�9��o֧��:&ƙ��}��잝�Y���p��j�c||�c|L��T	N�Uz�TeeeҩS'�&����>;v�(@S� ����1 �RPZ&Kvy>Z$�TVY勭{�'�    ��p_uQa�2}@s���;�o���%�FU[�#��t4���>��k�ޖ��h���Hs����Hnn�>^;w��/]/��U�1$1:R��ל���}����ד��> AO��LHH0��������`kyy� ����0_�IEJJ�׶C}�1����W�O��4���l�)}����] |���R�z�k�)�y��~��Bо�tIN    ���p_YE�<��2	f_o�'�RZ�1��!�^����t1{~�ZY��_�����O���\�>_?^�G���}�}��Jme��6ž��W+���i2�{GI����:�[�琼��;�h��w� =����'���&@��@��Z��\��j۶�׶c�O�t�*_�'�OiE�\��咁=et��Ӄ �mG�
彵�d�q���t��1+c�x�|2�o�d	�y    �Dϔ��_���5��}o��jN�|�s�xI���ֱђ)�%er4�@6�4�M�b�ïHK�됛]s������C��m�~�v��,�hN!�tk�()���H����S�+��GOHQY�dB�������������ҵ�@eN1�����P�֎}�
���p�s}�iӆ�2�T���K��^ |z p��1~i�    �Nh�E�~�yru#05��cy+��dω\s�I��}s6��p��}꫰[s���4qrq�4����5�]�9����)�+,,���X)))!��MG����Q�p���O0���	GS�>�X������Q�       ����;��o(ܧcyU���pZs���|���_�����;܇�� '�@��JKKh���Utt4�)�MkG����?�=�mP�h���y��       ��>4��������K�����k�����L���ᗘ�ܥ��***Oj������       ԏpܡ�w��}yo��௏W�}4��?� ���J�:�W�UUU��
�|d�X�=]_��L���_"##��n		1_����r���Dc��>       #�W�{��~�l'**�I߯
�����Zh ����t�+..�`�!<��[OMȳ��K�/��V�;4�t?�VQ�h,_�'       �5��А`{�����p�v@�;���d$/Z"N�;[�p�o��O4�/�    �!�u�X,۬V�&�����5$��vyveEUQ��Rj����KeU��]�"}l��m�X��XR  �} �x�� �(--���h�}hq��Uhh� �wD��^�����E}    �c�Z�ٞ�}f�ZT���/z�G=Y_��O����L��c[�b{&�$  �����!� �Б�f����Z
�<�S�j��ܵ�>�)o�'    �a�����O$$䵼'����L�ɞ�<�-�/zzA�|&2)Bη��F�V/�m'\  �_"� �#� Ю}:�W��@K��L'J4��8��)=>zk:p�/�    P7��g{V��k�������wyo���]�#2�vnV�=O���v�v�X�  �w�}:�巄� 1�} � �����H)..�%���c+WكSv�f���)ù>�    >��"ևr�ߔ�V��w���{�ؾ<����l)���*��Y,+  �����T�>�} ��> p�v�������P3�tZ�tDCc�"ا�I����    8���U�e)�U�����'l_~�����QQY�g�Xn  �W��k���4A�>��N���|�M볢�B wi�(�}    �}V�.��ȏ��zώ\�?'�z�aۗ����[�ˋ��  ��> h�> p]�Вhh�`�ѨO4�    ��V��sy����]�s�O�37����W�f[�H  �߰���BCd����^W�}=R��X~��ye�Ȭ�v����w� 7h�$<<�`��raa!�N�6{�.,,L���������n�E}   @P�Z��%���'��Z������=����#"�P  ~A�}����~t@�R������g����Y,�.X# ��` �A����ƚ��}����Unn.�)��>"WCS:�Wá�@}��4ا��5��P    @ӱ��J��Oܹ]�Ś���%��g�VYe�E$Z  �_�p�m3?3�
��?�[8��h�|�e�l������� 7h�E��ih�1�M'6�*U�|L�1�*/>��o�R�%F�>e���4ԧ�A�\z��ګS�h�w��	 �ԽM��R�u�**%��Ld�ɾ�<��.�{w�)}�J��8I���]fF��/����g���w����Ǡ��n���R�b��:��1;vGsd��#.o{R�Βe���~N_m�W���c�eB�N�y�vKiř��_���;5�����
K���)~�hX+[ML�Ն�E;�:wWz��ҧm�����|Y������'#��;��o�/�ťnߗ�����v���0�V��q��8�i�WVUɬ�v�7����~�dp�Ts�im�'*�X~��+��,���1?�����&��,#���6���#$��TrKJe��l3Rj��ò�D�x�t�vo�!u}�tt��.!��e��d��c�.o�f�~�~� �����0kŅYO�wH\����8�g�L��X?�X,�  ���b�������` �I������P��T_�/Z*%�z��;�j���F��:ՠ�*�Z�48u���o滋�Dc��>�����U�r�D����X�m�#/-� ��r֠���)��9K���Lw��������9�ǹK\
����N�����Ͽ�r8���L��N6C��K��7n�.���f��;���Jm%��8U<����҂3?�t�оr�9�\^ONq�|�i���l�|��� #�sӨ���i�]��y�䉯V����{��玨v���=���}�BC}�u8��7d��l\���.���L���v���K**��/^�������ޭύ#�KEU���z���k|���E.�K��������t�Ys C�Y�M^[�I�ʚ���_ێ���B����Ԟ��c�� �m<�)g?5S�\�*q��^p��$�}p����Y*���z�i!r��{a�=ϝk���vx�  ��@u� �M��:K���HUU� �H�Z�ʼ�<���c�4\b4GDDx�#����U}�?ӮO7��'׍H��Y'����brQ����kΓ�Sݹ\�3%I^�y�,�q@nymn��%��7�ף�K�>�r
��n��cR���o���:�:B}�~���C�;�fx�\=,]^]�Q�h��W򼳩]?����~���+�)���Nw�L.��D|E����;�q���c�/>Z(�B��������z�|����;�l`/���2s����?��n��� am�vnkN�M!�|��g�w�/th#��%�Щ��+BB�=yw�	���=}�ğ=s�X��D,��!  ��p_����[�
 �!� nr�k�"w���-������1��)���e}@s�ў:��YdX�tk�dFp�iW�;�b4���u��y� yr�9ft�������N�l�^�+(-���9�C�t`O3�NG�ιc�����uv��v,K���qrܤvs�3ڐNm�c�IGW��B�g|��e�w5�;�_$�s�].���y�tVt&i�	ҧmk���5��� �ar���Mgd���;����h��idٞ�M����2[O:̹����쪡}����:*�גc���^b�x:[�|�n��4�a�yi�wH�7]�����ԱC����<b~~�����"'��m���dվ�f��*,���(��b$�]�\�ޭ��[=��t�P�
��_]0Z>ް�0�%�j����S���ܧp�ӷX��X�`  ���?}�F�90��.�} ��(**�`��:=z������}.).>�&ttt������=OP�p�s}�ܹS �%ҐP]]���M6c{5hgw�������^m��!O_1�Z��[�7����ce�E�Ż�?l�aJ���v�[��Z׿}y�G�ʹϾmFv֤/�.�}�tԨ��M7��B(�#E��K���ۛ`�ܕ`�v��**�-GO4x}����X���ϖ���&I�dB�Q���kF��߾_�4���8 ;�tI���0��񲩂}��a���#�拷i����}˛���~�O���0�֔���v�{�W�i���-�k���1��q��a����1�㱃̱JO_<޶O˛+>���w~pI��{O�ʟ?_!��f�,��nkX�vr�������-��Y��2�
����j��yO��� ���1��x��m{�/  �{�oWf�����}�E?��� x�> h��g�Xǋ����#G��Z\QTTd�j����)���"##�< �����H޸ez�`����5��!1N��jJ�P��_|k�g�j�>9��we�3�xK�� ���:CL:���Ӏ��N��r_���9�}a�Z���q*�{u��h�1�,���.��3s�Wf�q���Sz븁�����.t�Ӄ9�%ĘP��Q�~�P
K���k{x�Q�Mg�='rś4���T�U������S�~�n�=���=x��j�������t��/)�?\({O���߾7IV�Ϩ�3D\d��n۟�C}�/���\�ކ�!C;���O�y	�ԌsL��h���Γ�v'���}s�))���X-���=q�W$r����j��b�   �oh��1^� ���` 4REE�x���)��c��[iFF�zw��	wh}��Z�Ǐ7� �H_���rn߮&ئ�t�hF��{hH�y,�v|ԍ�5�s�K��{�3�W?{��.��#g\��]�-kh��`�	�u;�r�>�lP/��^�$'�����:o?�c���re�?���/?^$���p�.���dF%��Y��p�s]�c�W�j�i L�}o����m�~��.15��~u�h����7]?���DW��A�6y��LGڶO�3�ms�j�_�2±\QU%W�<��P���/Zk�%�qF��'.�du�`s���c���s�>i��Z=�\a;�]د��=V�i�2y���Ͳ������_-@��Z�̋�zT���X��3�UV�Z�R    ?@� I������C���V������T�V�(D�|9�׾=�O�J}�^����td��A�w�
5]����j�G�Kvy%e�O�����s�8�?L��s����9�[3Nȉ�bim�uL���PuJ1ݶ�ѼB�q<یHu������z�}�c|Ւ 	�)���w��@��4�y��xd��� �v{ӟ���l�Q��}�F�u<	�iX��n6��Ռ��M�j��L�%<ͩ��;k��Ns3Wmq�4z���׫�9�([�v�Z�^6:��z~?g�L���щPC�C;��52θ�?~<n�cYǄ���g�
����uަ��/����Gv=y\��a���[\*�'l�^l���M��ǠS�����{�A��   �����i�T�=�@@� I��?����	��+Z�.]�c��>�ח�){}v�ܙ�D��@u:���S�0��ͣ��Nbvo��"����/�`:qٻ�]Կ�tno�i������g� ����t4��]�qëct�_5�����I�\�����|���R�t�;�*o�,(r�TR4�>O��N����1���j�jmjw�_�?�,�J� =S�Lp����ŷrͰ���e��"��p�\��,�+��1^��E�}j��l3Fvx��������U��?�#m�����i�E�����2�����G�0�v��m��g\W�z��p�v��Dn�]&�r�9�*&J�8T�t� ��#�O��?)V�}��W�{�f�X&
   �.""¼���t��*���m����㭪�4��p�� � ��!=�H�����\ٿ������P�b���Tll�lڴ�'۴�g׮]�O��<��ܼ��v �����\Q����^��-kg��*,-7c|�?�dw21�ݳs�ϖ�:��i7-�[[�-���;�[��G������$u��������v�� ��@�S I��狽������ڵ��u���}���2���u#��Cs�6z[:��_K6�]�����u��i�e��#�Ԯw
ͭ�Č�{k�VG�O��jhQ�#_�)����E;ʡ�|i�7mǖ�N�7>�w�Z�W�8��
�<��Ŷ��W��ɔ>]��g����F���ʶ�r��5�5��ٻ��*��  �/t��I<�wa7�i���)}��y(**l���� <����H�}T999f��I�����􉋎///�;v�d����8�ɣn����o߾]  ��m�\m9��t�7���ֱ�������l���`�۽C���Ż����q���j��ctud�v��@`��x3:��\ڧT��ܮ�ӱ�}ڞ����BA�i����eBe:u@ܗ�'������N�:���O�� ic=��J�iTG�8Y}��ISJo�ڶ?�:���3/>r��5Oi�<_�F;��J���Ε:Z��)f�m|�	-�r
4j8�y�e���
�:����]L��D���玐?\(@cX�����ς~�s�Sw�O��7m���   >�oa7{��[����C}�?� ��`�������RXXhZ?3������Tbb��]��g��>�c�vc�����8���ի�� �Jk/�RN�p�.*�ݙ��o=S�c;Ն��=�f��F`fP��Z����	st\�Ү|�.Xs��4��p�×�x��r|O��j�O��ݾ�`߸�-ۃ��H��0#[ݑW\*Y���T<����`��� �h�6�����:{c�G��}b�L��E�غ�����/,\#��p�Y֠���i�����T48h���U� ��o�n�#��i��7�����&��+�;������1�׹j_�#اuJ���/)q�G�뱧���~ s��L�x�N��U��`���&�
�igށ�M�@`UV�c�b�A,"   �		��8Z}��������o� ��0�4(���%�w�~���}�Ҁ�JHH0�)_q����t��j�� �1)^^���j�}�yO���=TgwЃ���ud�m���s�U���:�����w7�ڕO������� �s�M���>a�9?�g'y��3�k�w��v����	o5����o��/?^$��q��O!���L�aO|�R��F�W�o����v�q��6��/�(���fYG�z�S/,Z'?7�t�S��h�|i[gS����W��X�b��Z�:f���Ǧ��\�����j]m�@���dW���q̩����[:�0���5�����G��o}!�[��G�ݫx�}J��wmM���,b�B   �3�v�u�-�/�G� <���Y,s��Uvv��ܹS@p
����碣�M�>_���ѿ����>Q��O �5���4bVE��IZr����&?;��Z����/����^r�=���!%Kٷ�U�u�:��iW>�U�������_}l����f'��̧4\�<�W����SmjwM*W�[�2�tn/û�����/��W�-�͕�y���	�g���X��f%��mM��n��]���T[�j-{ҍ���\��j�����f��6��������Ҥ�SW�ں*�/��S��G��i���}�N��ʩqܪX�y��sq���]Я[���0��Gş�<�c~��.�W�+O/X#[���%V�܂�7�X��'lZ�  ��
�5W�-�/�C� <��>�}d�`5��蓈��R���3��rrrė�O��^�����g���' �ڳWN1'W�?�w��U��*:<��rY����=�fv�u%����|��>̫�>F7��X�˒>m�͸Ԟ)I&�bׯ}�j!���O��
56d徣r�����6���һ����l�����싴�檡}����=����6�g�.�	f�W��O��)�U�W;
�i@W�s֦��J�[���5:���h�tƱ�[�ê���B<U\#�Ys�vV��65(��S���(W��_�>���W�U���z�n���:F�{e� ��������6����Oݽ<��g��E�   |��a���������4lb������\�9b�Sݻw��Q��TRR����;>߾�>w��%ݺu�>Q��>[�j%����?hHGG��M1���t��]�~U�њ���"#�)8w
�/-�s��#�&�d��v�{a�鎫����m�Da�l�8����݇M��ܾG�j�>�nj�.��}�.X#���X����r��5�F�w��}���X����7c��M�x��Ι�}�B�q�yfYCu�{u��F�SG��۷�c���;������Vnv����u#��O�/��r�р�'kt�����rS���a[}��d��t�P���QGvm/��;"@C,byMP+�X߰�|   ����n�r���� i�D;���رc�a��ի�)T��)/kG�E��'�c�Ϟ={R����g��6Yn=���N��+z '�t��t����.&�MNQ��K̀Lchg3�YY�u�vt,��ӽ�ԸK�����o��x]�Ֆ\��|� s~B�N�R�ztr��@цC�����n�Ni�s뚜 cm?��S�ei��;����;G>߲W�x��qH�T��[���:U����l�{'w�^/���;k��ݓ�J�v�����i�Km#�]q��t	��tz�ۤ>������3e@�6f�Z���l�O�T��%Fy~̩9j��q-������]k�Wz�K?���wO}�Zn5@�O�@���1r�Pۑ`Sޓw���b	���D�  ��h�m���RTT��GEEIii��o?���H)++�} �!{�> ��8qB�l�"%%%��S�SAڭoժU����,�C�s���r�EQ�pp��իWK^^� @K�]�>ٰ��e��ԍq��
��(�+������=��h~�/<�x]{�O:ڥ�ޝn�S�oI�����wv�׎}�9+��@�������{��1��dަ�&�X������Jld���#A'?�l��4�N�j����[��8�}J��m8�У���?}�\޸e�Y�1ҷ�h����<�wV�	�6�M��z��	�|�����E����gS�ȯ��wj+Y�x�o�cN^A���5:vk���z��ʤ��:�rۮ���������//m�5�<����z�~�d�Ou�}�=��=����F_  @����w���u���[��Bş���Ik�����#� ��Q4���ѣGMxj����3�<�����o��{}nڴI�B}��� _**+?�����e�1�m��rﶭL׸�FvSû����ro�c����.}��`ޘn��y�w�V�Q����L�;I�;5Y�edI߶��ul�����Wڝ�Wg�?�LBC,.��8U�~j��$�����UC�g0�����jh3�ٝ mm�l�eF��hTu��ڊMn�ӣ�ڛp�]�~��׻ܾ?�E�o���A�np�Tywm����z������2�}_�m��{�$��㏵;inqpt$x~�Z��؁�j;>��]4V���/|>
u�Z,�џ�>    >G <D�(�:�tݺu2l�0�S05��
���rY��q�D��}���éO���~BO볢���� �>}�p�E���e�9�OW��qW��i_���::���XӼ�2I85*r\����7�̨K{0/��Č�˲݇L�Oi�?�Mpë�3`�Y�〼��;��؁fY&z����sAz7G���b�d���?Z�yg���-�On�ܜ�n��7q�<��2��q}�.����m��eyw�ЊA�����׳�i����"����ێe��rM���;�ͳ��
K�婯W�c��m�5Ly��^MR�h��R^nm�N,�2_,�    #� M���NC2۶m�H���Mp�+++��@۶meΜ9&<՜�>�n�J}�����LMM�ٳg7{}@��t�ja�F�kt�O�u��tq,痔��:��X��{�ѳJ;��S���O�4�SUχ�t�5���y�����Uë�O�}6�G?].3�6�2��y#e�-wk6Z�M����$�h�A��}����0X��d�˷�.���K�BdX�\9���s���o��ǲdω\�8\�68:����?sV���z��9y���%ا^^�����!��/-��k|�-��_ڍY�ݝ'�WyH�7�V>d   ������c�>��e˖ɕW^Ip*��q-33SBCC%&&F�͛'��������@�Κm�i�L�.���&��$��ttퟦ����C�]�ф��d�!G�O�Հ�]C����9�}��}Ў\v�����A��k���5����!��g��������X~k�V�}��n�����u�5��!1N�x|���T&��b¬���rߔ&��K���S�.Տ��T�[���m�~���?�v	�fY�o��i>�_�mػ�);��=�_��r��t�rYee��_��{O�Jک@����v�[w00����я}�B^��\��+��\;<]��,�A����ӣ	�=�c;t'	    ��>  �]�֯_/�'O���DFM���3~W��}�嗒��/���������ꫯ��>q���0y�����U[��@�J�+L���a�5`�����yϽ#�nt�ӎy4r^�߸����잝��4��y<G����RJ\����1.����k�z���!���?�0،+���Ԗ��a}͘i���ns{��nc���XL(ꉯVz|��8&�|�S.=��|� 9����37�8�Ү�s7�qk������M'75�c�9�xlo���ͦ���뷍$/.v�[�߯>O"BC���j�9�F;�j@���e��x��2������\��[���]��J���f�珔�1���� ��E��m�)    �C� �CK��hW��˗˴i�Lx�G��i'�V�Z�'�|"��������9k�,	4����[/3���_g4�M��ȓ�x�K�̛ҁJG��2z���Y��(�>����[�>����km�u<�?�Lf��#�F�j��+�T��׳���.��<.��\ܩc�/4��4\��H�A#�rfK���Ϯ����_��ѵO���9i��q�RAÜG�f����^�7�:£'י.O~�R��%�G>]f��z��5�v�a�F;ύsW=g��F��[���S���ph�x�v��������:.{�ҳ���B^�vS���P���O7���g��og/��v���d�#��3�}�&˧�w�\��&������G>[.��t�Y��a�f�*p�E[��   �S� �C��EKs��1Y�j�L�8Q�������<)..���dY�t��b��I�&Idd$�d�;��>u,�ѣG���>E��s~�_^3� �J**��o~&���J�Qú���� ���X>\���Q�r�����������v�.�������{�8ƥ��J{����>��9�^�NkdHc$FG8Fw�#��ĭn���ٵ��q��EkMPuٵ��C��Z�zs�֠�V�%��m�dtZ����g��l��j��#�=�Z�놧W��ӅPi�@���g��i�W�c�y�Z�lc�Fj'O���g�z�.r���fY�?w�s�Ü%��D���࣎���gK���奧�_�s�{�鵹��W�P����>x�m��`F����nh��FK����Ns<�ǡ\�5���P�j��j= �   ��� �j���dϞ=�`��>}:]тLFF����H�֭塇�\�t�>����Duy%er�S3=^�{6Δ���@���Ŏ1����u��ߛ$��C9���~@�62�K;�q���r�;_��}�g�ռ�KwמE�v��ZC���y� sr�Cs�ʓ_���T�k_ld��=iX�]ʂ��#�w$kl N�8^{�Oi(�)�}�ϟ��+����������uNcxO�׶����q���Q�|rL�L�����]x���f������������Wʏ�t\�#�����1Y��-�؈pi�'{u>#��a��_�#+\��{$�@�}�]y����Ki��{'7'Yj�-��3�N�ᡡg�k:j�ә��h�����sPz|���	P��ҵV��ŒO�   ����&@�(�4��q�#F��6mژ0Z���l��m۶2o�<9r�?G_j}j���ÇS�AĹ>?��S��O�Ve��ho-�w �����;���er�.�˓�#�S����5���Jyv��F�']��[�״��	�)�ULT�����f׾�(�/\#�E�3E����z;�u\�}���a��ٝ��wi 큏�Х�tl��K7�gi�p�t���h��F�W�s�O�8���}ME� >�����f�*������h��������ۻC�}�������1f�:��1�zj�v��`��]0���.�q@�NZG@MV	!��2k���    �;�  �4��k�.��/��o���2A˦�8�fF0��������_�7�@}�@�O D�����}$�zu��'6���KMڝ��.yf�j��j�=�a�_�G+n8tܥ�k�x��æۘ�o\��]���r����ˏ	Τ������{붋���{w�v��y#�y효����fi
���Q�M���G�ڽ�AB��xu$��'�t��yG|X{y�w�1��ġr��w�<:�&��c�u��썻�M]�v�� ��.�7��m]�TM�m>rc��������-�/{^�Q����XI�fb�3��v   �5�} �!	H�>�D�kݺu2f�IKK�+Zw��q3ֶcǎ&4UP�߯�k}�]���g׮]���f}���T@p������+��IO:tDZ{�/mb�%.2܌�<�_$��d�PPSЎc~���q�+�=����V�E�{��O}�ʜа�Vo5����g�ͩ.�̜C���~�b�����>5��t�3o������)ޔWR���vMN��:��Q�m�M����g��W(��1�ME���y��I�����t�L������4���t{���M���\���X���Y�ގv�l����u\ֈ0➮�O���   �[� �C��`Z�ݻw��}��z�����Tff�鄦�N�̙#�@����?�>[8��,))��s�
 ��J**囝-g�- ��]C��k��t��YXei��%U!�b}    |�` x�`Z���"Y�f�,^�X&L� ���СC��]�����3�j֧�     �����s�U�d    #� �`_ee� -Ձ��>�>}�H�6my�����H^^��������eӦMH�ϖ͹>,Xp�ِq=:J~IY��z�$9ΏLk/����]���|ٝ�4#1   �%4^�����
   ��� ����%
-�v�ܺu�|��'���P�r�����i�_�u	4�g�U�>_{�5ii^�yZ������5��'�Z)��L���v���RYEGc   ��UUJ'�k�֎b�e    �"� Ҏ}t�BKWXX(�W��~���رc	��:�T�]�t��\���%��3==]ƍG}����ڵk@�g0�,(6'O�m�,Q�ar ;_N��   �^Uo�k,�G    ����4�G��b�޽����˿��oY�l�dee	�Yg�%3f̐��dٳg��]�V���/� /����Ԭ�5k�HK�+3G�0gI����}G���0��<|��-.�A��z��;$�ɭ�����D�u4�{�Ʃҷ]k��;_����,    �����ˬb�M�>    �F� <�cx	�!����Hjj�:T-Z$eee��ӦM�>}�����.������%�>[��Z�v��������%�����:��.!V�9g�9��ܥbF�   ��j��s���,��$    #� �Ё�ʛ�Z��	M�7�Z�b�@���������|�2e�<���-ft-����)�&M��{L�    �a�X�J�����g~�#�Sxe�8	�_    �#� �`����r���5�^�z�����AG�_r�%���b�o���dddHKB}�����k����    �b	�
��3�u�)    ̀` x@�}������"S��{����B9t���i�HZZ��^�Z֬Y#-����>�J�։�)�Er$�@    �1,9G���j�,4�   ��@#�����UUU���|	�A�� Uvv��i`��ϖ��d)..�ٳ[�k���YRR"'N���`���=:��n�f�y쿒]TR��Q�a��G���-X#'
�k]�#�L���w�'�Z)��L    �1,b�j�r��V��=�M��G   �l���>}��'Yll�yɟ��E��@#i7���J����t��#dɒ%�;��v@���$::Z:u�$�=��{}6���c��ٹsgy��G�%���Hs���Qa�r�9����}���`    4��������ݫg�Z�n�Xh�  �\��CRR�9yoy���#����@Z�jeNޒ��+�����@� ),,L***fV�U233%%%EF�-˖-3���?���� �����;��	ABpww/R�n�[*m���֍��z�P�P�hq�$X�"����/�af�$W�ӽ;73�!g�w���=o�ܹdggGaaaB4��Qn��G��au���@^N���`GEť�rf6���Z��0�ʈn�X�g���0�0�,@�WTt�睜�]�L�gd4�������︸��W�"fd���}�0��}�0Z⩔�����>}��[8�___�?>988PϞ=���_o�����)_|||4�>�Q&�=]�!4"$H�W����]J�5����v�삛?w3��;�C ��13Zm�2�0�ѕ�ͥ�^z�^y�o�F8?�A?*#.��0�0��ف�m������ӳ�i:�Jԧ���E<6����D}z f,�?,�c����Q�]���3ʞB<�w�^�63M�~�����$JѾ�����͒��>�����	Q��ۧ����(؄����ɰ��K�
ik+Kb9�
lύ�KF�$+���k�����ذ��⍴��yRZ��a�a4�N���qkѷ��(�x��a���BG�Z�S�@
��V�.�hkM.v6TRV&���t~>5�N%�Ҏ�	-=jKKr�)�&dK�K1��);+K��M��N�.���4���Mj��[FѨ� �,�����J�.���h/�Y)Y���#�y����i.q_S����ũ���1��.��0U())18�0@����i�вeK���[� �k׮��oj�Xp��U�'���P'��>��վ�г��(����{t5��I���T:��NydeiAn����� `�p����1�X��~;CJ�!�>�d#-9M�0�(���饗~�W^�IO	��>�He4�t�0s�<9�'��#T���0����4�|G��臘�m3":��sF�������I�@�6�s[�6��l)����.%ӟ��RrV��1ǆ��gG��-�D'�\%���h�p��+*��R���I:x1��$�=0(���K�N��c�`߅+���;h��Db����=6�MoG�nΕ^�N�F�8E_�<B�E��-l.Q����i-^��a����<��e���2))I8���S�2MGpp0͝;Wt�۵k'DS\޴n��O��	�isd�1�ԕ��:Dn�%%��߇諝G(�̄~G_O�t7+"D88�7}�>wY1%[�����ۢ���k�ӆҮ�	�%j�aFA�tm]��gf-&�,�,��,�a�
������G���M�~���;}0c8��?�n�~���B
97�ooKm��*=[�N��ā�ΦH���Cf+P����l�I�`��ɬ�4�W�J�n@w��L/��%�?��R���+�π�o��{h&���_���ib��I��n)���~���1Ű���m�������p}e� ��w����x-������i*����e���aꈕ��p~�2�c}�SOOO�ׯEFFRz:w��N�:Ѵi����]|���^1����|�������E����ۧzAV�w{�7��IN#�iN0����be�f~���Y %����/���B�L*|�ޓ�\���Ny��~n!�]E��%T�;���o���a�a���H���h%�rg>i�'>/++��n}�TeNώ��-���I��_�"\�P�33���r�`cM.����L!>ԯuKjY�x��I��M�?ZBq��4?�[�ӊ{�Vr�3e�_�0��"6�YV2/��w��O����_�0�\H�VR�Ջ��g<z9��_� G{��'�,,�˹���@L�5�O��E��&�G��;S�I���::�L���������{��N"[��]P(�9�Yzp>��o|�W�zS ����p��YkHr���O~���a��X[[�_5.��'6Q�P��F;�<�%1�D/�B'���t��Q���'�� 'Q8Ѝ1B�9MMM�O>���p�lZL�Ϗ?����.l�F�S@EY�ǖm�Q�g�׻��}L�ό�@/���leLj�Ȑ 1i[��FQ�1����W�?^�a�a*��%+��L��H����,>�L����0�� ��iC��UG��7F֩�*~�]�=�?�
�%;Q�v��e�4/5}5o�Aԗ_\B�G�������Ԇڵ(w�C��5̠i_�0�l/w�=]�ѡ�?/���������|��қ�Ӈ|]龁�R���9t��k*�܅3��[F
�8����6���$7p�!� �ϰ�R�Z%�?��i�!���M���ıA.tW�����n�x����wn6r��qvv�)�+�x��>F^���a�XH�l�ż8՘��Ⱦ�ף�<)�ڛ呙�)�lv�֍\]]��ɓBT�4p�<y2u��U8�mݺU��15������zZ����mc\�ʸ`Ҭ��t�4Ξd��2<$P<���J�����c�tnώ��I�@�_G��Gd�/;S���ǋ�Y�@_�y����0�(t��\���#���G������0S��t�-��yk�>��L=�8Oc.�E��e}��׹��\{� ����L��ס��ri��EU
=/��I�"B�I����A8.�}h&M�bŧg�Ҙ�#T���v�Ta �R2���;��K�;�!K����ѼEҡKI�>'5'�n�~-�X0W�R�ߏR�jfX�@���%���9Yj�.&Vzυk���?w
�n� Ā���D���+��7܊dl�cccK���㵳��2���>�a�:`cc#n�|3c�ړ��/��Z�nM���t��a!�bʙΜ9�����K�.�h�"�|��.B�ϛ	�Ϛ5��>���;JH�������Ĝj_��i�0L�ӣ��x\y�4�gp>5����I��-[�^�g��H#��߂�}�0�0tD�e��Ь�F���%�!<��(����\��aS)O�:w5���ذ�U��,�J��Z�/8��M��ƤA�А�
���3�?�ts%Q����C1��L<��	"�����x&M�|�+	Jʵ��~���������u*�Q�|�;�3�� ��>v��
�x��.�=�������^O��&%0�c�a���n����H,���A$n�����؋7�o�ں{��:��>�a�Z�R�p���!�a��������AC�⩔�b�Oxx8M�0������Ǉ�}�]*(( ����'�h�>n�L]�vv�`W**-��W3(=��#��v�M`׆#	�B�֮�;ɝƍ׍�a�Q:�siu��L�WH+���Uq6����<�a�nN�Nf�� ʸ��G'�\��|��Չ��{�[_\j�?y���P�t�����;&Ш� �]8Ӛg��3)��%e�IsZn����7~�]��˸</\��&����C"f�T�9��]��5���}�kLj�-*��VRZ*ڇR	�o!��8�9V���<)�}�߽��>�a���}�0�n}(��*z��8wRSS����z��M�O��Su��֖Ə/�S!!!�s�NZ�d	1��}��y�������YG���]�vq����l���X��Lr�i�,tT"�CY��]0C}<�S���v�Di����1���;(69�Ԇ��#�kM�.b��M��Oq3��ҹ�DvJV^�?6�٨ܶ�o���e�a�<:������we���&� �Y�KA$�a3XVL\4�����T<b�i^<������ߋ2��~�'-�m���tu�?�AS�\A1U��䊓��x�O7�6�`Tb8�W����(nv$7 �D)�����C��ў>�9�fw�Je����6��_sբ�����-*��a��1����Y[[Snn�l��1�#�?m۶-����ѣG)=]���Ơ}��4q�D�֪U+���o��5eL(}�lӦ����}֞����!�e*���Ǘm!5c!��?wy9�������M�%:�<0�Ꮵ��Fwe;P���ee8h���}q\?ߩ-�;�҅k��{T���.(�,�w@8�6i �ZYV��S����=���PS�@�jQ�x�?��!��H<��\������0�0
EGTZ�����z��Ӥb\��p���1�T�Mp��ߺ�H�jh>���-u���W2�W)ꚑ��k����c�y�����&�W?mY!�ԏ�k������a-}5oMo/9W�?]��N%�N4��H�۪k���=(�⭎Ԝ|�d����Z���GNӮ���ڤA4�G(�o�O;̣�6�O�Rw�mE�6��X���|q�ï9VA�i�{Ue��z����Rb���\JNN&{{{8p �?�����������4r�H�ѣ�DFFF�ҥK��9p���>����D}`ɡ�ﱶ���獩����Y��524������gsF��~%��g����GfS���Ṷ^n�̨��+ȗf~���#�ޞ6���w���U�O�q�щ+W��V���4C����ɑJ�6 �����0�(��[WR�������p�R!�O~<���;�j7�0����D=})T�?6�}��`�?⧷�5�e���Dr�8���š�%H�6��)��G��u(��Ż^/D~�a~�����/W��I���X>΍�Ć��^y��±������V��f���	hFDzx�f:����[�è��^KGE��{G�y�0L���>�a���:.����/c�a�N^^�pG._�N��+WT9O\/,--�gϞ4t�P���²�����C�n�Ճ���}�;���<`¬Tf��0?O��&�'tnK!>b���t!hÄ"xc�^Q
��>��K��'�%�=���ǳFD}��y/�Õ��nI�:Ҕ���	�Y���Y����t��U�=�gG��v���3�c._�0�0���N����r��c���	UYڻ<�a�����R�l3�0L����=<��p���޴������L�������b� @@w�b"ɍ�	ׅ}][� ������]�k9�XS��[]u��������0׳��i�,�a�7�Ċҹ>.�fߓ�[@��=.�/�eV�yn���b�9�q���T�}�'zu�@��Og1���ٴp{���^!�T*������$e�s�Z�W�t�'%����9aa�0L���QAA��1�M�.W�^%+++�����'N����4�2(;v�XQ����O8�%&�o�G�p�4��1c(00P��e˖�豉�$�#C��IƷ7F����~&�l���:��X�� �*���m4�SQ�vh�V���molXk����#���Ng�в�'�+�X�;�ӥ��]�<�{|Z0�'�����I�ȏQ�A��U��8:(��EC�2�0c����YY��x棱��~,�T�����+�؜�a����N���MoL$~�ޭ�آ��Qd��MN����VVR��dceip��8����v������n�e����r��OrL.mL���L���.ec:ӊ#��B���e��������U8��3�+�$��<2�/�$Q�r%#�_��V��y�����lR
���"�%���#�]7z|X���  qIDAT�,}7�.�B;�*�۳���̾�n_~M��Q�q
�t5�'e���4',�c��kkkd�Raa������Ǎ��������LP�� 8d��i||<�9s����HKѐ!C(44�<==i���B4�4/�>�����`2�ށ����Q��orû"�7&�����.@�ci��	���b���E�bp��+(P��u�+M�c��w��"~~a��J�>=o�����
��p�ca�<���!�%��X��0�T�ԍ�T\B;���`l�;OĐ�q]��T*�����jW��a���ۢ��kʎ��eh=�.Ptޢ�B`%W�%��Oh�(���UT]P+kN��7���{���`>���G��A�	=�����y�;�#/(/��A��B�׏�؍�x�	�ůw%����j�.T�|��j�7"$Ȱ��s�a� ��a�e322��C� vl����1>�+J�2MG��B�+�uBZ���	QRR��ƊsQ�����N�:���[�l���ϓ��*���ξ��gp��=U��֭[)::�䎾}R����{��-�)Dn'���P&�[[��{҃��������R�x:������?�8;J9l��3���V.�E���i��]<BėSpc���>s���ѽ�L<͌�  �a�aF�舂u�;]��h~滏m ���K.Y��J��&cA�0� �����Q�iB�dgU�����y��c���(�$(g~9p���fg�0Y��Q����9��]P�2�M��k�t*1U���kݒ����HB2��q=�j����}��PY�o�֠ς�uV�P��ϼ���dx�e��->M��)�m�70��B�Dr�(�\�5\�������>*Ɯ�R����4>,�c�1�.iZ�Ǩ�B+;ҕ�Q��JCH
J��9s�����,4��ģZ4q��ܹ3��Ӈڵk'�Ϯ]���p�e^-������+���)3��g����q*C���%�g���%/,�\l1�>��!�[�G3�W*�����_�7,��f��d������ӳ��^�䶵�����mʇ���W\�x�6+����\J��l"'0yY۲3�!!]ޓۍoMe]�B���qߴF���'Ή� �a�Q)^�����>�$#��)��>��3L��]/�,�H�G�0�w��i=9�X�y�� oj��.J�:�X��M��WF~���ٔ4:��F{�_����]~8Vl���JHμ�z'ui�%���oN��RjN�!y�T��������}�|V/W�}.Al�N�J�hB
��x����ܘ�5�����#�����:�7���}�������E6vt$b2i�2�?i�b�2�dꀅ}�0&@�Xrrr�a�@��QV�pJT�pJ�^@u��eqN�����Ν;'J�6��ds��ݻw��={
����TZ�z�"�9yyy�<�����W�}fs��	���U��>���ű)	�@r��ޖ�?<K�0�����(�?�^�8H���k�P�����C�TT"��%>�\�ӽ�������7���4���/-/��LjN���dcc�u�q2�`��Zn��XZ�q�����w��vVZ�W���E%�tC�rr �a�Q7:�Y>��Q���{��T֖�nO~4�����ϮV"�0�	�:��l6�\[c���#�Τ�7j���|އ[��Sq�7�O<��]+�y�7�Z(C�X�؍����a�666�����%���H%'.���w�R|A`Z�hA������)T			B`%g���E�.]�w>�����ʫ\cJ�::�P�C�K���'��}6jm����}��3ɉgG�1��0I���YQ����]ۉ���{���%=4$B��W���MK�b��T��d��z����I�א�:�[��ٞ*��� 69��LRf���όCamq�(i���<-�(���b���%j�}�(�a�a��N�dI�G]|��M��)�=,+�^�g>
().��4��M�ӎ{
�0�0�Ctb���a��1�T��,)U\�0�(����2r��U�h�'ʠ???!FJKK�K�.QJJ�,��0a���+J���i�V��{��ӧi�ҥ��0���y�v��\1���N�O�����cy����ϐ����kI������i�W+(���_���HZ��L
����[<���Xz�͊�
�~�,B���m���[�Х$
pw��G��V��B�ߣb�\S���Q���l�c	)$g+h��f�u���ח5���w+�^�R��a�λ�_����l@/��_I�w��c�aFS���W`W<�����pL��^y�Y�����۪�pAq	=*��a�a�aF����a�����A���:.� �K���N�]��W8�///
		΄P�y���o��*�}�l)R��P.nǏ�}���ڀ���=����2n�@�s�399Y��m��DVVVt��5:v옺��І���$�Õ<�ו^Z������������O�� ~���_6P���T�Q�7~�g��-�k��I�ɣ��6_�adH�8����w g�_�*=\�����<��������|ţ��ay��Iό�MS���;��J��I+��&�aFti�B�ۉr�{��uS��tAT���%��_��o;:�{���4{�}���Jt�ORY�=���}�0�0�(�1�T �"� �(���
�w�x;�/��*H$R[p�^�z�𳷷7�nݚ���E)Ԭ�,!��{p��Gċk����(� �<<<���I|[p�;y�$��8���1l
K�Άbh�e�Xi�}����'Ġ�>��}��(�1ы���˦�茟�ߞc���AI˻~^O�Nn���^������RR��5���t�'���2�r�\j�(�kgmE�[���q�O���zR~q	m?O�|���!�;�i��C�f9�
�o}h�^ۗ�tmO��~�Ҳ����}'jt�d䅻���L=})��C�]�l��ƚ�KJ)���2��lJ:E']��5δE%ʻ7��;�X�NI�!	�Q6�n׊ZH��y���F/%��/]/��'�s��B_��	;+K��ҋ�����#D�H�iN��c+��?�����ɏ��~�1���ZZ:����/-�s�ʘ$ݘo�B�ú����v��YkOW�y6A$v1�}�6^�T"��H
õ�*p��ށ�ukO��B�|)-�6�\��F�q�����?$����W�R�ʥ�%���JK)#��Rs�)�RE^H�mZ�Ck����r�jB�z8�ؐa���a�\�"���QL�0z�:#������B����q�S���������=�����>�g\આ籏�������o111�5�G��PqİF�\n�$�&���Y���#Dj�݇�ܰ�.�a"$+�tu*��s)�T�X�w�E֚Z{���	Q����)�����Ax�R�ؔ�^��ӆ.;����kv	��RJ.k�W��q��y��/��o� ����n��@3��o�u��ό�M��#+��G?��}��X�e�Cowzql?!d���.�>C�Ey���C��~��},��f�4yS#����Qb��e�D'Y,@��F����t� 8��Lˢb��6��ցޛQ>֙%]��� ��K���P;���H����iBh���9�� �~yB�g@8Y[Vn��e�s�vК�g�Q�>����8�|����ăk�o��靍���ݼ�t��Gz�%��g���O>�(�	��XYnI}�\\�t�O|ڹLW2��heg���N�T���ё!�[������米�L�b�ӷuKzo�P���ex�5�V�M��nH2����4�]@�ߏh�M����O$����r�<1�'��*�51E� I滽�i���j�
��������b���ڣrgY5�3�¸Nmh�-#���O�Ҿ�+�fFK��߱�Z�g�T�+߽*<��1j�3��R�|��jF~��p_�����aFb&��x!�Q;�eu8�Q���h�E1+�%p������Ν;Gnm;R�Ļ����gȱM�>�}֋��3��'4v�lt��e�����Im,,b����������0��G����u�H ��w.}�Dڌ|y@:��Mh^�W�c����a4�?)�R21�aX�@�f��t������ z|XOZ����zg���|׻[ֳ��l ���Ή"fc�z�	!��mQ����	��}#���p���	��ʿ��]G�i���Hc;���o4�F!��d�H��2�L�v{�p�ڵ=��fI��5JA�t��x'�\��(N�H���2�EK�'��2ˊu�e��Y�e:�*sԕB�W�#]����~}V��yBŧ �Ypq�bCr�M垻���.����h��Sn8O�����c.���wO����f?+�͙V�?��~�X�%�8�~5o�Vq�pL�׸~4�WGzP���e��0�(
��q*�M��ni07Ѓ�͉+���\-?[�<�'�GP��-?c������P=:�;M��A��� �8r���L�ܖ�����c�	�YE��AGR(*>�dPQ��}�h�A<Q����DJ�l):b<�:���-���eQ+S#��Ll�ի��g$�sS���S�����'Sk��}2�)0q�RBZ�:�ˏ���p*��̙��z�~� _zdhQzJ	h-��{�=��҂�����/�O���kpYa�&y_�8��3J��:� � ��p-SL8�\����X��ws�N�^�}eס��su��Τ��F'�\%����lU�@�v�t^�	���߭NuJ�iCn�G��O_�֞nQ�9n�����RƎ��	WJ�鷦�e)V}}�@zxH�}���#�������!���'Mo/�Y�Y���8z}>g�h�z��|1-K��<\B"�e�~����ϲ�gI6�nLy4e�:�2ҕZ`�,�.]Ż����@��+,����½liT��S 6�M.�)�3з���`OW
��w�	?q9� ��y6���}�b�����%�o�O���Kߙ>�A���	\�~�c|��	��d�:�Mz�X��?�rP�.�H߇�k�R���6^n����4��մ%�"1�0#o�߁��}�E�����#C��q狫v��jB� o��/��O+����o���l��N�݃�$h��5��q�E��C1Ͷ��>�a4D}��l�h�6��rҩչHr�Ϣ�\�����L�)..���t���"K� ���([���z�����g��>��}27R�}�O�����`R[�pW+���aZQ�nf?���-)�����<R��S�	:~Y��Gk:��Җm�����ӗ��{}=����Nm��\Ey)9���~�M���*���HϏ�k(!��UG���kw��]F�`b�� eԿ�u�>�r�΂�v�}��	D�7d_�E�?����ڼ@L � ���Zn>�o�1���E-�sy�t}�6@ؐ�����4��v?��v��W'��kʂ�� qGx�����w�Vn��}�7����J�1,��;m�(���K��V8�up|>�5� �h��;i��X!�M_��r��-�D�<y_���7�Oz��������ā�����Sy�̔��n�kyeh�g~����{м�a�Ѭ�4�GG:\�θh�qZ�|K��Dֿ�?E>0C��kE�=]����(����^�����D�zpo����R�	b����2�z�X�_��?Cڷ�?�9����H�`�aF�����D��Q���D�/$��i�4Ni!�I��l�#���g��3�������C�#�퍑����}���N�o0����op!ĆD��lc릆�}�h+++!��ӆ�Ø��э�v-���/�u�U���$*Χ�Rm�L!���Ա�bH���8����RJ+(�܊	s5�X���Қ
mtT�e8��SS��>m�S�";�t��>�A�,�h�EZk��l�`���m�j|����)P�u{HNh�O�"BDY����~��Xd�B308W#(%!�J��rB�8�1A�D��rՙ<�qٰ�G������+,2E���F���zw2,�c!�M����BL�&���4[Ƌ�:�k�N:v9�e3�w��~�'�onH��LJ�p{�`�p��_g!���Wd�7(�b�x�)��]ڊ�w���q��NW2����p?z�0�� ��ڇfҴ�V(R�?�G�X` X�xk�>�k�/H׬���42$H\߰�2��?o'á�ѥ��sK/!&B�H�ȡ�S��[Q�[��O�� L�{ߗ;���?��2mfH��V��<�T"G��|�^��s����y}�����v6tG��bñ�=*�~�<I�|~ʚQ���	3��Y�z�i��;�y҃�#(�ߛ��r�q�6�	X_��Z���E�6-e'컥{�!B=�u��~=pJ��!�G_{�m�x�]1N��ǯN(\|p�g� �ߒ����y�Kk�L��a�K�h!^�S����Ʋ{���b�5�E{��1�)^\�S$+<3����+��.�����&�/�b�58h�O��j���8�AꗍY�L$6%,�cFs�+/D}%%%,�c#������Hk�����{	78s%_Q�;33���N��.���h�}F�J�sB���7��hc<�O���b�?�v����}x}�c��}��?���wue������fPJv��>X�w�?���o��ū��	�	)�տ|�e� hDɅ}q��G)�ڔFP(ɌE�u3�݂����$_e�j�.��%������kv�^�gd� D\���Қ�4�{���Ey���-ѳ�%J����ֆ�o�$�ӳ�\�(��ռ��a�n8!A�'��Ձ�� b���>t�����=9���y��B�j
�� �Xx�H!�-}�
�	���Qp.{t�Z/�,�k2��,���W�GJe�Q��W���m�����c�_�����牑'8�����?w��nı��K��ώ�CO��M;�Ƌ��k��y�k��iN�'h�����;�|�,�� H�� �1�±��W�v܋�@h��?&�d?�Q����-��p��=�}!�[)�'��� ��~�CC"H+<=���j��#������-�XFK}���[���f1��f�#޷�6����0�˕t$��15�����:�~���Q�����^�a�XI/OJ׭祾DS��m8cC���.�� G�����{?SV~!5,�cFS��rs�5(�2���o�l�u��Ud�a���N�f6�>�}bB	l��H��~C��A���m�#\ກ.K�biўc�/'�I"���@sNώ4Oڰ���E,�`{o�0Z�Xp�v���<����ݿ�X���w����P�;�Z�u���$��wE���~b�+�ֳ�B~����k�ff~!�LL��93�D� 69��T#��.(�۾_#J���&��?�N3�^)�)�V��s(��x�`
�~�s	�~��"L����#�l�$k+K�w@W��G;��+�ۿ��^�t��
KJ���5���C�B����%e�{���B}=�X��>���C2n�!�
��p.aga��f_~�̉�������sWkN�D2�1.v�#��a\\�����8!f���n��`܈$�^Ac��p?��!�0���M~5o��$��l�pQ�/\�Q�C�:j#�3cv�/���0�A��]����Rl�Қ6	5�~W@��*\�1G�;*�4,�cF3@�gmm-�����YM��9�QI�V�0�0j������u?6����7� %�փڝ"/$���D�޼"����Kp3{m��D�p��w����tZz(�~�b��pQ�1n�70��Ss �,<�"\�Ԅ���#��}�!�����Y@!?���:�F�LkK�J��4e��T�b����D�E%tW�."�~ŽSi�7����h[.��lPOB���3�On5vDr���pb�gWn�?����g��e�[��L�,ݬ(Qf}q�8.1R̜�ӘcF%�=���"�+%���kM�ڎn�F��p�\E���I����8C�c5���t�_�Й_�ϒcõ�ڔ�[����
��㱇����Q��a�ajˌn*�� O(\�j#�W�����&�\ '���YK��l�}l9(�BՐ���.�M��3������g�c~��`�9h���aM`aa!D}�(�E�a�a��?p�0�lTq�����Չi��XZ|0��\�&Qc[/7Q6�Q��ⅳH�B!��b�;ta}폣��u{��QMh-^F�ħg	��aZ�Ih\�Ή������TM�� k��[�DsC�+]�k[GN�U� 0�����Z�U܏Pb�����v5m��ir���ZZ���_���T�t5;O|'З�Z�w� ����Uܗ�]8����,�a�	zq�N�ȨVJ*�xm�=��u�;{�ڝ�<�u
IAؐ04+��p+�;w��>b;�xM�c5p-'O�z�������a���k�����'3_~���A�8�����>`����~��$?Qr�Q����[�cfC�+�sG�\Iʺ����~f�Q��������[F�\Ij�q悾���5���߷Т=;��zu��n�W��16F�c��16�����62$��R�Vs�;�ck��O�M��ͮ#���nbNgv�P���CR�7���Ϸ6���("��"/\i�[��t�a�F�w!�C�ݢ��3Z�a�a�1����@z��.~p?K��#�R��Q_6�Sӊ#��$j]K54��'wmG�׏�x]_|����p�2�-Z�%����}�}^���%JfS�Q�3�ӕޘ4��[��ޥ���",�����\�[�Ҳip�	0�����wPAI	-�S��.��$���j�;t���G��1��[ou5G�}��p/�=*�>�e��{�����b� ��zv���ڀ=��Ƶ�\�ҳ�33�+_L���� �4?'�\��^A��l�L�-�C��;��gm�K�G��C���Z�\�+mSs��U��5<$���RM.�w��^�/�D<���G�y�2O-����_9^�qLc�-�{,A�cC�j�����J�P�#^�u�*�$�����!�>�5\�q0_9wџ�ԜO����mZ���a�1�K��������i�P�a�a����N�dk--��
�� 2��,�4Ʈvp�B�{u4L�A����ؾt��kUQ�S/j|c�,��1X�]�ʆ���=����'��������hԥdzy�.E�:���P6#.5�u�Lr�D�3����Qx�7��y?m��X��v�M�Җ�ot���F���z��}���8�x���<����p����յ����D��	q�]�i����j*�T���su2����^bk��m@Ojv�e{��#?��Aύ�+%��*���\�7��(7Yb~ώb���u��cn��Q�K%'�0�A{��}π��4?�M��A�~�s"������Bť�b,xπpန(]�1�D��I�K�+�r�c��Ù��>.{���ʅ�'Ή� ;+K��	4��Dl�����[�d�γ�7��X����q$>��(��~���.-�{4Ak�jkqD�I�!ss1v$F�%�	������Ԯ����FT���4�:c�.%�}A�s,nX��0�*�C��
E�ݲ2^g�aF~8��Н};�?�uB���/�eQ1���t������G�/v[�^tk�0�S:�p}��M��S�N�fP:����N_WG�3:��o��g8P�g�>Zr��q���xmq9#��Z��>�e�X��׺%-�{�(y!��J����lQ��z��.���']����-�}zpM�����r��3v��+p�*�`b㮳	�=&��8�Ҭu�-�Z�[X$��'��Dm����pބ8b.8{Ն�F��K2R��ĸ�T}2k�pȂ�����]�Y��5u�������,8�U��1M2#�aԁ�k6;�5?���Bq�^C����b��c����i�����o�t�B���g��K�!+
hA3����n;sI�LˍeQ����^Ծ�����6ێ�񔒕+�M�fM��V���z�Q���{���8���-!#��~W��7�9�{�ZA?}h84u��T}?}'S}]�|\�Ԝd��q�>��$��~�<��b�@f��0�K�p�ק������u��I�c.�������(��f��>�aT�N�#KKK!�����һ�0��,<~3l%�zs`���t�O�E	45OkL��	.v�R�j"�A�hh�@��T0��֔�b�p��ㇵ��v)��/�~ �).)�Of��l .��B��Vb����/�Ҳ��A�0,��Z��۝�� �:��]�������aB����nu����-,�w�5��+�%��0)������Ld\ӔSjL���.\J����'�21g�p��rTW����#�}��Nm��91H3�����潿l���M.� �=[���"8E�� e��(��`^���LfQ1=��v�#Xd�����g��Elp���A�0,̛bj�v�b�C��H���,@��j�� ��J�.y�o/�/�"M���%�3�xa�
p�n��q�r���ji���gh��bLW_*_�����=FyS�i��$-��3�zӼ�;���#"����8K��!�	��nIc�Z7y�������f��>�aT�ޥ����rrrإ�a�Zq�j&�^�Kd���@)+���0Mɉ�L��tg-�g	1�Y���9�਀n��K�t�B"]L��1��GF?����	rd�b��I�o`-��`cMS��ei�	�$�d��#gh�Y��W�/�X�"^ĭ_�h�(����#�$�8a�hcMJ����*+^F�Y�sQ���qO�pJ�f�1���I�(>�E{ϗ�����'��p�ؔFrV� ������q���Ծ�}�J�J���"A��,Jp��^��缥{�CatR�b˶b�����B�ҕ�:�x#q���p*N��ֆ��%��9�W�؇���+�W.�a�ȁ��4�ӥ����"�I?�u���g��U;�c0������14�K[�����Ab���m�>���6N܃�c���x|�!V4�ЧI����� �5���
��Zq���q?���}_%�3���uC�ZK�b�&gО�U�熎#p~/���E��qS�3ƕ��bd��<���]-�=쪭R�fo[��ɯ��MK�"~~i|1�jJ�@�ݦ쫰��a�A\� 䃠������LH\��%��#h���\Xc̃r<��>N��0�0��M��uZA�圞����~B�7�G�,�Erk�������={���o��Dj�[�7��og�ѡ���� e�0ٛS��id���"&Q���Yr(���bn��PSP(�-V6�B\��Lc�{�����g����m��;x1�~���[�t@�����?wR�����{�	�
\��-��;&��

).5�b���޸˲p�
��ش��vY�Z��8����7@	:���/W4�g�%jił\[�JUN�j�(�G��+���<�r�� I�ޱÊ�X��m���y\mF�@P;E�Nc����U��`�SUІ�o�~��P�������V;+��r.n���&viK��Z��n�v"�����(J�a<�y\{��ҵz���]Z�g��V�<�����mk�LӒ��o�w��(�;�㕞��KD+�z��/��s	Կ���cz��hj*�ňzG˦��}�(}�]l���TP�tO�a�a�����~B4��{~��V"�ȼ��yZ��Q䙑������рZN�����<P��J�:q[bf��p�q�	:{5�� �4Q���Q��diq���9(1��7E_P��2Ė��qi�ūBd�o8%��O@`��qYSF��mD�8�P�?[)s��%�^^����w�bςb�c8|!q��'gR���h�Ԝ<���Iؔ�rV=#6�a�aԇq�#�7P��J5�p��<Q��!�>���ݴ��Yb��p�m����4e ��QzA��
��.�0�0��Ҧwk/��Q�c�n�nmb�Ȋ��N��,��щ-[A.vzqBCڵ�Tj.[b.
q۟�ΒZ�S�s#�k�����ȓ�Z�b�a�iL�V��a�a�a�i1Iׄk�{�+z� �f�B�O���a�)�Å��ׅ�h�_���i�yOE�릀�}�(}�]�1�0�T� �?��g��7�<��J�:O;��!A���v(FlZ�6⶟��e��@un�(A ��{�����P��ۛ�7����PBf^��¡��ee���]�[Hq��ϑ'��e�^˵�=��=�C|��hj�t�sY3�V7]�~�j�p?2�۳���>��Nm�|����h��(�=�k;��-�C�ͩ���{ht�`Q5���'�s���w��JM~q	E6Rŀ���>�ad���.��%wY��0�0�	�p�;�0��˶ӗ��/�C��l�}�^�97!n�Y��p�<��b�DOIim��@?E���N�5�m3Ls����4ʨ7�:85�=�ٯ�X� +���Q"���J)Zc��=��w�
ڳ9L���ʎ��˚����q���*�W�����n���_��땢Qc���p�����k#��1����R��B^N��𐈛����8�#C{~�q�	�+*����}���3��S^^)��0�0�)<*l�ZL���v�4/�,=}�"J�bB�)�M	�Ջ�Τ�Ӳ�r㥴,�2(�зuK������;#E6�P[�8�qs�c��Am��{|�6�}W�5������U_��|.k>��ƒ�Ϥf8^�WMp��W1BxŔ�/�{3@�Ýn �����и���Zn>55o����vmO֖Bط1��M�w������S'{�sna}�� 5%,�cF�E|�ǒ���1��1�0��+�3���PCp����y�V C�&�P(W.g���_�����I�H}s��@Y��MXn����颔vrV.��WJ�̩�������Aݪ����bzg�~RZ����+��o-��e�/^�$�a~�tk�0��=�0�kLBz�h7��i�$����+DLPWq�~�4�&]#5S�㫦�A���}��V��c||�t.��9Ә���ʛ<� ���Z�<e������Jk�i����ʨ�~dL��*����׫ʨ���)FS�Vi��vS?��_7ж���@��m~���y��b��Fcp�j����g�.�dkC������k���H��4\�P��?�o�u �1��@�g,��cii)���a�Q=zqL� �}���5��O�@4������ÿm"9���9�i���Bz�ͤ%��n)Dn���o�Ֆǆ��/w��³�����L�K�C��7Q>(_�y0q;-�=��ّ����zF^�;y^����qbRW	�5�����㭌�UK�H�	�p�p�H63�q���7&���GU���U����H�l{���w]�m���b\��\	���Uoe8^�ū��JJ�)'����e]�Ȧ��V�/wN"g�0��Yb>��/&QjNe�H�yj��D��-Du@���#i�Ԗ��ujK��-�\�KaȀҾ����f<��˶�Ģ���}�b��t&��Q���|��=��Pb�>�#�0�0���q6A,6��r�!A�9����|� �<OJ��ʒ
j(�9�c0=7��A��0r`Z���qk����?���ǖV>���|r��F�'�nrfj����E%�SP$�@\��?��o�b�C��)ĨL������z��R�hǦx���}5����B���:�1Jȼ����������P������bD�֦��� ���^Eƫ�s��^]�[\_��&�{�<8C,�U�G���z�CK�TZ�^iK�ݗ�ڿ2��G�h�zeea!�@�_U��^)-�֝<G�'�h��c7�߀xo臋�9�hH�V�9���VH�����5��@B2�3�Ֆ�>b�	�]�\���}��LF,�c�_�����R}��Ղ�i�ƛ��A��n|�0�hd�틻,2�>�1��,\&��-ȟx{�Q~
ْ9CrDw�Jsz���3�E��O���[�ӥ�,�{�����}`bIO��Āyk�|��V�'��S:>v��)�UT}% ��;XZn>�O�����*,��L�!�(T:��vDV��Q2��D9�����!�t%��E�������`��F�j+^/��m_�Z\��ѷ��n[�������.��k���)�I:_�f��P2�U�H�*_�^?��!&�gFt?�NNS�GMq�Iq�H�"B�ϧSҨ@���}��f���Ԯ=��+>�:�d�_5���!����GM�i��7���e*7E_���b� �Ӆƅ��V���u��C����o�Bfc���m5�����W����.�2sT|?2Fk�9�r��@_�H��I����c���	tw!-���Y�v�i��1�?��"i羁�B���`g򽨈q@�~�~8�~��m�
	�ٯ��n�R�G�������IGR��#�6Jc�����>F1���
g7������2�0�0��嵻i݃3E驵����%��{�9e����aM��[[��{�������:I���4�K[���r:��J�zu��NB�o��Y��\R
(]���Q�޸+���--�	��7�Ǌ؍�K��z�sl�E{���1.���Hs����D/��/JT�rF6��ϝB�)w����t�rG2w��B���-H� �6�o���5mef�Al�k�};�r" :/O@ύ�+�Q���cg��Q��߹�X|Ջ8�����焐sۙK�'��a�C��9� ?Â�����P�x�*�=�����V���B�@/؃�����^��_����O��U�������sl��G�{4���7��4N:��o����۪F+�����Q�x{j��q�JI�����j�^�h욬�3]����otߩ5���eе�|R3H�su��"�j�!�kj�����>���$�e-,t"�s�X�m������ǿ���z�����Mi�:�a�a�a�	�{�2��=���~B0����\�9!k->-K8`9�ڐ��uiقF�ьn�7d���zɕ��5�� z��FrV��d�ws�w��Wg�Lx��{OA_|�;�ӽ�-�{�p�3�o�-��$��/b��XԗWT,���ʒޟ>\L4�qT�.� �����C������Z!|��Q��~DS9z;;�gۣHδ�r��(�Z_���NdmiQ뉬�Fo|c��,�x��)�}�u�.~���u"]d�c��$~?�;aR���ˇ�t��ҵخJ�!܃6�\�N�Y�J!�ߛ*�չ��!}\K�v���YE�UWjs|��=�/\���ڳ9����5v.�9���t���S��7�?�x#�8r����b�^���6q��{h�o��*�v��Z;��ڿ2���C#hR�&�� f� 0�	�]�"Z��;�3����zEJ��Ʈ��@�dlL�SZV&ܱ1���a�a�a��w6��PϏ�+J���[m���=��%l��&����Y쟽�N��Y%� [t�-���� "�����6+rЏL�����p9�v�1��O�`!
���ߕ��U�������t&%�m������AB��ߩC���DP��Hό,�a���ZjN�(���&pmD�yB�x*N�Γ@_>��ҫK�%�=��b���
�ڻ���lK���i�x��oJ�rKע\6�7��c��zQ���a=Ć�}��8-��i�(��y�U������Җ��KJdV�����������Z�W�|���e��RpW�M�P�������Ϙ/v���>(�Pz��Zا����ڹ����X�:�E��U�����Zc������ݝ��VX��0�0�0����(w '�Q��7�E�
\�>�E?�?qC	*9�����,x��*�� �׻�н����]N��_���y
kbP� Q�<�t��(���c�c�<zzd/!x�j�w
Q'�����	�����"�!AB��T��bE[�8q��V�����"��R����	dci)�Ϯ�Fr���̪��u���1��9�^��gEk-޺`\��ݹ=;�-��452�?�9�^�4�^_�W�g�{� JŨ��%�{w�UW\uEk߃Z۳9�p|�#��p�v��5�����x<�\��C��db�p��rr �����m5���#U��{߯i��x�ܞ�_���6�0j��}�0�0�0����I4��(��E��B�/G{�ǫk�yt*�틻,ܠ�,�ӣ�@���B����{I��7D*V�p����Q����A����������1���A��S����ד��)V�'�>��%���g,�3f�����P�p+�ß�I���~��B�X�s�ϵ��\��ޯ���(�b�=�@��9.\ˤ�6�[�R��P���7nδ�ީ�5��\��s��T:(w����UW��=��=�ÿ"^C�Cƫ�ҳ)��U8x[[Z��X��[�'���!���[�K��~���mU��s�-ޏ��;E3�ן�WT��+ՠ����6�0j��}�0�0�0���k�b3v{S*�N]�2;�RZ�a�p-]8�
&���KITjBu��U���Nh�<!�k��NJ�}w��XQ�!�D��]#�}�Z�	�>�N.�qbLOG{���E�+�g]�׺\�x:9M�]}�v�ٯE�m�:�oc���J.����!7'ש�ZY�啱�9u��XZr�E]R�}�w���B�xq����XZ����Ju�W���~�t��=����Yz��s��_$X�?�T��1[b/Ҁ��"1dz�7$Ȝ�r�z�R�V>�J6����N�^b�rF6��]�����e���́����W�׫��b��ő�W*mϵ�?+�z��F����a�a�a�i4�®�ZEF���哒��w>S�d�Ǥ̜jK��D0W�L	�K0�	�ju�M)/�l�ӑ����ﯹ��+��=}辁���o���p�A�V �J9�x�ⓨg�/�;�k��=}���s{��8�x�Uzn~[b.#?�x��	ɴ��tg����-^C9���s[lr-?+��j����u��� JƵ�>�UW�;�j�j۞c��ъ#�U���y���e�	��G�^�8P8}���nx��ȓ���;�t�������ː`$���֮WZCk�Z�W�������:o����x!`���z���WQ�&3��`a�0�0�0�ԓ�
�J(�B��W\Z��H^Q�x�N�'w�U�q�����Y��ݬ�惡�~�q!��3��?W�R�/�������\e}�����l�Mvg6�$��;$��"rA!X�U��r�V%VI��4�V@I��hZ�
R
�`�"+
��@�E�	���n��˜��I6n ���3g��y�I����>�y�s~��wbm�/���Sw�{��ba_)�^�����q���o;����_v���^ˮ�wד�/os��vx�mć-`�"�fOr�{�[�#gI]����S&�M.��c��g^��:���\�s��}�a;���5/�/�ي�q���ah^[Xp�����YS'mן�*h�l����
l_2Z/��ɒ�~#ͧ-Sj��O>�����{�'����_-�����E=I�����x\�{��ێ]e��.>w��?�U��t����͕}yPR�W;34���x1�;g��`L���} h��־�0�b~U�\�vׇg&lL\@a     {����������-Գ'.�n����;f��U�UZ_\��^�cJ��mE�;��ޒ�Dun������������8�t����_>��K/U]��zO��Ж���ӯ���ے��œ��{s���{�cG.w�O��+vآ��cSe�>��_~M_��|���Cqp���ݷ�����<s��m��\z�/>h0ח����:'�uҐ\���:d���5R���do�?�����'�vٟ����#oߺ���>D��>|�ݿ�w�;Uf�r�����ϐ�v�߮�_��UY��_?<�����KO{�4�>����+�������uڶ�e?(�&�����̵�M��jgl�����/����ھ6��*��h�Ǚ_1�:���և����    "b�,��#%���{����K�#��������^��?���/��g�Kq�՚u��������U��'����{�����3��?t�R�����Ŵ��O���=�k��uK��������yg?�lW���{�(�ٓ�ϯ�?=&�If�X9|��r�����wV\EƲ+��_~�T�ߗs��]��y�v��~ڻ�B���>ٚb!�yǾM~åvm!�~�F��OT̊@�=[dl/io������B������f%�~���Χ���y��b��^�)��Fʵ߃�{�c���]�+�}��wl�{�����}mQ�?lm����VXݜ�1���.����#yh���:I����v����T�	��´��#����?T�y�q;�6;�z�Z^{i��N���P��_1�a������a i(�    `=��r��i���{t21�y��C�|���g^�$��)�좰��,�WʊnϬ딿����O}H������R�ӓ�od/k��%{��R����եv퉶�}�x�;~��v��F�؂�{#K�{TN8xzqE���W��0j�zl����K��GW�7�j��7r��3�k��ھ;�Ƽ��6����ü/vy[%K���s[ v�n�מ�\|%����}ٞd���wʇ����i�?,3���@��>/��ò~c�$�k�k�:�������$�����Չ�l�]�_�8^�j�\�y]{� $�}    ����KZ�eWΊ��7t�4c�/Mk����sR=�J�e&�Qaߙy�L�_<�o//g���W���n��{E]{�T�G�����+��Ѯ�vR�M2�#��ǿC2�����׬� K������*r���}�� ｏ�?Yqy����C�ϑ�7d����g/���KK#���v{�+n�K3�C/=5#�;vՕ�}�yy腵R	�j�������H��}�{�.o0�}��ˌw�>۾�^ִik�U��睱��� ��i߆��U���
lߤ�˶p�ގ�oo9��/�kWﳫ�>w���ƾY�>�~��Xt�� ۦ���0�H�6^��8������θ�z4�����Ӱ7W�W?_�����	�\{� T2
�     "����|��dw=�|�撏�ǣ�����*��Y���*�S��aW;����Jb?���'�'߸��r��{˱�#S3d��q��n:{z���s��^.�F�W��Jv�wJ��4!Yy��Rۊ�6��O>�%g��/l���YS'�Ǐ:��R�-T�dCs͜2Q>dJB��Jj��L>�kW �7�"�<�v�$E���G�y��a�\�\����k�مף���_�k�����o���k}�4�    PF/�p��0m��߾��T����m�jvA���[WҰ����wk�y��Y����ʥ���������-�+�Ԯ~54�=�S�ݻ���7鿇�炟܊��~���~)�~`�����˾���+׸�/'u~�3.������0����*1\��@%��      �z������oF��P�۟x�xK���)�~�嵫����oI�Ǿ��:��x=J4^���?'y�����
�              �
�              �
�P1������GTU D����g��R������:           ��Q؇�a��@ycb�-           ����             ���             ���             ��� �0�l�u�])jV{Ƽb�Ԧ��;F7V�����x����N��'*������m"��           \��Y)FV��*c�+�'�Ft�=���R奴ƞsV1��?0��Y��33�g��AŢ� �&Pџ�{���6�5���j�[�R��`��MN	&iY          $��b�
c�F�ޮ����xK�k��ޥ��V����(����>  ��1&L��G<������QS�mw�7>��۷dn�غ1�`������y�          � �WD�c��뮾M���_��.\8�%�+�r�b�%�dMߦ��D��9Uk� 0B[W�*c
׽��ܳ�o���K�{7��<�}�EK���&Q3GEk          P��:#ڪ��\{Æ�����sr����-Ӹ����*�IQ#�%
�  &c��*޿����~J"_��a�Us_	���4-�2��c�AU&           ��yUE��������l*Ǐ�om^�]0���(�|�9+�
�  �-�/F��9}�evKt��=��l�EK�
W�].          OF|Q�w���b�z^�K�C�7�_
�2����^����S�Aa  �`��o<�l�U�Hm]�����%�������          @��&�}6���1���+���in���,ѽeGa  ;d��F��i��-g$�ϻ���K��~���?( 'g:�ؚh.^~[�^����W'?%�!GO�&�Sd���RN���=���ap-�� �*�F��*<q��ٌW�Y�x9��F�~���WQ��x�[�oD��*<��"w
�����*r��B��	sm�O����^���↛&�k�7�67���eEa_�3�HGG�$I6��t��]s���ſ�<�x�������ߍ;v��+
RUU%�f�k���s-�VH�r����?#��~������ Fa��N����Qmc���D�ڨ�Sʫ#¼�1��I�и�w<y#�x����X3QV�z��b�Ǝ`���Qm���*4��"�Z���QXƓ7r���������OW�b��x���\�2�
K-��u2^�f�y�'L�gs����cr����5,�
�qIßd��ӳݓ)�IDU-#~�[�*�}	�aC��]:555;-�EE��b_$H�tuu��L&S���b��
&W�I�ֵx�j�Hj�-re����}#�̰� ���z�&F���=Y��7�'+7��d�F�p���*)����+JfۗQm�bڷD?yC|�r#o�OVn�����0߈-�{�#�7�'+7��d�F�p���*(/U`b�\��gN�-j��T��r"��6�=�y溠U)ԉJ����Æ�ߣ� ����ߧMᴎֆ���mXT������}5?Rլ           Bg�S�@~Q��p]�7d�/y�����5������>  �X���Tո�:�>''	�����L����_�*�          �Y]��n\��'I�ܢy?�kn��/zW����,
�P1
�5R3Ft�8�B_o�祂W���M.���.�k��JY�쀗>=����A����d�?,j�`�          @�c^т9u����ڰ���Mmg��rQ��JnE}�hT���ϐ��Ӆ���Qn}�@Ƽ*���M-�*	�k��7Ӵ��U���	          �d�Ȇ�I���>�I����g��><�7�x�TvR�gQ؇
�BQ��
^ ����ښ���˷���ls�;��_          @��~��u��p����6��CT�	FoE}�}  g�/�[�G�j:���t���           �Q3"�s��$��uW����#��	��n��,
�  ��;_�q��d�TӢO��~LT'          `�C����\;�_Z�1����f#7��>�¾
� 2}�tI���*�0��#��Ζ�/f��/~G �D�	�}��+�K�ͥB�xq/���J�=C��
yGǵ��1��X!��7^�;:���c�ϱB��!o��wt�/�7��H_A���B7��ښ��4�_<��`d�Y�gQؗ �ƍ �󯹖���Q��y��4-�d0�~� @	��/�6m������S�.)�B�d%o�H6�탥��?�3Ǎ-��k�)%m_���8��;e�Ԓ���Ul�1^�&����;z�76_m�?ǀ�x5j���5�W���y�#�����Flx̟G�P`�QQTZ��?%���v\��x~��8F0<#(�(� 8Ƭ��v.��Q��^|��`��\ ��كRUUc���v�a�}�I:����ޒn7��������{�}�+`���4�yKݾ�?�mVW��Uq��A�0�7��o�9��m_{��j���W.�k�����ui�u�}���1}=��R������t��4�����'���b�*3�^�\�;ձ��a�q�T�?�J:�|������&.[��7K����+Q)ݥf�j�E}'�+H0P~���	sS�{㬣o)�vٷ �V�f�+���G?*PnQ�o���7� (�8���e���E��ГVa������fa�Sq�Ѓfa���;X�����}-ƫ�z���Z��-/�oi���_�+����R��3T��\6�W�4�Uٸ8^�����e���K3߈=5�u�.�����>�mj�5���-ع=(���*Ț5k�
Pwf��F�{�w N[�q����y*�}�OO (��|R4�"�Aq(���� 7۷��y�8h��7����Qe��^��k���U���l�i��E;�����I��w��v�}]�f�*�^�\���둵���7N��F��Ǝ����7��x��ϲ=F�f{X�g�� �a�kr��To����t���6�� @	��`C�'q��X�<y]k��<��(���N9�2^E�y]��e|O����2>�.M��RKӟ#C��ӼE��_����]1��*q��u�����;��g�7��>�� ��.�=�����*Ba��+���rQ��X��y]k_��ż���3�U�(�Ny���w*�9�o���92���Ѿ�9|�N���#��o���Fd��7bňl�PS}]^0����x�mg�E}�}  '���9���t���_��mu0՚) PbQl�CE��2���Z��7,��-�'��£�E.���J��e|��9<�/�Fy��v�����aQ��K3߈�y��9�_#�6���y������((IQ�Ea �	��/�!c��`~��Dq�AcTDa�W-�7��׵�%o���|�JO)�+�t����[>�����o鑷|��7-M.9�O����a�)�[6�-=e��[�1�v@�jۍ��K�u%*�(� $�1O�jzT�c��L.�" {��P�(}}��lƌ}cu���,���������O���a�/y�˵�7�xUR�gD)�xUR�y�-+���eE.���u�oiMg�-+�򦃼�о��xU^i�ee�y����"�7�=s��ۅ}%,�(� $��_�N��?��x����C֭[ʶ큆�y��׋��Ǽa��i�%n�[:���xUv��g����~��P���l���a����;�����kO<��U�L��x�h�6^����4����k���W�3���P�;��t�꺪qU������A��Y� ψY!�5�+��(�}          �#*�
vɞ�WQ�
�B(�(� $����~��`�L0	U��	          `{F����'�5�5���T�gQ� H4#�����y�.Uyރ�/          �72+�[�s��II߃�T�3B,�(� $�������澒ij˩jV           �է�����R�iI���J҅\�gQ� H6�U�a	&W�wG	          `5f�`Ԩ���ջ$�"(�(� $�Ê}�et�(�}          0�����"HMna_DE}�} �D�|]+&�b���          �m�x/
�ň��س��Y� ͤ]�a	&X]��`         �2�s�y�����L�E}�} �D��c�5LFma�          ����[0,�<�\��>��> @��}&X��?e�ďN          ��3�e�+q��T�gQ� H��*�$�ф}r          �=QƢ>��> @���F0,�J�          �P}�~�`X|�j�$\���E}�} �D�R���S+\�          ��y)
��IE2R�bP�gQ� H4`�5l��	          ��z\)n�Le���IQ�Ea  �|��aQ��X�          ����+5�_Şw�QQ�Ea  �Te�`x����          �2����eDfV�Y��Y� ��&X�T�,          �
��Ǩh{�-(â>��> @�ӆ��5�q��hF           �QU�;��K����F*IL��,
�  ��Fߖ�ⲉ�+?�)ة/��
��          D�V3�}����;U(�	u�9�E}�} �dS��}���;L�N          �����I��[;��승
ő�,
�  Г�¾ݙ-          ��P{N�¾]2��*�*��Ϣ� � ==�R/ءL��C��C B��r���~����Ǎ'qs�!�H�Pe�q�k����
�}���%N\����Z�q�We����۾|�p��l?��y���e�q����L�Ҋc^ƫ�GF������t�y�[V.���xU2�h_aTN+~5�7��o=<�J�UHQ�Ea  �T�mn=�kq�o�^�\��؃'N����P�'��������ky-��fy�C�CA��sl�r�������a��1�*�|��\�G>�|�\�Uy�y˃��<�[�����Q��.Zz�����Rz��]�Y� ��IqAaߛ�~n�N@ �Ԣ:�be2��lp-�e�}��о�#ox�[.�W�Q��А7z�y�G��d�oDN�ϡ!o���F����0��%�`�yg
��Ĩ�%��Y�
+�(� ����dn{�,��l3���=���`��� àrl o��򆏼�q-�k��:�F���#ot�>��Q�s��򆏼�!o��o�9{��4�]8g�`�l㒓��$�*��Ϣ� ����1�ɜȵ�m
�M�����T����q����!o���ϵ��Q�sd�>�F���#ot�o�O�ϑ!o��򆏼�a��cA�d7vm�t�p���<�/qU�E}�}  �\"\'2��4��U�|X ���y�aP��=򆇼�#ox\���?G���!o���F��Fx��9򆇼�#ox�=�;c.��������z�sz�k%v*��Ϣ� ���j�?�%r�@RF�̭<���A�AQl o�����[>�-=��F��eC��#o�����[>�7JO��eC��#o�����[>�7�,h�ٮI��D��1�eǪ�
/�(� 8��t���?|���G�mnW0�9+��+ �)N�y����G��!o���t\���?�yK���7�������Vڷ�ȋ=��We��[:�-?���!o�1�x3��>�͛�-��[�in;Z�����	(�(� ��.M}1�_ �Z���n���mAJ �<ϋ�A�A�`C.�+�6�a��&M�$�lV�&��qn_{�����d���c��)�ƫ�����r*�k��a�Wq���W��g)�Ul0^a�*�}]�r���}cc�}��y�#�񪒩Ⱦ}�.~Q\u��)�W���U�R�gQ� p��%����uU�*qP�{��/�8�I�R�S���������׵��y큩��ω�b�J4���5)_�ț\�M6�&[��F���i�?'y�͵���Wɖb�Qa��n~ۍ5�NT��+�wJ�$��Ϣ� � ��Vκy��rvAR������\�/�2�H���p�T^�7�
��D+оH��o��7�țl�ER�/$y�����D#/bK%m|�V.��D�vN鯻c������:휰�>��> ��T����.ȉ|Y\q�5UFzn�O          �����|E^d��bn�X-�M�R+q���>��> ���\�ij{ ��p�8 �P~=�Y/          ��P5M٦�s-����cLk��H����Y� ܥ��5MKN�n��R����|��A�/          ���Q�^����\K�c�`��%sD�?J\$��Ϣ� ືx��=��t~�Ꮢ@��K>d���P�          %��sW�Em't]���$P]S�������	/�(� 8OUg̏3��Oʷ6wH���o}����AH^�          ,�S���1a^ۉ�4�I$ۼd�1�!S�Y�� @���x�x�'6-:��e��� ['W�Uu�           ¥rh*-�����Ԥ��gW���ܤ��$)�(� ��/H����KO�l���T�LS�9b�u��j�           "���/d��Oϵ�?&,۴�SF̿i\j�*���K  &�I�4_
��6�������4gݜ���K����6�           �6ը�/����\K�-Ri.��*S�s��i��p��Ϣ� �7R���q0�Z�뮞/���
0�yٔ�y�� ��� 0Z'L���u樶qr�C���Kn��KV�L�r:%�!GO�&�Sd���^m}vо�Ԑ7��]�]E�H1^�'y+�ƚ��7f3^�f9�U�\����[;�_Em6�Uhne�1"��o0^�g9�U�Na~�[�_En6�Uh�7	T4|�9��v}�)�y���G*�ĦE���sS��x��KE}�}  ��,����|�����ζ�'%Ʋ�m+����Ǟ* #��'o��'7�xsŊ�mW�ɛT�M6�+$�
ƫDsm�r-�k�V0^%�k��k��m�U����*�V0^�R������3K?�o���ĖѺ���}і�t��� �]Qy��~�mj[�N�^���K�$F2��V#K��          @������6��� M�-�_��mZ:ӓ�o��b��>  vG����/��h���|�~G�����G�вO:��Wc��lc          _*^�弔I��mn�Ƙ��5�]�]�)[�z���KD�~�*A�P� �0����[�*s�6�-J{���
~['V��~�q          ��S������S���݌I-�r��(�����zF.5��Xe�?� 0B�:-�k(��<��~{0Ź~CMǝ�p�@�7�qqu�����|1r��          P�T'�ȿh�Y�������Ԉ�K��=a<]���&J�Yb��"�x{����FaJN�f߰:' hqż�Lp�vM|U����VxU��ί7�q���`��ݔ=B
���<�����t�z�s
           )T�_�0�wF�ѶLS�}�fE��������ow��1u�&�����̖��w/���z�Y}q�}(9��n�� p������D�y��J������+U�j_�����1y#^W��F��5د�%5A�ϊ/ۘ�Ff�.sX�8;X�W��*          ��NT�3�g���=���s6�+ŘU*����2"�g�SF�
�֨�5��OR#�ՙbd�v�C���������<���1���r��lm���-��Q��R��)�l��L8������Y����          \�"u��c��cdH��}�F��f�!�=x���_�$/����w�~�Զ6O�	             ���1�!*����            �-�HN���0�h�C�,             0�<&����0b�S�f            �=f�����P؇P�I�����Q�j            �=`��bݲ��1�!믺�+���?�ÿ             ���q�}���?ԣ�            ��#SUշ��(�Ch��we��U�#             FB�՝_��Q؇P�1����U�             ��1fӀ﷈�(�C�r�?�4��P��             ���MmMk�Q�!t�x_��<�"�             �`D���v:�Z�EaB��2oe�qI�x��             ;c�f�x��}�0
��|�k2�mǩ�             ���ɧs��=.������q�g2��ͪʙ             C�8���F�}��-g2����K�T��             �J}F�9�ҰHPDa"�Rks�,X��l��o�@             �˘ͪ�\K���P؇�-\8��S�����Y��5            �-F�ѿ۰��1�v(�C�t-��~R��M]!��	             �~1r����K�-��[�&���:Z�_���6�}ψ^�*'	            �2�F�z�W�[��v��>�B�����L�ң��?)*��            PٌyʨސN��ߨI�[�!V�ms	��곛�G��lDߡb�{y��f            @|�/9��c�S����>,E����������z��    IEND�B`�PK
     �9s[Ìs�    /   images/01119c27-1bad-421a-afe4-dfb48490a906.png�PNG

   IHDR   d   1   ,�   	pHYs  \F  \F�CA  �IDATx��|	�$�Y�u�]WwW�=�=�3#i4�[��e+�����Ƭ/XL�a���B`vp�^0�k������XcidI#�Gs�1}VwWWWu�w&��2������z�TV��|��?�����;Z�/|���N�tc؀M���5-Ð����j,Z�Av��-��.?t��/�K���8�q�>v�쓱Z�c����5�����3��곎�����z�v,�0:Ͽ���n�5�
k̪���<�E�Z���-}q�e_n4�������÷*���b����p�c!��v4t�Mx�XA_ȏ�l�ZCM�j'e{s���\���/��W˭��B���/B�Z��`w8Q���J_>�?�F��q�ܨ�����P��<^?�͆0T���E%����a��Ɓ�ga�Oӛ0($d�0�f��h���vh�\]z8��.}M�g��*� fG�.s�?_~�ݹ�:!�ނfwt�3���G�G�4�38��5l�F��������Ş_��_H/-<�s�[8�z�\�k��ƻ�?79|�]s�s|�+1D����'�S\��M���F�Q�u����5O˖�T�Γ�l����4C�X�����!T�i�e">���U�#3;��� r�*�C!l$��߿ٹ9D	�J%��6�f����Z�<�����'p��E���3E�p8���yLLL`rr���(
h�8�==����A雙�B`x���J���^<��0+��E�h��ge~������8�t:�J�0::��7&����|A�G�J��������(xB�)�?�����j5$}��� �o8�t��B�G���~�ͭX�
JCL�D;8y��-�=���L���\���w�7~�M��;�**�3 :�u�v�!�7rk-]ݏ���ڰ(}>��H_[W��7v;��.e��n�k�&,�4{��J)�!2�5��g�1,��x�!-K��Y[�Q׹�����m2��DXb����[Z甾%���K�X�}GP�Lc�>�cQ�n�
�gX� �����?��ba>㫕~Q��w�&O�w@b�t5�x��Wd�b�'��FSm�V%%��TJ��|���kS(y��S@S�p��)�#�=�B@�K՗�� ��e��h�L��BU�M������8c�0&ײ���U�h�<��G����/aT�Sr�)c��v�Ŵ�uazmC�@V��y�\9���h�TAB�o�V�^,)���3MQ��L���������_mZ���0�ޖ��@4������c�` k�u����V�#�ׇ���p�ʁ[�doDT��v�CSV���[������|
��S��\@"��QG1G��ƚHN4�n1W����}�Z���y\���qKo�I�a4�z�*ĵ�WL�KKk���F�eq�M0��)-�e��f�.��&�U'����9aT�e
BE�p����H�C�����s8��$�_�`D�Q��!Z���ǔ%��9�u�QJA��pF�x�P/^^^�W��)��g� �4���3H� ��_��f3��5"���S�6ӱ�	�@m���M�{���dM��r��L��DЅQ3�
Ы��Qj�@�E#S��$Z��]��<�*P����9ݵbY�a]��3a�ߨ�j���zS�Hk�\U�E��0��y�\N%����������?ǒ9�Q�m�9�zއr�<ޏ~��c+�X��F�D�E��E8EZ|�1�Q=s������u|��Ś'��[���z<��dʺ��b�a� !��5!a({ɀ�� �t�.�r��coԇE2�0}ۅՌ�.��-�Wkj����E�Ma���i.�v�w���1m�5�Y9�����J��<�<Ͱ�O�b�%���8�ܚ0���zՆ��$�(�� �|�o�W��T&r����P���f8e���/�������?6�ی{]�O^J�^?C8��l��`�9S:�Vj-3.�$C���{�Ȗ(r\�ms�����t
L��e! +� &�u��>�NŨV�V:mm��W}�������3K�ܤ
%�6�D��A���~���ʜ���ķR�tî��R���?$2��3T5�� R��S���p(��S߷��J��eٻ�ĸ�h���6`����/�3Ֆ&F`%y��e�$�q�%W���7�1�l�d�d	��ޒ�xb9�PdN�8�����c!WFYƦ��~Ś�g��3���iJ�Z��@��\S|м�3j-�GQ�#�c���C�������I_r��4���oX������#~�L�|�t�{��;'��&�A���!�kkO-�KL�'X��p9	n�<��!��&˄�n��Sb̸F���]��·�^����%ARvض��W��L���E��c�]���}ne�h����\��/5���>錀j��FA!1m��d��)3Z����!un�b7�o��c�5L�#tu�:��ǚvE�i[�O3��dM���s5|e�Kb�k`��nÍi�SE�X^1^�I:x�$������K�I�җ����c��:�t�M��7��P,�K�4R{�;`�1/w\?C��F�i4[�<�W6���`����A��E?!�ib�L�eݢ�$;�I�#����7:��{�V�.+��)&�rs�'�퀽���EK~Y��G_1�0����� �� 4�-�tzv�8�P�s��za�����ϡ��Ys^E����d��vR��e;�]��G�{��Ag�W�!LQx3�����Q�����:U��Q�8rНYa^��1�w��V��t��;;�Vi:~�~q΃���xj�pE���7���K��-2��
��hKc	��V_��g%A�@��Sp�J�ߢ���rw��r�1ix���s��/dU�=,afװ��|����/���l?�G��l]n��"�i0���S
�a��L��I�_�	\�{�JxP�_����s�W�dYΟ����Όn/�fU�Ū/���F������l�\���(EPu_�)ߖ-e��g�`�J鋻��i�����BA���K�1��
J�@�[�[��^׸�É�Պ���h�P�'o�nce�o��}��"g u��V���g��zO�|?��BX�ޥ]4#�6���i趽�sZ��D%�+Ҹ�!?*S�~z۽��}�J���:/��p_9Y`pR�C��7�	{�ư(���%�45�����A̷}�Ӧ,���H�6L��k|chǕ���!�����*81���f9���f�D�*V�:͕f���}oQ�p�hk0��ӄ�[��L�0�ef�RŲB[��w��gU�X,����aa��E��Gp0EIh3����L&� ��݊m乲�~�W �p�i+���0���ʉ�r\nV �H�C�)�h��?t��%��JC��L�8n ��l��*�Ŭ�6��p����!�[���~�|��423}��{��>?��|�1�u9�Ae]���!�w�"X+����������<[��Um���\�ن�-	:ͣv6"�+L�RW����Q:ն��N����0_�&V&qܞĥ�"�#T;��o@��~x(���pO��"dv��6� �<�_��	p�62�Q���XTqX8���^�53�*!�c�=��b9t���ﯮ�A�vxg`/M����Vwy����)�k��D��2�pV#�i�<�2g/ �o�D���=R��4�\RS�a^���e�ޜX��6���O�oH��)��k
�6���࣯W�I�����H?�m�!|���Ԛ[�Wmmػ^��+�j+��[����Ѵ�:^��U/�k7T��eg"A���Sj�r/�J�����e��؞�A��/�w�7�3�׶e{��%8��:�- ����^�)��X^�U&+[j�,��%�h'E��$��8�������n9���8\3�낽K��{wf{�`A�/.� b��U͐�j�NL/����*b�VA�R�q;�����c����G|J���3��X(톽��ӹ��Yx�2�1G&2�g��L%Xc�Q��EK6MU!+�������5��0���YC��Q�"�LcW�w)���zS��*f��B����m�m
�#�,��;/������X��4���kSKW���W{��d{u��-5n���ՍvL¸B�q��:�(�f:d��&�5�r�]�\D�_�X;�o��P�?sI��?��z���33�li�5�v��ỗ�ϋe�{k��C��.�E^��P�{f�Y��!�������W3��GY�'�k0=#���6��Z�a������#f���Q|��8�T%M��U�_�2���o�/��f:�Xo���;�wө�1�%fqk�CP`�9�ʪ��낽N��S&�?��0�!�O9��w�ϕ�X�q�o��JW*�Ğ�a��H"�_{���0�%<�͗��Ϟ�;�<����"7�O~㟞ŋ�)�|��?��验��0U���"�= c�H�����/�������ٝEKpO�s8��\�����a2�;�xk������qV�}v��t�ƛ-�l��KS5S"������N���z�&z����^���2���IUZzl������m��[��ǩ�e싄$�+�ҟ�ۅ�lq�]���؁Q8+.��7��r�ٹw��k*S@hW���^a�rVP��R*\����}4%�)�;���~'�t���Ԑ�m��C�QlT��ҙ)��G��W�����*N������Rk6�k���~o=6����V�c�Qe��BC�7�X"z�p�G��}[E�,�(�
��=�l�s��a��^��7	��(��i۳�j��lӜi�鲎��6lߧ�`㼉�g�凞<�r������?q����ןW�;�[�aY+�K�e�OC�$�OX.���?�iS�A��*��l�~�����*���I�}˕��������%��Å:
�*HnɠCn�h܉'jM�k�����(����3���|�\J��<V������G����w>�����&~�i������H�*{e���iG@L뎧�Y�h���x�
9��"V>�-tɪ�l\���px��,�!j�TMǲ�Ơ= �;l��z��	3Z���F4�ɧ������/���ˊp?��ĽB��X�B�q&�V�Yt�,��V�
��2!(`�)�xg��+"�d>�!��p�]���%Z��^�@�˔<��(�*�0dllO>�$���b��7T�����g$�L	�#��b�?֊L�הu���4j�Afe#U�f��|O�R�r���{s����7���"�E�i�茹܁�Ūz`�E�Ip6�D�&]�QK�|a�D���amm��_ɗ�\�¿#��"����:�Fc7��x<�_:}O�Z�s�������N����kw;�QɌz�$�8x@��xqj�� l.l���O3w`g/�c� p�{�w���3�f���X̠	b�A�8W�o��֮!�J�Ib�H�ZƠ��5�(�̥�E��S���l�g8�߭`/��6�|��d���f��ѽ0	��q���:�CG��w�"��l���$>��7�[�*x�ܩS����XtE����w!���/�O��	���Z=C�4e�z�k5��)ֲ������/*�׬�5�E�vE<�C��ү/�m�Mk��9����^.�]9�i����e��2.�a`���8q��Um5'�X^�vc��P���^�����p���R���:�u�>��x�A����O�|����g�����ދ���!\;����T�Φ��/�;k߱���wY�	�V�l�-[�~���r,")j�M�G�)��%m�-�^߾[1.1Q�Rޭ!.3E�y��e/����-��i�)��K��g��aUL�n$>W�����
���C����~��������R�jOp9�u|P:W�Bmif}j��U�3
�ejVu��A�y���`���̌	����W^��-������֓�����z����hTU�l�^M�+���_�\�`��;-aH�UE-4%z'#�80��#�6Q�d2�6.o��i��Qw;�9�ŝq��`}W���G�F�r|�_f�ͬ\�����!�� �e8�	E)�iA@�P@WK��ݶY�!s����?>�����RY�޿��)l���	:@�Dz�KD�(�Y���2�bA�5�D"��%|v���8�Mn�4s�&�e����o���!_(*)�Ő�{���g��F&�G]���t��;�sZ��^��H �Ŗ2>�)��P���Z>sE�`}�1�3͘C#��k3�)WI=���|A����JD����?�V�}�U�UG��������'.�L�F�.�Pr�ן0�vp>ݡ ����� �^J�"ªc��1��*C.�R��iZ%��!k�@7�@[q�./�|	T9hb��*H>�["���R.�q�P�9�����?	Glo=,w�р�n�3�cj�sY�����Oͮt�����ߌ��Q4�R���P�i�l�g�@ӷȸ���,��n�3zf������>/̯��@�*h��sp^��*zge&�Fs�_����@ȋd#��kߡ�n^�7H-��m��2 ��~���l���%ĮW�۴��R�M�f��SG���G�M�$����6������"Y5�2��d�N��Qo)���{���\n�� �K5�UjUo��+_���b&�2���2����!���Z�xĤi�EE1�>�ݒ1\n���[����u�� �Ί)��Z���|�ӥ>`iv��[�0��i�����pE����E6�K�^��>������b�!Lm�y2mCΟ?����TK��F(,��N��-��@��xI�d��a���I��l�Z����	Ֆ�@1�pf��a���W�^�k!A4ׄG��2�9�� �Q�Ii�H�G斻Ԅ?:�b OE���\!%�Z�ѱO��,6�����iҷ�x1+?�8�X�9J_f�4�A���~8�W]z�2琚??���!v��=5g�O�
2g/��K�e}�7�˹ϊ��va-:��gu��_�tB��#�|��E���.��O&oz�1��M�px|ΫL��|f�2�7��0��d���:*'����U5Aoo/f��q��AL�̨�y���%�>	�A��%�k)~�x%�N~�`P!��TJ}{�� �HR�U�.!/.-�o���%����f2j�nwaf]�	��>�^a�駠W+���o�\m~s�F�5?.��7X&ϟC�����BW|�G,j|H��5�i��!���hU;�E��q���Y�Fe��ڧ�j�����.xD]}bj��F4��H`�Ѹ��.�E��:؆�;{P	��:D�ꞁ,9<*�l�_��v�3�v�D�ކ�;��u�HBAvB���!��{M��?6`�+d��!�)S��B��M�}EM�����[�78��pWe9�u�ǅ�D:�"��v����v2-�ɦ��M)g������+��&�׬"���� ��ˑk�/����U;������}��b"Ygu�v�m����Ik=���l���s0�04�Lz������u�o˷�L�õ��(�dĄl�Bf��_  ���rF�    IEND�B`�PK
     �9s[�e�e�  �  /   images/3d0a314b-f708-4b2c-819f-35c414b123ec.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx���	���}����tH��$s�F��`.� �v�aBf'�O��ēd���`q��$��Ɍ3;;�M2�0�F�@�!��!�9BWKBg�������[���V���<�t!d�<���[����l    �8�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   � ��c����Je^�V�ӨՎ�4�����T�ޓN����I�j�S�F����T�֛�Z��ߓK�7��r#�*'�k��p�K!��6����!�5�H5��S�dv�����J��յ��5k� h �Fޙr��|�~b�RY��V��V*s2���T���fh�����K/����sJ�L�X�fG>2��J.����n)�ӯ׳ٗ�s漺�O�� ��	t :ֳ7��[ڿ��B�zN�Z=&W��k~����{饾�oI�ȥ��B�s.�Ri����E?�6m�|��C�|~o9�����R:�������G�ԉ_�B)  G�@�#<�|�	S��s2��ݥ�)�Ri~����
�z&��z=���<zBX�#o�������W*�����\������N?����7� 0a: m��U�Nɕ�Ww����/4?�޼��nE�V3�������3����/�x���7.�x`,��B���t��K���  ��@K[��O��;w~�06vy��؇zFFNȽ�ڔ����V�z�����~e����=wd����������7uw?|��5�  ���ʧ?]|��k�1~y��ة]O>yt�V��]�\�\.�9y��d����fK�]r�c����r_�����`��N��o\{��Ӫ��=�×�=��IS��hq���I��'%�Y!|��c.��������e�k.��W p�: �y��??::�dR���gt���M��j4�OT�tɶ�du=y��S[�;o�p_�����{�;�.���� Da�7����w㤑�kz^y�t���m�@+zk���k���֭���|�������}�-# ��#fݒ%��J�>>ytt��_<��G9������}�$�����f�%�l�2宝���X��b �@`�={㍽�={�?�;v�e�[�i�7����<�d��y��˞�鹧�����֬) �P�qw[���0ix����?�J9?��VS��]�<j�쯿r���4c��E��� ��t ���˗�0�R��i7.ΕJ�&�J��Oݳ�����~w�ԩ_ߗ��ɥk�n �: ����򱱏Oڿ���[����t�w)W,N�],^?+����K/�ށ�So9�C�J��� ڔ@�xbժ{GG�ɴ���J���T��y��?ع�7^���
�岻�� ��t ޗ�+V��>8����^;����*g���iɪ��t��^v�3{�L�O���_3 @�� �k�6�����h����[��M�L�z=��`���ƅn�3u������w Z�@��=��?�wh�fn���p�#�gx���㦭{����.^|gc֬�x�-��W��$����q���*?3mÆ�ɤ� �)��Ξ;:�����7�x�U�N����c{ �"�xG�\��ģ��~{���%ۊD.S.��ܹse}Ϟ��P�oߤI�w�w� �t ~��Wϟ28����L��~V�r��j���Mߵk�����o�N���B��y��=�������}v�o,M'@�K����v-n~]_��UWݿ���sW�y�  � �V��1wt��gnذ�� m&���l}��o�5/\s�ݛ���[v�}C ""�:س7�؛۹���6]+���r�{����O��=�d�-/M����׬� ��@�PO/]��_~���ccSt�\��7g۶_��ۻ��e���u� �� �ѥK�������l�z\��522縑��{�%�|j�QG}���o. �"�:D2 n��=�?}۶�B��
����{��/]qŷ��:���z��  L���W>�����/����w�~�z=3}׮�'>��ŋ������|: I����˗��>�Ŀ�Z,N�!ɖ�}s>5upp��U�~}ѝw> `t�6���ճg����Ӷl��a;;�'�##8f�����+�x�4oޯ�}�-# Ƒ@h3�t�9�7�j2�����^O�صkqyh�ѧ�/���s�W ���&Y�jἽ{��o��3pX�K���m���W.��cCs��+C� ��5n�)���O~f֦M��T�]�q��{�\4���o<�t��s��- �a$�Z�c+W����_��9CC�`Bd���l���.�l����i�wl pt�������͛?�qu�Sj֬L������k�;j�Z5��L޻������^���<wݺ�
 �>	t����fN��S6o>7��0:Z�_tQWH�R�^o4����|���ju`��ؽ����d��c�n��KW\q�L�_,~���x�:@y|ٲ��6l������ �Icd�����LɄt:��>=�m>��'���o(��P��7o�V7n�&�7�C����v]������U���{�x�:@x��?�޷��3�n�.�לq����@;������|�?���8p�Vk���b��zSatt�����s�\s�^xS�曽���"�"���ۺ���>:�8�o�V���?�ߛ�4)�=��QH���w�U7l�T_y�Ҍ����t����}�Ͽ���|k��z�=�� �	t��%���l��+�Z-`�����N��s�f����K�{��*�X���r��gO��z���	�ſ~rŊ����k� p:@���S���d�-�4lig���7FG멞�����$���睗	��U߽�V{��r��;re=W.��e�~�k�r�׾��  ?�@���Wϟ���e���B{�H�;��i���HϜ�i>�s\Еl��|���ꫯVB��9_��zz���׿z�e�=��Y3 �t��<�bŕ�l��Rir�	���/Xp����T*=~��|�?�Fm��J���M���r}۔�{?�56���?��_<��۟ �6:@$�[��Wfo��ϓ!S���֭�����*RٓO�'�ܞ=���ϗ*/�P	�jۗzat��y��~���K?���{� ��xp�={㍽}[����[�p��|�֨T�\nB��g���/��'w�E��K/�+�ח����L��u̶m������Щ]�YW���	t�#���L۸��CC�8����ع���?BoH��ܙgrg��OΪ��}�\{�J�no4R�v��Ć�:iݒ%?���� �p�<�r���7m��\�8=@$�C��@���Ϊw5�]�j���;8T�MC}���g�V����+n�t�����'���Ǘ-[~�֭�W�\���{��0KϚ�),[֛�S�|�;����_NV��M�����V���+~��k�
 t4�0��]����l��k���d�P�7B:=!����z��{�\PHΨW_x�ܨ�B;ɗJSl��W�W��7�֮�3 б�8�@�]s���ٺ����(�~B�ܨ��]KϞ�k�ԤI��G?ړ[��P~��R�����=w��-��;�����O���_�v�B>�{��O۾�� ��m�]��@�W��=�P~≱��/WB�H�뙣�o��/^u��S���_ t�(������Sz�o�J���	Z@2I=�uV!D,5}z��tio�3*�G�������Fj�Ν+_��)']z���6��"���߬\9u����CC��Z�-����O~2[}�����ط�-�v��]�ox��5/���p��5� @G� ���իg�߱���������H�18XKM��	� �Je.�g�;.Wy��R����a�ܔ�{�
a�+����'~�� @�� ���eˎ=f`����QZP2�=�*���L*w�]�Nȕ~�X}����	�N&��{ցg���go��cg�r�H ��	t���[˗/8n��/7�|V�u��)��CJM��)\w]_�7*�*6��Zz������ү�~��V}��;�� h[�0z���N�?0���^� -�>0���ɖ����|���c��|�����{8�F�GW����w��f �-	t����+>|��m�+�����޽���h=�ӓ-,�˥�_ܝ=��|�k_���ٲ��3<|�����z����Y�- �v:�a���U��ݶ�ϲ�6�܇�]�����3fd�����Շ�u���=z��>�߿��5kv ڊ@x��X���9[�~)[*M�F�۷W���.�"�9������7�l�JO�O6��|����.Z�fo �mt���[+V3o`��\�4%t�Tww�Q,6m��B����33]��d_r6���S�Po�r���s�<{�י��>:�{��s~������d����rg�](�}�H��7�2��;�y�F��H�q�v���_xaw��>v｣�Z��{���7޸����^���D:@� ���n�9k��;�FF����s��.�NM�t�<ra�Ҟ���<���z=4v��o�m�?&=o^���þ���X{�Jh1���'|0�/������׬) Z�@x����O��i���##�B�K�<������@+�]+V�6#=�J������@-�Ɓ~Pww���Sy��r��(�� �I���׳��y[�?�~͚�����]���{g|����cC�˞tR�Ќ�$���罹O�t7��x�#�x��CS߼�-j�t�����}�T*w晅��ٙ�u�FCC-�E=eϞ��J�Y��? �,�p�7ݔ����y��gK����W^ٓ]��g����>:��䒮�7�9hK��[���r���K�OM��	m,=gN���~�o���Zj���ݻ/�k����}���$��K�>�'3��]�X�Sr��/�I
��Z��Ї��{�ԫ����m*�V~�R��̛�͞yf>{�	�d�ZhG����{���O��F��8jǎ��.]��{�����#��w/�쌁�e�]5���teO;����W\���'����V�&��7��ʝqF>{��l+�T*�]�Y�ҥ��/�r�%*��h����'W�x���k� ���3<�t�����Ц2��e
K���&O~�[�3�Taٲ�◾4�jgwyo����+��ח2'��ϟ{n!�K�Lv��|���̌�u�H�|m�����۶}����.�瞧 -C����Xq�1۶���|��M*r�ߕ?��� ���Iw]{mo1��^���j#�_2�<9�P}��r��=�hQ!={v[��HϘ��ᆾ�=����.�L��ưo�ك˖��rݺM���V?@�GV�Z�`۶���V�Ӷ��S�%Kz��{X��JϚ�I�H/�];�J�v9������R���j%���r���f؆6�J�b[�����C�V�����p߾�z����}�-#��	t����u>k˖�j����LfΜLa��ԤI�Oمs�f�U��m��;Q��H�n�PɞrJ>ᅅ��Z�p�Q����N��W�%��{����n�t�m���ݑ?��c���^����=22/���9�
�\�5�ӷ�m�={jɊj�3%������/��g�]H�S���֟����Ԕ)����z���'����]]����3��	t���#������CIe2!�U��SN����͈)\sMOchh��c�U���Q�<�t���˕��w�N>9�|}��;�|�Cyݺ���1v3w�X��O��v�_ �%����˖]?g��O�6���I�/��|��=?�=��������;��p�|����^�毸��Χ'�9���}'������ڶ�X������� @�:�[�^��y[����_������W��M���{����]�?�+_n�UF�_m۶���x {�y]�E�
�}�b�����v}�}c_��p�oDe��¼;�t}�Ջ֬ DG�4={㍽�6l��L���Dr�Ua��d%�H~�s�����)�w�h��ֶ�o{,&׽xqwj֬�~=r��f���~�H�S D�0::{ڮ]�|�� @tZ�"��ҷm۟��P�ܹ����~��!{�����ݵ���� oi4�&Fo�u8��r���ʫ�i�2=�_�W������`ԑ>iϞ=w�5�s�׾�� @T:��x�oM� ��t:�/��;w���ݞ�aP߷�^{�5���;�z(?�D��ys��dIOjʔ�=���<9���O�׬iE�sv����W�xn�ڵw �!Ё��|�z͜-[~!����ڗ-��.\�1J&�/^�ӌ��Ʈ]��#j۷�F����WvgO<1ί�C�������WLΤ��o����۷�ރ˖=s�u� Q�@����+�6_��A�^o����S]�^ۓ>��\�Xr-U�u���!�S��h�R��n�h}`������V��G�������pĈ�����㇆���M7-N�|s��'@'�@��������C�Kuw�����7�Z@��ص|yO�_I�7Ï�<�l�鵃7L�|Dn x�F�'>�;��/G=8�op������j>u -�b�p{f��_��u������%+u����[j@z��\rV���C� o��曵⭷(,_ޛ�?�%_���z��^3񎑣v��_֯Z�Т;�|$ pD��<���K��8gǎ_-�+t�:T+d�ػ����xIԖ�c8����N�n��H�`�Z������r9�HO���}�x��/?��[F G�@:�m�����K�Z�
-�Ӣ�[2� 9g|p���M� o#�3�����޽��%�t%�C�Iϙ�M��$o6$�>1*���*l���ͧ� 8b:�QNٿ��{���v0���{���e2��%KzFo�-��q���.���z���zZqx\�M?�|yoi��hg/�x�ͫ�����Ϲ��� G�@:ƣK�^q��@hao���%��C���Nw�X�[lFz2�;�;�|������Hr.=� �����G?�]~��Xg/���#���G/Z�f[ `�	t�#��ս�������W��zzRݫV��T�&9�[X���t�]#&���$�!J_��pr�;ys'���g���*�חB���r߬;����k N�a~����bqFhQ�R����ZmZ���=��\㢋�ʏ<2২��Q����dBz����"=��]I�W_}�"4e��3��.ι��� �Ph{�W��d�ƍKC�Juu��>���d�9��ܹ�{�Ԓ��~���ݵ�d%�������T*��暞���pm��(���y���<����k�� L���dj���[��U���2�еbEOz֬���ߵ$\����>88\�2\�G}Ϟ��HOv����T��r�T��z�_��p3ԣ;ב)�{�����O. 0a:��N޿�s����C+J�B~ٲ������I2�T!w�Í��Dz�;Fz>���;����'ׯ������h������gM `Bt�m=~�u��޼��Т�_ޝ]�0:P�����b�V���ص�6v�]#�d�{�MwOϜ�)\uUwiݺ��F����k�o<{��ξ喑 ���@�:j������Zr�9����YgBK������t｣�R��$��J��3����j��gO<1_߾�Vy��&����;����_ Ɲ@�ҳK��Z�m'��|���]pAW�`�$C��O<]���W�=��ha��d�Ah!�K.���U�m�Z���k��G�.���{�}( 0�:�v_�z�Qo��OB�uT&��-�)y�������&��3U_z���4i,��ݡ�$��,�)�z���H\[F����}�~���K�_���F�q$Ё�3m��?�T����ח.\{mo2�9�wޚ�^ۻw89k�g�<�T)=uj:{�i-uL$�|X��w��ۇ�Qb�=22嵐�_i>�| `�t��<�bŅӶl�(��l6սreo�=��7-�������/h��Ƶ�H��=TLO��Iϛ�2�u����R#3kV&���g�����^���qǛ�q�2?� ż}�~7َZL��+�;���(5yr���c_��p�]���kd��G�o�aR�bR�7�����wגG�3$	�F���O�r�g����6��� ���@���ҥ��o����;�B�S:�:�w+=wn6w�U=����J*�oi�ڑ���Kv��O�Vk4�7߬%C��;v��V�>pƞ=W=�bŇ.Z��;��N�m����6mj�k�2��e��́C����h�N�WR�$�ˏ<R�_~y�x�Y����޽�Z�Ɋ��=���v|��9CC�k>[ 8�:�&�����i���z{S���{Z����/������qctWR�ʳϖ�s�d�'�|�v�$��k?�E��k����w�S˖���u�n Vhy.[v����W�V�J��%Kz�����V�N�����/����(��)=�P13wn&5eʻ��P�7##�ڞ=�z�M=yT;}X�={~�����O_�� 8l:����t��R�)��?�+}�ѹ�{W(�˗�o��@htt+q(��F��{G�����q�J��O��љ����6��^ ��@K{|��s�n�z~h!������k�7b��1#�=���Z3��O=U�_pAWG�g�w�a}��Y3 8,:��f�N+]����>�5;٢x_���ʓO�U7m���_3/�X����)S.������� 8,:в�\��ɯ�~fh!�+��N����
Q�V��~�T~��R(�l=�ݩ׃8?|f�޽�U�>��w�	 �ohY3�����-��=��|���w�^5���/WJ�<2��D S�v�IV�- �	t�%=�bŕ�6o>�U�OS�&��]�����uk��������Cdf��}�W���w��f �}�@K����7��X=O�T[��;�:xwJ�z��G�*/�P6��ܢ1����l>�� ��"Ё��~Ŋk&m�|B��Z����]��.U�x�R~��b����!r���Y�~�깋�c{ �=�@˙�o_묞���s^�8d���z��(V_y�������8��ͧ�< �	t��<�|�u��7/-��Lm/Z�̈́T_z�\���)���g���W?�z���ck �=�@K�58�2�3ٓO�e,���PT���=Vy��R ZR�V�MN��& �t�e<�bŇ{7m:)��TWW*�����~�w�J��;R߳�Yshq���fݒ%���w�P �]�@˘=:��C��{��袮TO���?��-�_�z1YA@��T*=h4�e�� �kh	.[v�m��- 3{v&w����;jT*����g�}������_�� xW:��˿�������J��e�u�t�%V���dJ{��Gj;vx�m(W,N_02��ͧ�= ���b�x�y�i�v]Z@��S�|���w�ص�:z�]�ax�yshc3����A��k^Dћ�h�r�\��Z6��_pAW�mU_{�R���Q�͡��8p�˖-9ݺ� �L�Qk�tSz۽��
- w�y�ԤIý��sϕ����m�b���?k~� �@���SO��c��!v}}��9�?��h����b�g��(���?��+N�x�ڗ �D�Q�64�B�_|qW*�3�����*V_xA�C'����J�_j>�L ��t Z��Z�p�ƍ'�ȥf���N:)�;I�?�`����s�`S��r��>�[���JE�C ЁhM���
L����p�U�;�Z�t���8B�\��ٶ����� ��:����3��x��̜9�����@���7Z}�Uq4���䨒@8^TQZ0<����ؔ��v�T��y�^o��[7Z{�5q�P���iɑ�K�� �O%Ё(M�!D.3o^6{�Ξ'��g��9�������O5��z ��@t�q���m�|Z�\���]����㏏�����/n�t�o�n�� xG�Όb�b��=;�=��C�*�?_*?�D) ��|�4��'�\�|z{ �yq	Dg����!r�.(8{B��W��*��a���?��@T�X���ܦM�C��3f�����g�k۶U���7� �L<sݒ%���w�P �m	t *�GG���.Z�������=��4j� p(ҵZnn*����� x[�ʤ���C�R==�܉'v��yr�����6FG-��ʤ��A��#�D�U��ɿ������gB&�ѫ��o~��lo �R߁���ʕS?z�]� ?A���9p�?D,�Ʉ���C���R����NxOҵZv����5��� �O�@7ݔ�瞨��gN>9�������T߽�V���Mlޗ��� �ޖ@���SO-]P*M˝uVǮ�7�����w��jչs�}�<u�7�\t뭻 ?B�Q�:6�����ٙ����=��o��� �>���L~p0��? ~DǾ��qp{�ڵ煈e�<�cW��[�T*/���9p��8�ls� ?F�GܓO?������|>�9�Ď�F����׊�ag;p��8p�7��{�-�� ~H�G\_��4D,w�)�T3�C�<��h��[ہ�*��^ٻ����[ ?$Ё#�wx8���'�ܑ����^�T���J ��Ʈ
�Gt��zt���=��>?D*5mZ:=gN&t�dk{��G�8�>; �#:pD����z�w�gO9%R����^y���訃���)�3[����� �A8�zFF.˝tR.t��޽��sϕ�8�[�� ��"Ё#���N��̛�MM��q��K��F�Q���6it�� �	t��y���?rR�׫e:p����k�ڦM� 0��������<�5� Ё#hZ��,�*�
�:+Ы�F�� $]�����U�_	 t���97D*3wn&5iR����C��gJ��!w���T�"t��:pD��ߟ�~��cB��'��Qw�'תU����	�S,F;�`�	t��)/�]�E��<��v����sϕŢkՀ	�5<<�9t���Q/@�x��˗�H�f�J��w���F�l�8bR�zfZ����{@����],�"�=�����X��w��GTo�|i� 82�GG�He�=6ڭ����s �ccg :0���Ss7Fy�y��+��3�c��W�="�}����M7�S7��&	��	t`��T�W�He�9&2�T��Z���3Vρ#.S�v���n>�N �`�p�b��!R�CT_{���zD��ZM�C�@G��@<���B�2G�1���=W ��;7 t��y!
�!����7g����SS�t����޽�ڶm� ��bqA �p�P}����^O�e�=�c�'V��v��ȏ��|�ӟ.���/��t��y1
ġ���P�Tz������\�Vy��J �H�^ϼ�qc�3���CuċQ ݕ�I!R�y�:b{{�WʡT�|D��VKΡt�c	t`B��ƎJuw�R�'G���p�����s J]�ʩ��	t`Bu���Jϛ��T���������aP��:0a��b�1�M�zB�2s�v�����P���#}`�t`���R�He���@�����@����GW��}�w� :�@&L�T:+�(�
�Y��>�mob�h4R�r9y3��@����*�?"��4)
��g{;�
�����\�t$�L�\�2'D(={vۯ�'j��f{;�|�r\ �P�0ٱ�!B��j��u���@����Q�C	t`B<��ߝ{����m���۫�Z- �.[.� J�"S.����=㙙3���y��9�"�Ҵ С:0!ҕ�)!B�L�o�ĵ�ږ-h	�j��5�S	t`B�k��C��M˄t:ʕ�åQ.7�;w����t�|j�@:�@&D3��e�Mk����ρ��U�����p �0��ryn�P���m���@K�T���$Ё	��Tf��;!�w�|��|��� Ё:0!��r�Sy�0 ��{�@ZJ�\� :�@��m�����/�����Ɓ�F�� -$[�N H��nA�:;4�MJO�B������g��s���j�(��ow�J%�q==�������a԰�hA�j�; t ���t�e�;�f����h͚b � w�o4QNp}}��v	t�%�FG�7w_ D��.[��Juu����P�7���@*d��$w�t���\�>=D(���ց�m4jЁU��j�8w�z}j�Qww[oqo��s�e����t`�e��(=����+�����t����q$Ёq���'�����Ȉt�ee#=0�:0�R�zW�P:�o�@�@�J7�B:�@�_��1���=�mqZW�� F��.�hdB�R�Bhg���,뛻 �H���q~��f�z=�JVЁ����!Ё��f���#�T�oq��ha�:�q�|���t�[�C&�O�)���-+�u*Ё|��]�g�S����+�Z�@�r�D�zt��J�C۳�ha�Dw�����J�
:в��/O���.�@o����z�ahai�t �����~���^w:���6'�'	t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@ xc�z��h����N��t� h{ ���̮ry֑��q>6�P� h{ ��f2��lv�`�:5 �8�  ?Ŵ\n�Z�gF��I Ƒ@ �f
���R�T�w ' �gH��8�P�5P,U! `t �C��>��k���؜z�  ��@ 8D�T�zT����RiN8�� ��@hc�f@��j��\W:]ʤR�����;�g����k ��ЦJ�z~W�4�B.@�I�Gz�щ�3]��x� m�X.wm/��[pis]�tqv���H�ٮ_�p� m�V��GJ��Z�b�m��N�%�Տ����5 '��&��jn��:@>�.%q�:8j��q� ��@hq�F#526�]�ם5�#4_�T���w%מ��~��E���J����Usg�����)vN���C��5 �ТFK��r�jK-�q�M����HVғ�Ut �+��b��Z&Y5o4� "��d�:�NWB��Q��Y*�� �����˅�JŴh:M2���B:]J���!q�@ �t�P����cc=�F����1;��ՕN�B�!�v�J�Mp�p� �s}�lf.��'�)�%q��T�U�� �)ק���r{�����7K��c�zw ��D�D��it�������p�ԮRiF�^����J�D��it�f�N��B��T*�F���  ��@���� ��t���\n���Je�jur �q �"��4�;��U(���T&U�S ��p�>�V!�����w'Pr�����޺u���־"6!�@�ق��8�$�U,���L��=g�9�%3��ɛ����x&�M���l��xc1#��lf�@hi��[�w���/T�,KH���ߪ��{�$Cw�������C�ðk$ �"��Ev��w�f#8t��mW�zސU;��<�0��Vg
  F�@�q|�;�eUM��Rf�� �&!���8>���&��qn�Db�ry۪����+ �It h�O~'��pn&3�XV(�DQz[�B� ��@���4�������m)�
�@~�t����  4� ��i���yڶ}1PE��JeN$��
 ��#��A�R����ߣf���=ۮ���(�u��� Z�@ � Sځ=��<�8e1���-��@�7�  -C� ��tݝ9�)������R��+�&� ��"� @C��R#��T^T��J�W ��t  �0}��h�뎋��*���(�
   � @Ct��Ā뎉�vT�3JQ�  A� �i�y~���C��@>�  ��  `Zem����j���&��W  0�  ��g��ٞ�C5��=cA�/  �@  �"mە��7d�6G7O>�F�`P  0�  �,���M��bfwT�3  ��  `J�`^&����@�0�U��  ��  ���Q���m�e�b�ry���  G� �Co4��\��@�(r�U*�U�}  �G� �C�t�{�]�Q��Z��!� IB� ��R����ۮ��B��Qmy<  �A� �I��N��9NIG���\�r� H ~x ��6��]�S�8�\*�	D\  �t  pP�S���T*/R"ֶJeV�i  �t  p@q�������(�  	F� �wԝJM��j{�2�EY  �t  �_9�.�tݝb�8��Q�%  �  �SƶK�<oX����Q�#  �	  ���mW�x�v����<#��7} @!� ��o�s=o��8���� �  ��  v�o�y�̐];V�<A�5� @"� @M���r,+�0;��3 �6E�  �D����͵�@T
��P�:Kj_*  �@ ����<m۾�Ei� �	t  :����=ۮ���(Jm�Tf��|  �� @�R����ۮ���(r�T*s#G  � :  j����$
�r�V*s�s @'!� �@��ΞT� ��܎�|v �
  �@ ����R�}�;!R"��s_��  �at  :HO*5>�cb ��*�Y�(� �D� �!�l;?�uG�PC���re �E� ���]��y�b��ʌR� �F� ��<�.���b�a�(DQ�  ��t  �Xڶ+s=oȪ-�6�N���^  :  �*�!_59��|�g<�  ��  �!G$���ٵc��3]#A0(  `7 �6Gy8��9���
a����  ~� @�D"�mb�Rf�W��9  �@� �>T�mA�"�rl˒�R��W�y+��ry۪��R{  �@ �=�l��q���ݶm�+�ű�(��S�]�[#��J��U*�9  �@ �d�h,�T�@�\EV�+���r�ߧG�u�����r��Q��q����  ���  $���q�W��c)�� ��)ǩE�mw��!�o/T��Z�̉j� �wB� �`^M��*5����n�W�������1��1�r{K�<'�~ ���L  *E��*���^���G�-�*��@hY�  ��B� �@n�^�@*��e�G�9  �B� �0)�ʙ(�C�l�/��  �I!� H'�*z�v1T�q�B��  L� @B�QT�EѨ�d۽�ee   �p���yٶ{��
  8d:  ���
rQ4"����S��.߶s  ��@ �`�Ra-Ε22Ϋ����v�  �)#� 0�R���8�#1�oۙ�m�
  �:  R��8�m�B1P`�^ɲ�,  Ӆ@ �0:��ȹ�T 
,+]�qn��  L'  ��8M)勁�8w���oQ�  L;  �d�h<��(��T�8 �at  �ḫTYY�S���,[  @C�  �����R%1����8 ��t  Z̍�B:��b�H�.�qG�#  ��t  Z(E�L��@J�*;NdY�/  ��� �ERJ��Q4.�һ��q�
  h
 ��������綝  �4:  Mǹ��:C��/�,O  @S�  4��T���U[�m������  �t:  Mb)���[VV  @K�  4�RQW�#=Ul�ˏ/  -C� �h��yղ�U��  �R:  �bq���J�b ߶3��  �r:  ��\���(����J��g	  0� @��K)U��.�6q �At   Ec�(����8w����9} �At  �Y:'\��b�вR%�1  F!� �F�(�{J�@�e9E�˲  �@ `��QT��� Rq��  ��@ `�J�2Q4!R"���8�  �"� �"'�*q����t��g �,~� `8~X@�ahEJ�	W�����:C����8w�������D hk: L#��AP���=G)?kz��vZ�h�ue�XLg���� �- ��5��8W��w��:Ȇ�U�En�����	�F�ZM�a�t{��h: �' ������wK�0E��y�qz��ڎ~#P��g=/ȥӌ�@�!�`
��Ӫ�;Q1j�)��jq?��ʶ��[VV��J�JJ�)؝���e�F `�t 8DLi�<���<�C�@e���m�K���M�S��T��7�  �C��!`J{��q�G����V\����8݂��gJLy�6A��$0��c�8M)勁|��Tl�Wб��w=�ޓ�2� �@��Ĕ�Ε���8Ϋb�����m�	:��գ���d2�� 	E��A�@ǹ#�8^��q^��-��w�P�g��H�#=�F�  �? ���+�i�Jb�вRE��b�P.�a�]�Ǻt H ����-EyO��(�,�8ǁ����Ql�K�� �`Xo���q�{QT)˲u�K�(��ץ�f�UǶ�t 0� {�q�G�)�T��	1���mƏ���A��Kכ�q^: ��@�=�͉��ޱ]�D��m��8z6�>/=I��ccG�s���;��� @� �`6��lvU�Y�b ��8�#�r��y\�z.�6�(r<��������o��� � : H{ĹU���퍠�e���߀"�o��(2rZ��[Vƶ��V�,0J��H*���3	;�{A`-ܰ���>��n�� m�@���i���mWu���ʶU6����W;�-�<��M�R�tM�𮧽wg2���T�z�'߸��%_��w�
 �1@�R���U��_�z�w1܌��t��G_���+g�������CE��H���8���q�z���\��H��ysߋ?����e m�@�qt��K%��8��g�'!����ү�}����B �� :���8��t:���tJJ��wU?������.�����
 �@Ǩǹ�e� ~_=���t�2�U2֜���?�ɇ�r�M�	 �@G�q>^*��04�� ZLG�~�4}$��Xt�O?��{��r��h':���wk�Mk'����n���s�l�y��{���$ �&t mo�\N�N ��{�\vM?'}�sϝx�y������� � ����L}�) �I��[���<��)�Nɜ����q�����A  �t mKǹ�� �!)W�)�a\.�66һK%g���7�O� �@Ж��M%q SW�TR�e���b�y�7�\���{�y� @�� �N9s}C) �iQ(�]'�t7���P�=��}���W����� H(n`����� ����_[��k�m+1P*������{���&�^�T:����:� ��!�ۯ��l��ץ�h������>?=Y  �t mC�uE��w� ��0�E��g�/|�ٕ�|��]q�-� H@[�;�s�9 4�>�Ro�i���nI�#�|㟯���/]sME  At �ǎ� �\���>ct4=����OW	 $� ��H;�@��9]ǉL�4n�sϭ��������w
 $7� Ko
��T� Z$�kgw1��V�s��#� �@�X�ƐM� �u�����;���@�6o����>t�_�uק �@�H�j���� �Rz�t*ŗ����>��Ǯ�����k��, `8@���"S���J%�r�Ho'��.���/�p_�t� ��t �����r�8 ���F��������Q�x���ꭷ�% `0@�*֝��j��=�C�{����3 F�H}��y� `.}쥗J�&�6��7����/�{�M �P:��`j; ��ԣ�����O?}U�@�0� ��I�����l���;�5nW������?��5}�]	 �@`<}���M
  ��k�>z��]�g<��'���K��Uƭ� nx�@�@�(�,=ս7�5n�����������~Z �0��0��&�G� �(~��rS�H3���?v�W^�(: �� �)e��U^�  ��;�JU�0���_?����' / c�q�1 $�~7vø��� �at F
�M�� �x�n�Gѯ��?��w��9 Cp��H�J�3�����+9]�g�z��������: ��7 @[�3��4wǶ�E��}{���;����m��� �t �)2� ڎ��ޓ��b���^�j�@�07� ��G�9V �O5���a�q�:vmΦM�x���ꭷ�% �b: �0z �K���mX�;Q$=o����� -ƍ0 c0z �z6��[��������]_]��  �B: c0z ���wg2F�E�V*vjh����O	 �7� ���9 t=�����s��6n�3�#�����@��;��6�>{h���.8�+���) �"�h�0�,�=��a�(���x�6���)��et -�w� @G���q�P2c�Fvr�R:���g�
 �����L��b���y�}�on��j� ���=��� @G�v-orS)��E�n�����@�:���0� :V%�}��7	 ���e��j� �����K%�k�����g�&#���� �H���Qk�3[�|.~ �4��e|F����BM���[�	 � ��%��@l �K����c��LsH}������  �D:���p� `�3!�Nb��qj���?� ��@�Lo ��YU�N�I��m;^ ��t M��v ���4�H)ˤ��������/�����# MB�h�*�� �������V��7���~Y �It MWe�9 `/&���� @� �J����v ���4w��X�9?"r۷/ h"@S�9 `t���T$��߹3��W\�}�k* M@�h��N�  �E�+bL����Ro����� h@S�͗  �&����� ��@�4�ctX ��[ˌ�! �$:��	�s ��ah٩�9�>:�# �$:��a�9 �@L[�ޛϻ��zu�W׮- 4��iX 8����>RQ$n�pq��� F�h
}�-�� ����s!�4��)BF� A���7���cc�
 4��)�  p��Fqb�t�0  �:��	t �A���k��c���3 M@�h
�6� ���,�q�]��� �� Ma�zB ����+ˠ@�|����|�]_Z��y�"�4;� �~Sל<�*΍t E�h8F� ����5-�S��) F�h8F� �e�ώRi� @�� �t �d����*� �@�p� �$���$��� F�h�0	t �����S.g �@�p�b 09ƍ�W�i�#�  `�ݭV]�#�4\|��: `RL���\@� δQ  &ˊ82@��   0�io�::�& �4\��pW H2F�4�   �E �F�@�8�DJ���|VmO% ͔��R�?��T HČ�h@��x;�&e۾ hk�(4D��M{��`t��1 �G�h8}�e�] �x�&Ёt ��M `Rt ��@�p��a��� `��g�Q�nY�_ ��t �( `����� ��, �!�g��C�h8�v� �Oq�8�D�h�0�t ���o�_b֠h@��7Y�pc ���7wt @�: `��04*�A�:�����tZ  8Xq�S� :���|�FA  ��Ȩ@g@3� �M�  �p�
�C���ᘦ ��H��0��t Mዸn� �wV	CWC�h@S�J�]�"� �!�� :/~ ����k܀ �@��g���s �bԋ��U��"� ����@�,:���;� (qL<bM	 4��)�Nm�6� `ߪQ��� ��@�4z�8ϲ� �~�?+�[�w �B�h�J�=�!� �U�V�?бx�4�M�ۛ�
  �cZ�3z���z���.Ge��V��| �?P�2�G���t M�o�|�tZ�"  ����ƶ9�@�� ���^�qt �(��h:��*V�i֡ �E/��� ��@�T�j�f: `o��?7�kОt M�op*Je2�U  v)�~F���sF�4�����j&�y: `�|���� ��@�t�rٝ�yLs ��>� 0���s �@�h:�� �T�}�v%����%�� �3qz;�h@K�i�3=O  ����q��5F����%�4��RY��@g+A"��s��f ���D��e�; t��r9��Q�:��ɗJ���c+
 �㔢(��q���s �B�h�|t�:θ  :�x���0R��t -5V,z�== �,A|Z�T1�� Z�@�Rzj#��@���~��@�J:���S3�� d�T2ns8��h5@��e'�fݔR�  �^!���(2��g�3�9f@3� �0Z.w��� ���Rɸ��5F��������y�Tm�  @�*FQ����-�>��s�f@�� �1����;* ��5Z*w���N��5��q ��@`��b1�����J� h;�(ʚ8z~0S�#��h�1�<��jw��	 �팖�F�v�����h�QF�E���߶�� �6*Je�ժq���������% G�0�E�V{Y� �eg��-�rmy�N� �@`��B!�30��� �&��禎����X�J�?
��#�ig��3;��) �DS"��B�ȝ����̞N�1��#��P.�*���,�, ����� ���`Gϵ�u+ F�0�p��=���@��
�)3b {��G�̸ @�� �������l�  ���Tz��&���zˮ 4��h��|.��W��5 H���7Q*�b�Ɏ�ka&�U ��t F��.��fzވ  cG��#�:�@�L�e�#�O�����l 	1���z��HǹeM~�:;��_ ��t ���P�Y��SS3 j|�ԍ�ɮ=ע8�+��� �@�~X#�j߀�
 �X;��>S�K=���J.~�[�*
 4� 1F�t����*�Y� `��0�)W�FNm�e�\+wuU ��@�(C�|��������3 С�����|Vu�q�����)t �R�}k���� �1yj���P��k~O�F�& �$������e-��� `���oǩ�uaOϣ M@�H�����E}}[�P  -S���~�T�G��X�=E��- M@�H�(�d[�00/��! ��E���|�l����l6���� h@b��c�t__*5& ���Q*��Q4����q>�����`^�xC �t ��3��f~������%d�; 4�X�+��O7�T7���Θ� @�� -�h�Ȋ]9����[ @Õ���7H�`S��^����A��!�$Z�)��>�'8�؞��hX~�ɪ  F�w�m|��u�z�|�S�5�7��Z �It ��J��GמGQd٧������x��� � Qܾ���~S�;�t�O��y���z�w�� @�� �������!� ����g���׏D##�  ��P�4�����i��ZqΜ-��K �B�H$'������߯�v*w�y����Ǣ|��! H���j�R���k4]S��*3f�' �D:�D�]�R�tz�wae���;�{�[�R�� 0E�a�3V,��`�9�]�������* �D:�ı����Nz���ݝ���GT�{��+� ��)DQ���DV7�q�+�^w�� MD�H��w�KR==��X���>[ K�`�*Je��ǻ�p:Χsj�V�;w���� @3� �ժ���R��hQW�>���  ZU��2>�+�����5ݪ3f�- �d:�D�-Y"ޜ9=L��_�.]���z��+ 8 }��汱>��SӦ{�y]�J���� 4� Q�O9e�������c{��ձ�/Y �~E��l�7=εFĹ6�`�ȧ��z� @�� #=c��8��� l���ra8V�կ�t ؇ �7�:11���g�k�Xw^W^��'��c �F�H=znM�n��};u�I}�(+=�4[��j#�q��A`|�7jݹ����{{�V �t ���r�s�qS�8z$=�jU_�q� P�Gη��'b�Q����,�5o	 � � �N:Ilם�G�re_��$ ��j����DĹ�J5����p�ϙ��Ut Ƴ⛱��+��c�H/s��\Q �C��ڷNL��oGE��_ h��z�/�TW״�<������l�dY����4
,�ջ�')��)\�؂c�^wݛ -B�0[|3ֿjU�>��H���re۲"�PQ*�el�7	G�i�ܱ}O�E�n�� h����^q�9�9��B&��cۡ @+)��6>ޝ�8o��{*�r��+V���v� @�� �揍ɖ�fi�y�)�q6|ߨ��]]��m mh<{�'&���ޱ}O#G�_uUY ��t W��}�x��e���\���9���ם�Y��pN:���yo�I���.�?Wy��/ ����j�a(S�N��%�����s�mx���t.��<׭
 $\��kW*���+	��8�F.�˛n�G ��t M�o�� �Z����l�?Μ��^,�� �L�� +�,g[�0P�V��{53ε�ᇯ�'� h5@�LG�O<��D������Pv*��H���G�>+�c� $�oY����ޤ�V��8/wwK�/���V�V#�4���#}*jkҿ��ښt�uz�wx+��� I
QԵ}b�+);��5��uԯ������t MU_W8�H�Uټ~����ǔ�N7�n���{.��Y��tcAз3��$aZ���ܹ� A�h����o��[n�yq�;�L������0���.�q"{�T,U*�Zo��"ε�c�y���A �:����HߴI6�]+�?�q���6��R��֥wg�e۲��8 �F�2C�|O�֛k���(�R�/ 0��e�+ҫ;vȦ5kd�(oΜ�����X>���媜��Ւv���Z�ڎ��~���L � :����H�yy��k�ݳ6�nO����S���>Bm�XH�v��q9�-�L �0:���7h��N���\��n�If�}��]��)w}zʻz�;��h��R٭cc=Iۥ���q�y��׭�O �0: cL�9�*����y����f������w��(6vy��5��}��BZ��q�l[£���<�� �it F��H��eٰA��Q�s�9?+�N����y���3��Z �U���^?��V_��jÇ����~�N ��U �2-�˿��2�#Q�������o��~��t �E����~�H������L��0�RGu�l�  `�ֿR�>��0���)}��[oɛ�]'s�H�.XдQ'=�^�+��p�C�[��mb"���)q��8�g�r��{ eƫ% ��8�ǩFzm��u�d�=�Q���ִ�� l}�� &�F�5۶w���Z%��Gq� ��t F�7vz�E��O��#���j�����?�f�K�M0U���B�����5���tS�Xq����� �� ��o�t�O��tm��g��}��=�<�h�hz���l:͹� �@7�H��;Q*��p�����`e�I'}T~�C �� ���Q��Ou�ʶm�u�����c�m�U�Rq*�j�+��]�� bQ�3<1�M��{j�1j�2z�	_��UWM�]^ h0@b�#}:vx�*�z��RڸQ���?;�j��d��[�b1�n*�yL{:�>:mG��S�}s���I���id��Kׯ�� 	`ޫ( ��t$�Vkg�O��SOIy�V�{�*=8��!}$ۘ�g��L�q݊ ��eզ�����ή��ܞ�TJ�-]z�<�� @� ��Y�#[�Cɿ�Ҕ>V%�7���d�{߫�W�j���R���Sߙ��CfYV�Je���ߨ�������YM�aw�Lg�L[o���+V<p��7�H  !t ��x�5����·������~�������\
��������jj�ק��7��>��P�d�#��t�W:I���l!��0�ah��)0q�y���Y�E����ɏ, �:�D�o�g�!���Ֆ�n��X���+����q�2��V]G����(�v�O�ǲ�_ �Ӂ��(��ü�֙��(��i�(���+W^q>�H@[�Z��Z��Ϫ-����7o���
ټ~�t/[�f�}�8�L��@���Q��z�>�����\X����.{���y�������{Z���׭�V  at m#��g-^�Zm��Od�駧���/�(�M�d�?���.m�0Q�Z�˖v�0��TQ���;R.��K����2yJ{]a`��-]z���� I�v?8 t6+���s�tq���.	�S[����{ߓ�NP3?�����kU�w�+K��j�07}J{]};W����o~3/ �@m� ��c����-?����xc�o��g���2���W�˗����L}̡���,���r[�W%aJ{����ͥ7���	 $T[�  ���}�3j���d�=��
�)}<�6}�w��j֟���}}-���w�t�j[#�@3��jqD&Z��{�}���iGI��^71kV�O<I�W  �t mM��>p�)�Y�Pm��v�w���,��7n��SOU���.��:Գ��F�8�۞ڻ ޑ��>��:���=0P;�{���J�8�a���:Γ"p]U8唏�񵯕 ,9�� 0�y�%����~｢GԧJ�������K2�O�De-j����=�2�㨬���HU L;��d��9�،������e�����Oҳf��?��D�d���춝�����[.��w� H8@ǰ]ך��J���P|�7����Аl���Y����\������a�u˲��y��^�(��J !���p��I���?ܵ�אw�g{�;��fϮ�8�u�-i��u;�>���o��S m y�� 0E=�c�,Q��[��qlj�������/H��Wj��N;M�T�������ܹi5oތ�Yg�W��'�,Gccl*�A>��u�q9k�<��堿��Y���_���uW�ƤH⨹V����?���_	 �@Gr<Ϛ��K���j�~4-�]�i��='3��^�}�1�5��Bq�KU�-[֛:�؞��7%��o��Mj�oL'���FFrf�t�ҥ��ҥi�d�Vm����F�͓�_�BTd��I5�B�Q;���/~~ݺ- m"��� 0Mr��֦���/e��G��F�����&���|�>����u�R�,\(�ŋ�L�(᫯J���%��Y�aEQ����,�稣�q�Oz��?�ޠ��S%3��z��Ӳ�f�%uԼn��U?��7�� @!�t<�6}�> =K��Fӫ;vL��-o�R[���z��3B=�$�dD�;N��6���kRٴI��twѢ���]]�a����R�ͩߠ[t�%J�iW��cHҹ��3t�1/��	 � v�.\h-��R5�a��|�ڔ�)SJ��M�h���W�g�����T�:n�"I-^,^�b���-[�S��Fr��={�Ҝ,]�Q}}�{�f�-Ouw[>�鷏b{��}o���:̓r����͝[�,Y.<  �nt ؃�JY3�菤oŊڑl�>;-W��;��S2��sҿr�8�tq��M��k�=����$}���J��z-փ�+��RG��������)բ:���͝��~�������Z��;Y����׬) �! �����{�N8A����6�]�ʏ<�Hm���U����S���������,[&��k|���_���u���,ϳ����%K�j�|7.Sc��Y���fά�Vn��k�0�B�U#���Wq�?# Цt x]K��6�}�	�q��U*��q������2��c���o�z6+�	���]]"˗K��Dv�h�f�n�(A�yF��{zj#�jѢ��Q�G�M]���9�Zx���5kv^z�Lg�-�����S��o�� @#�� ,Ǳ��^�L��g�z�q-���Z�����POuw��j#냃�+�v�,і-���T�x�6�h�8����۲xqV-��̙��I���O��/��C5,Γ�;��l]��ы���� �� IO{_�яJi�f���{�G�t��Qu���}+V�F�ݾ>1Um'�t��f=u��QJB�6I巿���Q�~�牷h�8��y�J�R����0�T�����96�ȵv�ξ��#��z��~v� @ �`����[�W���믫�w�-���i��z�z-ԟxB��K�>Gy�1����vWs�_ݧ�&jxX�8փ�[ŏ/��m8D��I�(_�@��{!����>�\��@X*�����KX.7�s�0�W�Lg��آEc�O?�HٰA �� nb����7��6�u��V�s�S��>+;�wZG�t�N<�|��.\X���;��D܀A�Nz�?���/���##m�.�okG7N�vhKvW����+�q�*���2P��-���ܩ�mzԼQ��n��^�g�.�����ϸ�j�� �:��[��h��7�o��%m&�1����Y�L�<�h�����H���i�����ś=[�N:Iz�;Nlו$�M��Ov{�cr���ھݷ�z�Rݸ1�n��zt�Toomd\_�������愱�ߝ��שX��Wk�`�76�ko�0�JՑO<������#4  !t w�w�����.;v��_�ٱì3ŦI�֌3ΐ�OT�zӷ'���Q3=�~��?�����+�o�Jq��%Itx��g�࠾���*�Td����m���P��ysML$��p��L��C|�,q�G�yoo@(��<L�f�Q����k}��m��� �Ogog����+��ºu� �0:���������K/=���/΍���k���Y����eƙg�����y>�#�z����裏֦���t�d�,I�hZfVe�̜����|y��J)�R	Վ�54T��m�-[�(�'�&��#�ٳŞ1C��3Ŏ�<�㲾�[-��?Ae۶��o�=7���{�0ׂL&�8����v�} �mo����k�}��V�>�~��f
���jxN6k�<�,X��a��ש^~�v�t=���jKu%w%An���o����n|��NP��(�\~;ڷo�:ڷo���q%l@�zzd<�;��!?�ˎ�\��I^r���Y�h�>jq쩧��ysC?W'�����z�_��ڵ7	 t(@S�7^?�#�������L��֑��C��䓕��ڈP���Q��/d�HבGJ�'J��å֨�F��Kǖ9s���E{ZG�����P����h����
v�؈�1��q��Ċ/[_��qGd�Ǜ%�gm��Im���gd��g:Z�uZ�k:·�:�?}����. ��t MG�m�^x��f���g; ҵT.����)�(�z�F���P�/�T�����˥7��3fH;��"�tw��˓��Q�8�=ێ�|>��x���@FG}dD���ؘ�j5�øf{^mD\o�f��j׮ W��{���{d<j��A����?/z}�t��?�暎�g��w�|� �p:������oב>+��L�D��d2����Gf�q���󡇬��lRLL��Cծ�������Ү����pwݔ�i����Y�ʉȍ� ��P�T>X�bǼ��]�s�������J�Ƿ_V:-V6+v�ˉ��8���R�?�#��������@^y�6R^|��R�F�]��g������? �@�::ү��g.���_^�J5d�R�x6}��У�����a�O��՗>�]O}�9�X�:�(��H��F��N�o���A_���q�t �z>~.q�I�Y�J���ڣT*�}W�R�J�W�\�JEſV���M��\W�L�rzzlg`@?��^���{���G[�1�+������G��I�Jg�G�'^x��S�����Z�y�����+�p��`@K]�nݍ��zuiƃ����3����8��U޺Uvơ�#�Q�v�����r:��z��w�KrG!v��$��v���jI����71tTբ>~n����~{����h�CO_:�j��a�k;~�G�k��a�DGZ:]�������q�ڙ���?������G���8����n�5��v]u���}�����_��o~#a�дϭ�\��w2?�����%7�� ���wc ��פ��g>�'�6l�I���+*3w��?�\���^y�Q晆�S��qX����k�u�wsLm���F���y��_���^C�Z_���\ϲ}���4������d�2�;u}���8����7�H��^t F�|ݺ���袳Ԇ�w��tt�}}��R����I��e��':�]ӣ�zzo|��ܒ%ҽtim��+2�$�Ǣ����\_a�����������˅Cg�y��7�p�  � ����Y�ȿ^x�J��c����Ѿ;�$���^+�����#���Xo䨺�G�wO��m�,\X]���Y�0]�ϫz�7n�Vl��4�?T���G�8��?�f�O �O: �\~��/���a���#/��f��F�6���}T[�F�5�����K6���c�+���a�Im}4�bz������Rx�U}fyKv�g�|�
�f��O:��ϭY�  ��@`�������W�����/���B�n{��O���l����L�F���d�'j�]OϞ]����Eb1b�&�GG��T���:̛����0Z���-Y��]��]�M  �@`�_s���^|�?���'�<��?���T��#��&o�G�+[�֮�j��Qu}�/����ǁ���gs�(ׁ�J�~D���v��o�/?����G �A �풟�����gw�~��?�رz���j�ժX���x�3��4'��̂�+�p�d��c���6I)���[oIuǎ�L[�;�OB��jۊ�����N�_�J  �@`��w����?�ڰ�
�Ze����a6u
���n����4}��uo�<��?_��d2�yB� ��А�u��*���b�|���g�)��~�� L
� .���/�ӟ���o�v�Y铡�BO���ꪅ#�z����K_��@I��8�k���T�hoc��?<,�-[���H�A^��\���B������T��h�������|� ��� ��n�ޚ�����<�xN�Gp��4!�k�ϯ������]�-=>=c���̑�5wn�h7��������Q�U��}{-���Vn�?�(g]��+VFW���Ϯ[�1j p�t �r�7��ʚի�o޶�Ł-[x��q'=IF��.z�q�%��]�����*��>n��8sf����@o�7m�w�J��8�+q��_+���`����y�[�-Z~��u; p�t �s�ڵ��aњl��eo����Vi�h�8i�s�HO��]�W^����p��S�࠸z����To�>���,,�����W���^{�Ϥ)���ק���[��X��'~���e� L� �.��ι�3�����z��g:��S��s�`7et��pף��8nK���=�קGߥ�_:���~q����_���E���z3����s��S�'��h�i�}�����
 `Z� ��u���������g}�]�܁O�=�F�3֍�=(��y���}���_q��Tw�8��=����l�vD������Ӽ^��G��|^�BA��һ�����;��_Gժ��z�3u�q�z�U�>��u�� ��!�$��֮}�_��/�O=�̱��u�щ*�u=֣(�g��u�:H�(/�q��X���qqv:��c���_����ka���z���?���>^=j�8ֱ�{��^z���{:�����֣�ah��"\�o��jA��9ߗv��9�䍥ߞ�y�1o�-Z������ ��"�����[�B�]����#{�+�O>���T��G{҃�����Qg�a��ۼy�tZ�X���շ��i 4�����喿��'?y���w�sĪU�n?w�M��`Oʔx��5�f(̜Y=�O^�n� �0:��s�M7=������'���1����;�x��lﵿI[Î�!���,[������]uUQ  E�hK�UW�֧}���������y�c'|��$�{{=҉�ζ�4u������Fç��O�_���� ��t m��o�/k/�t��l8fٲ9م) �Cl�h��B{�3�O��E���˗��%k�<" ��!�����^�1~�w]_߿,ݺ��9'��P���7�J�'#����9�ğ|�G?��<�  ��@�1.Y����r�%��v�=�8f��~o��!�)ܵ����{s��,��3�p���ҥ���7�' �� �t��_wݯ���]]7����u�)��8�E�k�|]=������o�
�=���F͟|R  �C��H����O��E�0p�}?;v��Y�E���6r0Q�������~�d{����#:������˖�Ǩ9 ��@б._���a�����^��k��;��r]J�CL6N�����Ow�����������6F�NG�W���;�8O�~Z  f �t�o���5���?�x����>��YFӱ{�/!�D��qĶ��G����_��  �B�@��|��a�.�ે���Y|���TO�m����+����JΪ@����:{w !�@� ��sʨ��TTF8#;�g�IUu'3�m�򠻪9�9Td�ħ��qDf�����:.@P���;�T�[�փʖ�Iߪ��ι�ޯ�!��!!�|_}������<�v[  =�1.\�������Æ:*�{���(d��P�V�������>�`�+�y��[ �� �e�W���5מwމ|�Y�d�ܙ�.ҁ�������g��n�r  y�	�s�շ�i�U����E����>���:f��@򆺺F}�����O}jY��7 �A�<�w�[�7k/����6|����_;��uv:���i�j��7�8�ug{���t��a����]w��6�v�-K������;Ϋ��$�����G���E�\|� MI�솳?��{�t�u�{��/}��#=�G!ҁ��86��~�s�;��k�) ��:�8��k�1N�?z�2�k_���gwM;�@��3�<pp��ǿ��O|��� @�� ���7��8}���O��E��_���?�c���:��Ξ=���n8�3�9?l�4;@+� �u��[��}ߵ��~��o[p�1�Y��:0a�b�o>���{�ao?�� h9`�d}}�8�=�z�;������3:��)��B�c;f��|�1_�w��o;K��4�0��C��u��v�}w����ccg.��nzl��#�ڂ@�KN_�~,N�X{�K����?�(�S�:�T�ۯ�(�M;,8s��G ڄ@�������ƣ����+�rgt��:f����m�3gx�s�s���g	s��$����G�/h��N;��j����wN?�� ���c��G��N����' hS`��~�����'��÷/�ַ����:�,��:��Z>=��?���}��m�v֧> ho`Λ~�϶o�#����
Y�ߞ��L�V{�#~6�x�;ξ�����n �+����Y���O8!�7:���'���p�a��|�:��g��r��_�-��3���  �C�$���~y���q=����4>gN��hQ �K-��.ܼ�#n<���.��r ��@H����Gq�d��p�~s�,	�3������MK��9|�A�������O~2 �S� �k<����c��Z-�w�]a�#���1ܳ\. i��_�[-ڴ��C?6#�_~���c v�@h1 6qĮ�;¼��$�j<��iS &��Y�F7/Y�!�x�Eo���[÷� `O	t�&4<sf��B�c�}������0��?��� �]cS�ֶz�C�]s�1���ϖ0Q:@��~����'���+������4dc����2�˅mlٹx��p���~�54�~N ��#�ZD-���,�5��?�a�ڰ!�ݸ1�C7�`�eY�6o���!�|;7oޟ���>���� �[:@�:5<z�	��/�l	]w��k�/~B��'�|�ܹC�/�04g��w�[��!���}A����ٳ��/}�1}ǎ0#�z�����C��:�z#���ܱp������Y7�pS�� �k��͜�����)�_�X�2�G?
��󐍎h������ڲ㠃���?�笫��ݝr &�@hS�7�?��1�g����������)��Zͮ��|�#;.�%?wn錫��/ @B: a��#l>�]��Z-t>�@��яBW��·
u��ӄ�]ڱ`�O�x����˧�;�7�  E�ߐ�r�>���zU�24�6n3~��0;�ԭ[�jdƌ��<�}��[k�g���7�{t�&!�xR#ӧ�G�����y����C���u�ݡ��?��;L��ԩ����oZ��?��s?p�7��� �	t v��y��C/yɮG�gn��� ���8�}~��h�ap���}��)S�\��ғ/��t ���k<?x��F����`����a�ƍaz���fl���^gdY��?l[�0�8䐰c��3^���X,�/ @� L�F��?�/x���Mٱ#L���03�Y7��|�|~t4�[ƦO�<0�xֳ�ТE��|l֬  �B��W�̜F�:*l��^�_V*����s�9)�u���M�^<�G���ó:��E{������A�zd}(�;��i�6 Ю: ���^��8}�W�ߺ��)�o�|f��Л:6o>nʣ�.���3����<��OUuu���s�Ё�
�F�Ϟ ��$��t/��ʑ8]=>~�K�.|xӦ�;�m{Un˖%Ӷn�;m˖S�o�Ȅ{Z��0��~���cx��0�x���9�>eJ  ��@ YoZ��q��ߌ�_�詧��������m�߱�)[�ԱeKW�iS��}�wt����a��ٻ���!�3��P��F� {N��tο�G�t���7�u֬Cxmmh����O�28�8F��8��ǀ�>4��FF|��q4�t͚����{��q�Zϙ��3���G��RN��Ƕ����������ux���Ν/��G憆���?�s笸��1<<5?4�1m��\nt4׬��5�)�M��bX�Μ�k�� ���a4εF�7��Qt �T���k��+N�q�S��[O;m�]�����gg��!c�Ë���룣󲑑��cc����N���2�)cc����)Sj�ldl�#�=S��~}�9��ƗBG�Z-�?��,�5�6����\-�kYVi\g�X.���8������)�cC��S����cӦ�<�SkӦ����?���xI �: <�ׯ�ӆ�U�VT��N��{ ��@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@ �N�^� ��t ��dY6�\.�*�J� �� 4�\.w\�� �Et �)�j�7�@� @Sʲ��8�? @�� @�z^�Ryy�X�j � ���U��q� �� 4�,����������� hr ����h=�˅6����z�����  ML�@���>2u��Юb���Z���� hb ���ٳw�vV�ׯX�j��/_~ �&%���=���C����,
m*~�����>C��u�Y	t hr}}}��J�Ѹ��X�7�}�(.� hB Z@�^0j[��U1ҿ�lt ��@����8�\܇)�z��+����y�{~ ��t hw��@#����~����5}}}; 4	� - F���w�=�˺����H���g� 4� - ����o;%F�Uqo��fw ��@�022�aʔ)��qv�R�+�� �8� -`�ʕ�����,�~Cܓ���~�X��  	� �:�%����^��Z�>T(� H�@��e��@\qo�Z��Jej�X�> @�: ��[�ő��F����k��r�T*]  1 ZD�X|�R��G\�0��#���j5+
� H�@����1B������A��� ��8�"�~u'�\.�K��G $@�@��yG���b��4�T���H�R9�X,V L2� -�^�_%П��OY��1��
��� `�t h13g������������Z�.�����o4 �$� �b.���m�r������ܮh���g,[�lg �}L�@���Z�vNp&��z�����c��#}K �}H�@Z�|��J��ٸ<5��^5<<�����7���� `� Т����*�˽y�Eh솸e�����8����� �� -����;�r��|]`O���\�TN+�7 ��: ��,��:�g�+���HG��� �E ZX��[c\~:.��SS���u�r�٥R�� �� -ntt�='�����o�R9���ki4 `�	t hq+V��'�e%.�x��߲eˢիW��c� �h �@�e�5�E��a�g$��kGFF�r�e���bŊ{ L� m�P(���R\�L��vtt|5��J�� &�@�6C�J�Sq���D84˲��=}s�X�j �gH�@{YZ��/��aN��.��g5�$ �3 ����Ň*�ʅqyS`BdY6-F���j��B��6 �� �fb�&F�uqyv`B�H��H�������] `t hC�|��ccc���&RO�\�ܶmۻ���j v�@�6t�%�<Z�VO��j_n<��0q?/���:������ �&� m�P(|�\.������1�s1��� <] �X�TZS�T^|}o8��k׮=c�ҥ# ��@�6W���4˲�屁��G[�n��z��-[�lg �'!��͕J��J�m1ԿC}��D;eddd}���D: OF� ���~P.���7�150��4<<�����m>��� �.�R�K1��,˲&\��7wvv^#�G��x: �k1�?#����.��]]]��z��q] � �۶m+ň\��������8_ �1: ��_���3�,�%^�,�7��R�<X,�w �q ��7�W��7���������-�ˏĽ��  A� O�P(<���r>��j�<<�7������� @�� ����/�ks�\#�&T�e�8n(�˯.�J� hk xR���?�T*o���_�1�`�͌���_~��.�䒻 mK� O�X,�G������/�&ڂ����]z饿�r��M��$�������;��r���eW`BeYv̔)S�a���'-[�lg ��t �i����z�Ry]\~>�������W��� @�� �n)���>˲����PqO�)���^*�> h+ �m���_���z��Y��W\���{OO�W mC� {�T*}�q<X��Ɲ���	�sJ.�[_�T^\,7 ڂ@ �X��oƈ|M��/Ĩ��0q?������ޗ���� �<� <#�#ت��k��-��L�������j|�� @�� �3V(n������s�&ҹ�r�+�R�#��&��	������/ϲ�qN�с	�t����7����3 в: 0aJ����j��Z��x�����2=�����/�yt��%��	U()��'���8^�1Џ���"./ �$� L�R������;;;��a���D��J��o�b�� @�� �^���7#��鿌��,0!���n����I ��t `���^��{*���bX^C=<#qg�qݺu�^q�駏 Z�@ ��b���Z�n���8*̟?����}���s5 �2� �'
�µ�ryS\~"˲�g�oW�Z���˗o �� �3�R��j���z����{,˲i�Z�ڵk׾t�ҥ#��'��}�P(ܶjժߏq������3�[����� MO� �\�������|#ҟ�c�z�}�j���B�� @S� �����o͚5��1^��#�G�/����}��[�hR �4_|�u�֝z�=�����
�Ϛ5�q�P �i	t `R������J��J�sq�.+��7�J�_ ��@ ���w��vK��q����� @S� @2��J�7.�o�����j�zm�� 4� $�T*}qժU/��j�������������k�>��� �G� �i�V�VOl����vǱ�7o�(�W ��@ �T(~�z��W������'��\.���/���K.��� @�� @��-[���������5Y�-<]�����sO �it  i}}}�qzW�\�Y�/u�����q�>X*�� 4� 4���18h��sJ�L��o�8; �: �4b�_300p�O�ˮ����tF��===�	 $O� M�����j�5�z�q��'������� @�: �t
��7.���W���ޒe����9�R��X,o $M� M�K.�3F���#������7��) �4� 4��w�"������獕J��b���d	t ��uww?p饗�����s1D_x\�w��( �,� 4��+Wn���?)��5"�����-�V�:n��� I� @K����#�1�?c���oˍ���E�� $I� -��W�~�����w�]qON��˺W�Xqo  9 h)˖-�#�u�����cu������ @r: �rV�X�9F��1F��e�K���իW��e�v �"���4�'utt�/_�%˲�###���_ H�@ ZV#ҫ����������~� ��#���V(Y�z�I���_Ͳ�@��V�Z���˗+ �� ��e˖=X�VO���_������q� 	� @[(
?xm.��r��/��,�N���}w__�p  	 h����Y�V�R���)����tvv��� � ���R(��\.���%i����  h;�R���s�,�?�������.�l���� �N� m)F�+��qY�kz>���8_ �t h[[�n����zN\���ۃ@H�@ �V___������|��xy|hCY����5k:/���m�I%�����ӳ�\.�9.�cu^h?S� xY��� @�+�J?�T*g���B{����A�L:� �ś���_gY��L��_ �t `ܶm������1XO�������{zz~ �4 `\�q�W�>{dd�����F�,k<�.�&�@ x�e˖=X�TΫ��7�h�B���r����I#� ~K�X��\.0./
m�^��$ 0�: ��ضm[wWW�k�����,;��.[�bŊ{ �B� <��������vy�=�˽8N`�t �'�����J�rU\�3���@�t `Rt �'�eYw�V{s���s� �K� <�B��H�R���PhqY��  0i: �S8�C>z��w/�{Lhms�����_J �9� �N?���r�����Dhq�z��8	t�I � ��b���Z������e�q�v `��  OC�z�\^�kC���$�  O�ԩS�W[���`�t ��iٲe;���5qY-�t��#� vC�e7����� L
� �
��w���q� ��Y�I!� vC�eq�J�qyFhM`�t ��T���=�zKz�޺ �B�L�����-��'����5�Z�;� �D�L�+Vl����t�,k�@��۴�k�NY�t�H `��  ��X,��l_��k֬�ܺu딽��\xᅣ1� ��@ h_|�}��\�2 ��	t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H��@\��@PD    IEND�B`�PK
     �9s[�kZ��  �  /   images/6608fa58-7afa-4488-b64c-2b761d69d6bd.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  �IDATx��	�U�ǿ��ʪ>�/�FA��V�i<vD@YqWCא��Y�q�Й1�u��	cw5vv����@Ggt=wW�G%D9�� ���>��:�z�}�UM�4ts��������ʪ�z����/*%��@$S�d*�LE ��D2�H�"�T"��@$S�d*�LE ��D2�H�"�T"��@$S�d@v,X ������u�a�y�3!��sp����C�\��0�$-�P�������	���ǡ��2�YV0V�JqS�-��;]���jl���i��l:�L���*8g�z�����A8�pǁj�PUu��
���bg��Q���ld&.6S8NW˅~�p>ö��5�̄L��i�S^6n�%���f��ɓ!���0����_�����\|���wr����(AQT>��G���H"���5l/ۺޮ �C]�ee0���@FI��W_�h	.��:aiZ=��?������'�
��+�m(�(
�;�<�V��<��7��{��&���`綾��@6Ȏy󠼵���cS}���m߇o�`�b���Ex�+'��)��{��8�@:m��Zfs�����5�~����?{6�ߴ	dRA��x�����t�������=-ŷ2^C��\&5�lV���!jn{�koݚ�7o6E"a���h-W���OWQ~�ZW�~g]|��;["(�u�"(9xЃa�j9�U�a�R�x�C(�Q!	�!8����J�WTp��!��Յ̵k���m�/�4Y���b��?�ٽ�Ν%��
���҆*��Yy�ʤI�~商��Y��O�L�Nl*dI�	�G��ٳ�|�X�
�����Q>n\�\��a�D0%��>�Pno>��MQ��_uL��(�
����]���R۟#�� ö�6kVH�??���,W܎��� �A!k۾ݴw�/Եy�f��M��0/)�w�I"p��2���Sn��`�2(p ��.�ҝ;�MA��d��� �A�K/#Ë�7B���̫�&�x�����;PUF�%�rZZ��u�EYY��R�?_�%堘Hw"Ɣ�Fm���0��ud̡C��؀���џB��@7�Μ�!�L��n�P%�dI4��	�J�A=��к������o'�˖���C����Q\��%�ֹ������l�5�NC�8�/�L��E��{�3&�*�t>f��/X`x�a�u2��L��f^��&'���	�k1��LF���ffv?ʆ����v���.�Ik�B�(���c�u���Ơ���:���+�x����qج?�)c�Y�F+�=)aǻ�9���yO�)�i.C0/�`^H
����\�Xk`'���ۧMө�;
����}Xy�4���;����4~�����(���D��;�d�=��"�Ǥ�!*�����k������I�� ��c�?����5k�
Ⱥ%K@mj�[�yf���)v��(��*��h	��ۡ�"ﶾeѾ#h%�s��|4&�R`@�����t�������UaFt����[��.�A�3'O����WWC��DY�w�I06��r��=��+��lֵw�0���\�9�55L8RP $��*Z���x A�-}����wWT�S;� ~jr�B*�6�����  ���6fL%�7�#*Ԏ�����r�P����D�ߝ�)0 X	��f�4�[���A�+��m������:P����)/�*|�^�	�c��}�uM�چAz*�T�K�A��)<E>ӓLR����~&�+��<�:�qL�87��E�!�uZ��X�ǣ���\���7�.K���0�
<S�Ϥ��1�pg:j����)���jBUU��� �Ud	���*'9�0����T6q8W���)�ӾaT�z���t)Ĳ��Bb �� B�����8
���4�,��n*U�F�㔠�U��%�� ҫ�Lw	��ya�Q��oK8N$n�U0L$����1
ap�:=$1^��f�;�*�$�
���鵴ㄆ҈ p��Lg2�S.˹w�k���4�`���������EuSҊR���p�A�@Y�"�EnK0�3��i8a��R�0�𣆖C��o��9���B���s\�H�=���}-�K"���	��ؐ.��{c�LF-	�L�/�k�bY��1e
���W�
<ǎT�BP�T�u�s]��{���ڜ�����k�
2�Rð�
����o��f궽�v�xv�,�~c#���33m���,�5�4���I�	&9�>�Љoy�FxӜ�;�G���w2t�RzY$b�"z����0�����[*��U �CI��J�ٱ���;u2�y(����e"��
�m�뎋:�ӟ�xc�w��G���3a��_BP
���?�MP'��Y�����1�h)d�]�۵L�u�]����y����x�3w{�x�Π3n�ݧR��a�Ŷ��]W���{�Z��ر
�#�sf���ꄂNj�/ʼ���=G0�̜�c�\�k�}�l�+�CB�J=�N*9�rA^��]�q�R-k͝㮀�#0 6����g6P(2�H���3M	�cfc�uu [�@
q��(�e^ַ�A�{'���Ye�f.�H�������E�t�.��P8'_f3E���!N����I,ӹ�W�q��w]�9�Ht�tP
H<��V� �g�:�Y�ug�;�[�D����"�p}�����bY4�A)0 =�ࡇ ��Sj)�u��x/ZB��P(��#���}��Gi�;�%�δe�Wsy~�>�U�io�]w�h-kۚ�(4(rUx��{:�sΦ��� �S	�6Z�)e��l4l=��@K�٬�����^J�!Ť5�����@�(�y�)ӄ]���Bt<��(�����h~��ؾ��2�KK;��IOԆ�R�L�̿�� ƒ[����R�4I/;
��*��H� �	��Exh,-��3��r[�2:�pVd4#�aP0��h�0�fiG��w�~J��cG �UU��^S^���,����%m���i��Y�Q[�ɲ�mCɥ�?�7�o�W�\ ����uYc�Q�����}�Z�::��E�X*Y�2�P�T��"pr��'�Ώ�>G7DIE�#�.�j�ca�u�h��][Z*�r��BD}�:u��ܷ��Z%F-\�J�;O�3%����_�����������pnG��ŪT��ٶC+	��h�e��H��)T�7f�>��P�'������K��w킠�T=���a�;[��bU@ۚ5��[o	�t��3Q[��	J�%K"��_���2��Np����c-�!�*�����KU�����	a>u�a�b���{�ݸQh�*%��?JWQ6���>d��C)���<�$��w���������D��d�5�l���]+�^~��&b�fqc�d�>ܞ--%X�"�EO-�*h)A�q�������%:���~��jZG�)��1�`��A����=��E��
 W��WV4zS��9M��<k�HB�E�0�:w���TV�H���p7�%���.]��x:6n���^;42iD�9Bc�j�	u"so�9ArmD�4N+C@n���Hߗ��K��%2MM��k
&�v̀Ch[�R5�ٯ�&��+�@�
H�5�@����)S��k��Ic{�l����ara�1��3��7���م�;T�D��g��3��L--e
Z�7I�������$�]]`b݀	8�8/��m�p��a�7������;�D"N0�'O��?�
���,�Yx�?��իa�����{�Y���7E�����\/&�AA�
>��9�N��--`�Ҳ�U�c}��Wn�k*��c!x�y�a<:������:Yta,��.�h�u�ʕ��'w��y�>��g/��g�����w��c��s<���{��π|X���z�6�_�=={>�:�2��n���*�Ĩy�����	gc�Xtｎ�l߾���ӧ�_0�V���)�ӹ�з�#S�9?��'Zi��[)�-A��5
��J|�^(�
6S�W_�?���5����:5qH�ZU�#�[o���;�t�c,�9�޲~��{�:4�E�E�ob�~/��҆n
Z������믇�o����S�\�
�x�	hŴX�ʙ�#y�Y�8�l��tҕ_|���u�c�!�����She!�|���Ucq���b6�����A�׎jl��"T1M���`�����u�OkS��$
���,��ĈŋW����aG.�L�/�8����$������[�lT�����̯�us�Y���zOj�88��� ��W<����m�@FI	�W9�%�����8x�F zg'�,B��CsC���"13'%��䢮�Ј��Hn �t㧟����G�+d�&|�V@�?�D2�t �ʼO��< �k� 0��!l�`�9�1�� ��Z��$���(��*Q١{ 4����Z����lB.�E��g�����a����l�@�U�
���j،~�o����O�7FB{ ބ6�������6r�?�?���!���@V�X�ulN�`�۪|��Ѥ�_H٠{ $��>P��?-&(��}��m3ZWa/~������/�o��؜���fc��JFR?(侮��_��`s�ӀҬ_0��VQ@H���F~�����b{�?������B�5‐�A�3����!�(E^��%Y�D6 �F?���|���=7��dA/�$�ݦD�D��k4���K�����
�ŧc3��Uh�kH$)��0=�;����@���ө~w
󗏽[i��� �]\}%�>����C�&�� �m� < ��ȉ$����D2�H�"�T"��@$S�d*�LE ��D2�H�"�T"��@$S�d*�L�I�����\�    IEND�B`�PK
     �9s[�����  ��  /   images/2c98734f-75db-43ce-800c-ea69461525e8.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx���	��e}������]�st�3���#�b�uT@�5��!�f7	r�?	��pIV�b�ML�1DA�� �r�r�}�Q�un� YM8��y���~��5�pL�4����y�O.    {�@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@���#�^]޲��o�n�h���!˖�Bn��J����_�j��$$I���$Tw�����
!�{�%�B��{��ۓ�?������Ԯ��ݞI��T�ilI��ͭvcC֙]��uֳ�  E/��n�=�*�5:�A�4�_��[�J���U�i��h���������'�����6tS���3���\ҞJ�ͩ\�ٙud�ƏB{��b��%��n?��� ��@`h�q�����S/it�G�����c�fZXZ�؍;s#!����LxϑVH���P����������y��l�����ٍ����ܔ���Yc��b�w�~���Љ�� `�� �w~��W5�ʞ�ʕ�1r�n�����G�?��J���3�ܢ�v!��'���J�oXw۶\��@!4��7f�/¿�z�Kn<+I� �7���K��x���Px�l(TO��7'ɮ��!��v�3iq�[��Gxn��ϛz?��g���u�<X���ε��
��_��׎�+  sF���N[{m�ޜ}a-���*ϯ%�C�K�OK3͕�!w�T(ԍ�W������5UhO�Yh�|���^1=��_X�� �=B��W>��ۊ߹w��|\=Wy�}ii�V.��\=ɪ�l�����]��}g߼��{
�����2�l�e� �:�@�N��W씖�y:���C��[�U��^�J��dR9<��<��܎�3o>���
��o�3ۿ�����  �6�@t�<���˷����������1�.�� �mL�m���+��姽a�m[���kK��W_�j�ߙ �O����^�d�S=��yͷ�ʡ�0����G��s��	ݧ'����˺o.�w��r��=�ȩ  ���^s�_Z�,[�������KG��
Β�f��v�ѣv��Gmmt�˛����j����}˅��	b �@`��q����5�(�"ʇR3$�ɴz�d�������n�A�>�K�v����[ 0�: s�m�^�����Znd�M��3[�Ţ�]Z!-�HG��Q=zˎ�o����+5&.���_�� ��@`μ�c�|h���};����nr�����3[x��]p���w�K~j˧>���� 0: {To���}��L��)[��n�N�I����t|M:2��7��M�a�����:+IL``	t ���~�ۇM���ع�۳܂����h'!��F�;F�t�w��;�}�\m�y��	w 0���s���������g�$���93���&�k���[޺���*�����/�F �!�x�v}۴ߩű_ڐ�V�G�U����;��߸��-�o��?�����@�� �_Z�Oc����OM��u{)7`/����j�}��y�x����*����#ݫ@_� <�S>��e~0,:��OK"SK
�j��M6Z�����.�uv��ŧ���  }D����?.;��`��nJ��V r��U�fco�:�_�����S�5��}� ������/_����w�g_�NR�+�;�$)l͍�1M�v���//�6��E<A�5/� �7��w��٬�����_�� }����m��r����~�u_)�n������[ DH���������ژ����b��Ls��a�M���׼c���>��^|։; DD��3.��z�u֦��Z!��F��[��5����ε�^�\|��_X��  `H�r�5﹭9���\nQ�!�Hr#�sK�_ٹ��O:�z�/��o �e`ȼ�_e����6$�B'�P�N
+�K�����𴱰�7/x�17 �K:������F�hk���$$�7�i���N���9��o.�l���O��  �L������������%k����NB�-[x�T�����%�{���t �@`�:��]�`�_gK`��C6�5���򎅯��k~�/N?��  �@��Sνj�L~�c���tz���VKK+LW^�f����W���S��
 0�:���Mg�VXvF=ɍ���S��t[n�	����N>�?��/��  sD��S�^y�d6��I�9أiaѦ��ߺ�_ko�UC� ��ϝ��w��އ7%c�5���9�;.�#]xl-��I�}�c�|��� �A����'�x�����OMeK����'YuSa�{˺�~������O�C � �ЧNYw��'�n���i<-c�,[�(��<�jm�l����	<�����f��WO:�[��%|�� <M�Ϝ���%[��k7��/�̴:��,��Uޛ���1�jo�j��O6��Ѿ��j)�GWYesq��9��Wv<����	&��	t�>r�9_�C�U4��-
��L�۝����h1˺�,,eY�q�x�����f��~��|`g�y��fs��v=�O�Mߖ-<�4V��=k���{�x�:@8����l��){c��k��a���q���\��^�/��?���[��{���ќiu,�ẅ́�������]��#���3�Jod �t����]WΟ[KF�0G6L6��,yx���Ti��k{����Φ�f����[��Fg�����������3����y�����w �M b���K~��|�9�;o���d�H.�{�pU��c�պgk�q��z}���n��L+����SϽ�7.��1_ �:@�N[{m~{�}jc:����� slG7�g�v)��O��;���}{�Ri[�ٺg[�~���\Y�'��ŕ�c����/���� �:@d�{��6���N%��C��a/�8�l>r�|OX\�e�G����K�!s�o�7��Zo4��s�[�_5ݒ��y��3�9���w x "���U�z(]�g�$� �<�0�lu}��s{׷-��{��*w���hܾ�Q���Rߙ}~�S��_Zw��.x�17 x '�����>�`o�T��`�D멞C�m�\���o�=z��o�X��m�l����kIq�����t�տ���$ ���E �^vƅ�W���|c2�� {і�f���t�,������/Y]���ԹsK�~����A�c����ͅ����{��;�7]��O� {ѩ�]���F咩������	a�t��ۊ>��n.K�×�G,+zg�o�0[�w{�1�K�$$[�����?��/�|�Y'� :�^���/?rK���gCn,@$��ܚ�@�O�U�:�l}��ٙ{�n�O���i�:�����e��܇��/ 0�:�^p�9_��l���Y9@D6L��9��1V�e�88W�S�����;����,�ZZZ٬�œϹ�}��q� 5�0�N���߿9�����08�a��
��ü�C"�s�?s@�rԾ����޺����*�F�_�����N9��r�/��o CˋC�y�����M���t�'����wG�֩Vk��E��ZH�c��T��O�x��3��m��)�{��6W}��s�Y}���D `(E��`P�y捅�����t���\�>����P��ʳW��>;s��z#�v���Uy�����O;�C���7_�Ar��kސ�5�V�6L4��XV,��������J�����w�4�l���f��l�Mkοa�3�����6��"��л���E�ѿ�JJ��#�;z�����ܽ����_��1;��o�wӺ��p�7�󬳞] �0GN9��e�K�f:)�
�G�����l�5Z̲�z׳�^�/�(�����k��i�����n\5����5:�� ��� sळ������KkIqy�>�a��I�g�(�X��_�Z�퍾�	�Xv�#ϻ��/�q�����S��
 4�����?/;hb���=
K�����!K
�Ї��4{�!Ց�w4��[�M��{��dZ9��������eo�ܯ�% 0�:��������K��(@[����V-���Y��u�gfn\_����ӧ����~��s��֋>x�� �@� {���\�����Hr#�܎�v{��i��I�X�%��+��C��o�=3�y���ג��?��N=��^��c ���Һk��!]~A#d✁�q��Z���ׁ��E�\��g����}����~]M���}B~�߼�/.�g�����"����~�ۇ=���e=d�����E!�#C��]��qwmz�t�/W�{�'�־�K�����[ C�<���e�7��?_O�Ð(瓤����a^v�ƉVߟC4�w����|����������z�7n	~����� �C�<E�{�w�]:�����%!y��r�ˋ��cj�����7��M��V�����q��v?��ڷ\^� ���Ω��F��&�O%���m��)g��/��D:� � O�ik/_�>]򷵤�"���/Y]*W
ٮ�ȯ8�Z���;'{������y��\>��m��޲�\�矵`�wO����l�>3�V�,\���<��_8�g� }M�<I���v�t�kii�0�F�Iz��rﺪ���|�WR�~񇓓����l�D�5ȁ�S�%��ܲq�~͏fj��)=��>���v^��K/}�֬��s� <L�<	�����Ƭ�7�Iy�0�+�ݿR��������,�Fz�+�ON�%��zh��|^������������ˊ�%�,�ڝ������=]������ }K��3;������٩�rp`�B��tu��ߢ���� ��r��?��҃�@���;&]Z�<^(,(fY`�������퍾��#[|�;�}�O��}��� @_� ���u7|jG���0�YR���\��v(س�K�k�����ο�� �����=�W��3����Aka �v���j�{��^���L?mٚ.}��k�}��ӏ�x ��t��������-٢À�Vr��r��ŧ�����O̶۽���@�0�jn�{�Y�����P8��9����A���~��Ri���_�{��h����Nh'���_=��߼����� }E�<�w�{�[�f�Nj�H.;��J�ZL����$	�q?��>Y��>j�N������곇���YQ,����zq����Hv���S�r.���ٖ���'}�k^�W�k �ot����O^q̶����}U>p��ۛ|�>��Q+KŰ���ɮ���p��d��iW0OCo��m���ۻ����[Q*�U��z}�������ё��]"�4W��������.��W� ��`O:u�o��ҧ��;f�|����Je��=z}�X%�wp���;���p��~߽�Ѹ���Q>��U�� ��sIz�a#ի�˼��NnQ�x��θ���}��#� �� ��w���t�s�![��j.{e7���tN�i��B��}ۥ�=8c���zo����Go���W��s��6�zG9~�J��O�����ZR^}�L��o���7�# ~���]���u7]\KK���e������9��}Ծ���Z�u׶����=��oi���ڬ?ky�x�>�R.K�~��#��F�iz����>�*2��>w��C?�}�� @�:��s��k�d*���a�di^��|�xa^���"�g�T&�S����V�X�����޵��8zU����wB�_�vȒB����wզZ}P��ұ7��3���Ͼ�E� DK����?u��M�eo�w���U��G���5?͒�U��_�ejb��v$}�M5:��==}��z��f� �O�����ӑ�cj�7�>�,	Ɇ���y����೧��� @�:���Һk��P���AX�{D�����\�K�T���~�A��n��lit��O4���ɉ#�)���O��&����x5�;��/w?�c#����m��O[{���~� @t:@�^_�}�|A#d�0 X����7O��ߥ#����_�\~��t�����������hyq���e��8���ȗo�����%�e۲�_t��B  :}�`O����`���=gE���U�R�d7�����Z��;��Ƕu?'������S,�Oy·Υ�,��#^I�9ێ:ҷ'#��y����?p�� �"Ё�����;[�ї��v�����×����E�ʥ��V��M���7�M��=8;���V�g*WF��{6�Z���>R��-�S��#}ka�/�r�U7\��/�� @4:0�N=���lH��'�4I�+�TV/�B�zg�_~P���LNn��Lv�l�j�����ɗP)0���������#�#_�ujrG�+��,�V\�'����.��W� ��@�ֻ���E[J��q��j߮�="���ՇT+�,��C�z�`h��ś'&��zͼk�;���55���b�E����:@�7�u�WG�tk����In��h�Ϝ��pV�D�q�����kgCn,�����[�c}����ʃ��/�69Ֆ�<�n��o�l�^}p���6��Ñ>R���'�7�V�����;ݧΣD�/^��i'�w��6��/}��O��v#���^>����R����Z�G�e����-��8�R]1����+�7�z�~��ɨw�l͍��=k���_�~̕���/��<o���-����F�q��#F��:T��bo�wo�4���E�?�6=�3��ˇ,)D7�pw��<{�!�^�O5�!�Ho�i�9]�gg\x�q=�ȩ �^#Ё��K/�fw�>���J��������V�Ŵ/��/ޯ\�1�j?����(zw���ڶ��I�&�N�s���\�w�+�OO�"=�1
K�X��� {�@�J��?ڞ+�خ8?�煴����~�A����<��k������5;��_���}�m��<�R��S��^ؚ.~���{ͅ���� �^!Ё��O|��۲�o}���n����GS�%��V������� ����F�ޞz���j�F��g�[����R�2��IH�dK������@ `�	t`(�r�W�;����N��J�r>IN8l�o�Z?��9�WR����S&��z�!�|���	�V��7wB�9li��c������ld"���ݧo �;�����2��C���������۴�'c����+˥��_�	�86M5[�x���k�v���H��i����h�M�����tq��Y �Wx�Y{��<���.��B�$'Z�8�sV�[gZ��V� ��w��o��|��#��Aw/?�R��ujr�t�"�#�����������y�� ����@�Mmߺs��uk{�$��C���J�/?�'�.?��21Ӟ�0g���3�v/�O�Fz��"=˒�7���o�99Y�D7 ��d����G�OO ���lˁ�?](�
}�7�U*�Gs�0D�$$�!`_�a7\��y\�H���'�N<l��Τ�V�{��7�$�wG��l��:��}��~! 0/:0��s޷��Pa�Ч^��\^�8_C�����K����qm�n��r��������t���\�����55"�	�d[q�o�q��_��GN �@����Bҗ��G�[,>cY��Xo[��X-_�������1~��#մ��I?`,_x�d�u��zt��gCn����ݧ� �sH'���_ߔV}�������-�D���r�L�u݃�����`������T�tBE������ڭ'��������񉯿�/��_ �)����������>���j|@���\z����ΙV�έ&���z�'�b2s��r9��$�Mv/W���z;���ڡ�N�W���.��e_X���F�9$Ё��#Y���4W
}��uH����ڹ��d�re�Lk�w�8�����E�,=dI�����Y����/�65َlM--�[�z��u�� �3(����lM�l�X.	��\�@����:�R��-��F��~s�+���V[PJ�e#��y�35�j�[�3V�e1ޏ�3��=�����^��6 �D�|��3���ێ��K�����Z��W\�~鶩�V[���ڝN��{�#��ϝ�Ύ�V��#dK���:�nm�l�fZq��TY��-����� sB���W�wcZ9$��g/+/�ujO�ґ\�����wOGw%�����;���p��H����t���s��S���n�o��؍�~�>pG���'��Ͽ�W^�� �'Ё��K�.߾sY�]����zӛ���fƖ�f�WR�-ӭ�w���du�2׿V���l�魈wC���Vk�z�~�ӗ-���I�fJ�~���� {�@[��l>�8��J!M^y�H%ILl�^��R�1�i�hG#�+���7��{o��w��΋��E۵M�����w�a�L+�>����y�^�� �%Ё�w��_�k~�χ>�+���T��$����"9�j�7��1��(�����ڒ�,-fOv�Cg��no���[���S��+ܙ_zƙg���g���z `��@ߛ]��[!�딎ܧTZ1����|�WR��͍C]J�F;t���6�sG��<֮�A;/>�f��[W�����? �1�k'}�k/ؒ-zq?]���h.w��R_�����,[�0��՝ݱi�ٺ�������a8/>�&r��<m�<���w ���������k�JY����]ê�;�f�����<�S�����~f��-��a9/>�Ꝭ��~���� ����_<�cHF��H��r!�7b�nu:7o��~���ن�N��v�3F��9;�coz�'/;�s�r�� ��&Ё�5Q����&�:�/�8���ݹkK���k3S�1h&Y�^\�[E�� ��&Ё�t��M�ȳB�N�'�KVW�w���h4��o����j *;�Eo8�ܫ����tc �i�@_�*��V'��b���A���j�7u<�4Z�����gn�T���qj��X�U�[�� O�@�Ω�\���قC�e��ˊ��T{����h\}�tm�vv���l�kO^��}.>�� �2������Y=�����ʁ�V���ݵ��@_h���H�n�� O�@����^�ƍI���'�ݿR�璾x3!wo�ׯ��V3����l���=��U�9�� ������X߬�<V��(ok�n�]������`��l �R+$��aQo��� O�@����\�I���
Y��x����a[�ٺ����3mg͡�M�_s�_Zp�Y'� <i���ҏ�˽�/\Y*���O������Lך�`K;�f�U����s�� <i�'������ʋB�d��ˊ��cj�:�n�O�g���o���?�5� ��"Ё��Z0vF;I����[��~�����J��Л��/wLMm�jz�h6��m��]ݧ�+ �D�b�w�q[n����PX>����1l�n5�����)w��@��-�� ��4/"���]��FȢ��KB��}�����o{�qŝ��Λ���N+��o������� �m�ڙ�N��������O�X)d�=�[7��^}_���axԊ��� ���D��O�ԙ¾�!r�|�>{y��)I�k�a�Í�� ��t�9����G|�W_qK `�t jS���}�+˥,K��i�+ݺ�.�a�C'���������"Ёh���ʃ7�#��ȏ,����%�|�'����9��l��N[{m��ӏv�"�n�@�f������=��pV���	���5�s 4Bnt��Z�}zq �		t Jo���ljb�+C�Vs���
�����O/�/�sj����x�t~A晴@��R~�o/�C�^��X�X=D�kwLN߻�)΁3�T��;�t��?sg �q	t J3����[^�r�.�;{���;s.΁�wTi�S:���� �K��9�_9pSRyV��Q+K�U���=X�1�x,٢��t~��$i �@��(����
.��p�,[� ��y�m���=8; C#�/����}����$Ё�L�"w�>����!ܻ�Q����Z x�ܢ��@x\��ɟ�ƫ6��X�آR��8�������wMO�`�Lf#�=��/-���w �@���/X"������^���_�kz�ݑ���i�$�Y1����u�G%Ё�L�#/+����POn�u��ݵ�ZC�O�L6�sA�<&�D�?}�[��Q�_"�̥�b�������h6��T˪�z��]��y�� � ЁhL�+oY�V�-�×a�ݽ�^�y��Ԁ����l�pr��9��@�Q8��I��ந��2�/��I�׿ͥm�f����<=���k�@xT���~�u��BĞ1ī��V���;������9�LuJ�<m��K�?�� ?E�Q���%Dl��ec�lh�f~��Zm�l� ��v�f�a�w'�' ?eh_l��mo��w�(D�ˆw�|�D�q�s��4�Tz��:��#Ё��s���Fy���|��2��N�wM��k��ZR9���~��#� �F�{]�0���C��\���j��_��ltlm���4��SSo�>�| ��t`���娷�w}(W���^oܱ�� s��U^:�O��^uʹ_Y�))�
�ZXL�e#�lضx���_uom: ̑Z:zd �t`�ʏ��B�w��Vϻq>t�ۯ{�6Skt��}	`�$��_����_�r� �t`��	��B���Ð�1�j�pSc6 ̱�b�M�:��	t`��]�v�w=+Djy5ˍ�,�o�W��-�󠑎 �7�kn�ؿ�l}�a�^�v�xa�V���֨?��� �`*)v��_�^�'�n t`/JF�O��:�Qn����t����L �'���;##��6�*  Ё�g&)� D�7��RȢ^7~��>;Qo���W�l�A��"Ё���3o,|;)��:`q~��>�]�v����yW����"�o�+��g��Za4�-��@���?�T��i�̿Z���9t���P �I��!Rc�,�ҡ���lY=��v����g�O� ��@��zR~^���E����x�F�����ȕ^:�@����tp����3���9�zRzn @���=�}��'�(�?/dI�l$?4��o�zD`:)|f����$n� ��@�]#�{u�Ԫ�\��}�u��sӦY���^�L����Ƒݧ� CL��n��a��ʅ�3���m��t�m��B'W�݇.Ё�64/D�x4�ʡ!R+F����x˦�z ��lVzA rC�B�C��MIqY�-�V�I:Z̆�����V롉f3 D���
 CN��Y,��:i��0mo����-`�͆⒏��N<�l`h͋Q i����#�q�y�j��7� "�$dߺ�����k����@<ZY����ñ���m�z��j5 B�j��@��@�U=�"T�'ɂb�C�޹��9�VRxf b�W���o�вJ������>���Oĩ�����@�ͻ>v���!��-����{�7n>bUO�|`�t`�$�/	�Z62$�Ϸ��ī�FO9��e}�����i&������Ur趷��v�	�ޛ�_ CH���	)�i>Q�;'���vV꽙+Ё�$Ёy�L
+B��+ñ���m���k%�`H	t`��;�x�s҇!�ۭNg�d��v z���< )�̋�\zu�Ɲ�j���J:���q��l���f�[ ��@������C��g|q9���MX=��l�_ ��@�E��<#D�N�&I-~�?��!Ё��
I�Uk�����hv�C��vmo�reOi�:�MS�V ��V���:0t:0/:�����t�W�{w��;Ο������� 0d:0/ZI�O�Т�pz �#�;  !�̋f�_"��4���7����vV\ ��@�E3�9�w�0�+�[:�gInE B�so���l�ά"T)$���V{�� :�_Z![ ��@�\a��e�\|��{P57�+�[km��@��d�(���k�{��O�_mʅ4I�$�7��m��?�NV C(���IC�ܫ�t�ϟל?�O+$ŏ\zu���[ CD�s.IQNp�擁�-�M����O��ܽ+ �̹vȖ�s������s�� }�P��&�t`�t`�u��X�P��t���N� w�O�C�Uk�����k�tQ�P1z�{����+-��!#Ё9�N�(�<�[�'-��@�ju:Q�/�K�s�$?"4�gЭ�}-��Q sI�s��	�a
�����zK��+u:0|:0纕��ea��m�;п:� ��@�\'I��B6�3��t�k@�jE��.�\����t��D�V��-��V����$�:�s�4��kM>	�-;܁~�f:Q�hK'Ĺ�=˒�^bn�;���>�S���0����t�	���������-������vb|�>���wi��9п:��@��@�\����,��>�=�ٶ�����T`���̹v'�.Ї`��:��ډ@��/|��KBt�g��m�ہ>�	Itǣ �@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t ��Ъ�;�N�7?�$I�Y�X <� �:�V6�c�ҽ�1���Lelņ ���  �!W�N盍퍩� �1� �8�#�vtZͬ935 `	t �'PZ0�m��̷��  sD� <�$�-�4����V� `t �ݐ�i��x���-��v `�  �)�r��ek�֯��a �=H��N'i�N���P�MҬ5?�V�^Z�d�޾~��#�T�>[�ٱiI���`Y�<ջm>Mׯ0:� ����j��/��2�|�V^�l����]���&�H��JgjS�F�i�/�gʋ�mڛ��� ؓ:��h5����t%�Hs��޵g�������5 � ���:�dvz��l5�5g($i�譜��=p� {�@�c�F#W�M�V͝5g8$i��xņ��ؾ�\��� ���lm��l�m�ex����\.�8Į������S$��L���z��:�N`X$I��B����N��ֶmX&�x::@i���3�E3l:��P����|א�v� ���z03=Yi���1t:��K7e��l�Q���V�Mp`O� �s}ì�`|s�T����K��z1 � �b��4�\ad�|yd:D��}�Vc� ���w'�����g�S{�]z�����E�I�k^u��'��,fИ��Q3
�fU�q���M4Ƙu�5�d�q��;�
B�i���]j�:�3��b��roU=�����*���Kso��ճm ��i�u^yn�+�:b�~��b�� �T: ���0�r�Zӫ�[b(��:���  ��t 0ǧ�I���W�b(��6��5 `t 0 ǧ"�W��[V�PA�Y{��  0": Lǧ�ٹ��8�mY�;��X  F�@�	y��4�4�a�ٮ��/�e)1P4���- ��� 0n�<�vsA��8���As�8 �� c��i�wY��8�l;�� ?h,m~^ cB���p|pˎK;�8wb1P�^�8 �� #��i��XVR��~�r�H�D�;�s~f cF��q|�(:��tr^(�o���n��
 ��#�`D�n��Fp��P���C���@����ځ��\ &�  �D%L��k�n�8�ǹJb�T L�  FΫ̯��R_L���o,mM��M E� ����sk^���8_K�<��+ 0q:  �\���*����X����  `   ��[(�󕹦j�\^��AI  0�  6��/u
�-�b(��:� � :  �T�W�綮���N���5 �0:  �4v.?(�m[C�f5�6�  �  `Sخ��/�e)1P�NcA  0�  6̲��hr�z�Ake�  `0  l��D�ŝ-�N�@��/���
  �#� ����4�=�s'�� �p�[ ��t  pj,+)�m[��\$�� �o,m�l  t  p*��s��b�$
������9  Kt  p�T�����|1�Jb�7���  2�@  '�P߲�J}1�J����$1�8 ����  �0�2���=1�0�W�oWI�  2�@  '�+ϭy�ZGL���o,mUq�	  E� ��ʕjM�Ro��t��-mMB�   d�  W�Xi��1T�yh1E  �t  pLN����W�P���B��� � � �Q9�B�Xߺ"���ksѠ[  ��  �v=�8��X���F=�� �!� ���7(�o_25΃n�v�s ��!� �#,�	K;�,�N�@a�]:� `
�  �0ˎ��y�(�~{uQ  �R:  H��J�8?h��H�� yhk��  �� ���q>�����B1P�q �:  �M�-9^>%Q��K�D)[  �r:  �K�[9^�%Q��V��8 � � �Q��[(��@*���ځ��9 `��  � �2��+U�b �$v��4�s �!� �1�r���m1�R���$
= `��  ̐\���W�b�a�/mM� /  �  ���K�|maM�o,m��AQ  �Q:  3��
����1T�qh1% `��  L9;��-�����|��* ��#� �b������KbYJ����~�&  �@ `ZY���۬��V]  �� �4�����cɲ�D����X  � �ic�qi~�A�vb1P4����  ߃@ `�XVRL��vs�(���As�8 �(t  ��r���(�T�$�e�bٶ�k�m�:�x��`�4���-  �A� 0T�a%E�|}ב>���n�N�8N����}��F��Ł���s  � �Pn�i�npܿ/I,}ӏc	����mw�����S��$
�a�+e  8& ��SN�%��o�SVE�x�u�>뎛Kt�;���%��[;�=}�  x\:  ��|[�\\�/�w;�����i��]Ǻ��{�$voe�vIb�7  8�` �Q��:i��� ����rK,+�͋Jr  N� @)���u�@JT��9� ��C� �1i��-��PV8�[*�  � �Q��q�SE:��  ��F� �ʲ�b(�k��  N	� @Xv��8��PѠ��yQ  �)#� 0���H�Қ�D���l%QI  ���  L�K��&��yX��"  `�t  �y"�Қ������`�~M  �� � 0�J�W^ˊ�DI��pPO�>  ��@ �0:�U��f��RI�Ya�n�  l*  ���n���T��8���s  6� �A��oY���T�Zq ���  B9��ع��H)G��|Z�  �� � 0�r��4��b$e�  �� ��);�M�'R*��h�ƹr  �� �%�ӷ�|G�DYv4��k�  �/�  L��݁�Zb(�[{�9  cA� 0ʲqM1�>JM%�  ��!� 3%V8<�\ꖊ�  Ɗ@ `����4��,��Ȋ��$QA  ���  ��+��\"�"IX  0:  c�y"^iU�J�DqP���,  `bt  Fl繲�q�8�  �( �R)��kbY��(	V��  L� ���8��nّ�(���b��<  3�@ `TrŦe��H%�gG�9  &!� ��b��H%q�
�si�S�  �@ `�%�׶��@L�׊�sq �qt  6�r���x=1�R������m  �!� �$�v{�x]1���s  �F� ��\_�|[�DYV�O�\9  �E���(��P��q��8��8�k�  �k ǖ$	�p̀4�b��n�*�	2+�#;�"�q�D  S�@�ͤ�D酴�	��e�*�sc߉I��R�'�4�>���M/�/D�R9 ��"�`��Q�0�D����ͣ,;J�|����Ѡn�8/��?p�(t
�J�h: L' 6A�vȨ��Pb�bp�[�_�$*�NǖM�
�(_,1� S�@��PJ� p֛ό��ɕ��6s3�+��E�T}7�#�X���m�F ��� p���>{�^��Ĳb1������e�L�3w��������o N
� ��)�Gǹʕ�,�6sZq�8�f�J��i1� �� 'A��Li�Ej�[��b�$,X�_�,=�=�B�T�2� 2�@�Ĕ�٥�BӲ�@L�Dy+�낙�D�p�{1�tvy�l"����V��`�('����@*�sVد��{F8LOy�ץ��\�`�^	 �c#��8�0�#֛Ϥ��ږ�닉T�Zao޲�s<֠���ql��κt � ��#�f�r���x=1�R��8���bc]: d� G�z���z�x]1���q.¬�#��+��q" G����8�����3J��@�|[���y�[�D�����.]o�y� `6 ���q�3KY�/n�)R�Wg��9!�q*������������������ � �fp�-��@rņHǹ��\%96@o����K�o+�|s��e/x��n��;^�^�@��LI�[VlY��5�j8U��pSXb)�zmS7�� ��(��b%���	}W)%Y��=v�֭�����߼�����K `�� f����8n�#n��J��C793�~W��o��Qo��6�N�]�;��i�r%��Nپ�;�O�~�����^~@ `�� f��5 �+|'Q�U��1\ǝ����v�7n���4~� N�`&�R�����px[�Z7>җ�m�/����L�/ 0�t 3G9��urIR �̼��ҳ��Z���s������+�/ 0�t 3exp���I��� `e&�-K��~ޯ��w��#���
 L��X�s}!*.�� p��H/�k�e��;9�����u������ �":��0��N�K��ܫN �0�n���t?Wu��_����4�4!�L=�(��� p\�H�<�ww_q�V���[��>|� �� �L�~���� N���}���L?'�n�u�^��k>���~� � �L5}��/4 pR�9�bY�P*;�<�l��������ο��^}� @�� �����& ������,K�Œ���e�ۭ��I� 2�@0��~�%�`�Aߵm[��X��n��ԫ����;_�� F��:�?p��  6Š��Y���\.CݩN��_������{�	 d� �JE��� ���w۹R�8���@��X�wj������� d�`j����  6�R֠��J��o�f�Z��-������>�T  �t SC�u�#]  #�ı���4����ծK^�_�u��� ��T�;�s�9 ��>�Ro�i����ʭ����]��Ȼ_�J_  Ct �ǎ� 0^����q������� �@�Eah�c; ��ސ�vs����ݭv^�K��O~����� @FpQ ��z�A�æp 0!�9�\��=q\��~U�6/ �:����l
 �����{�ʕP��n���U���߼��/ � @&����7* �D�=@ܜ���g�z���-���k�}���	 �@�9q�A���v 0Ġ�uˮ�X�m�z��-;w��M�+ `8@��DI��&�� z�Q/}n6u=��j�~�uo�O �@�)~�˺s 0�^�n����l��古� �@�zj;���������M<z�m�_�����m �"�dS��|��f��~�����X:�L��&�� ��S�C����vuo��?��w~�o���
 �@`���>�W ��~��G�����]�����_��g�V ��`<}|�  �C)����J��qSݻ�z��ƇӇ�( `.zMO���% �)q�Qzss�Dsw8��ko�񅌢0��Xz͹��v �,�a\�>�aznݽ��7}4}�| �p��Xi�;l ٥��M�0�`�g C�0R�����( �8S7�ӣ��?��/���� ��/ #��.g��4PJ/Wr
��q����SzG�0��8zS!���  ������;�c�(���X|��������� �t ��=�� `���[�TC1���U���\0�=�X5 �>Q8qŎ�u��!g��/������]�i�	#���s �^zGwǭ�eˡ��G�ó &�a �`� �[�N�P�L[��/Y8㗯|{�Ϯ��+ 0A: c0z �/�]�\1j-z��vl} }��	�b�=�٠G���Rdڹ���O	 L������ f����F���-�_z����' &�b ǱŹ� 0;LEW�%K�w}��@01:��ӻ�
 `�Da`��X�?�c'w E��8}6�  f�?軦���:/x�;^�w�� &�@0Qz�\%�% �������n.gԹ�Ka����`"t >�� 0���5��@?��� L�`b�(�h5 �a&n�%��W]���~�[ ƌ@01l ���F�E_
���;��� &&�8Z f��(Դ@_U�� @���1�� �R�8�-�q����s��/]������_�	�1"�LD��p �����X���H#r^�>"���`"�� X�_�b���d�1#���� G�����I��7���~����7}M `Lt c��� ��a�n��Zw�t�M�J `Lt c�w�  �`�n�l�1"���ީ��� �G;<�]�e����� ��`�6� CG�k�1Dˮ_�w����W� c@�+�A�  pq�nΜ@���u������� ƀ@0VztD  8
�[kE��@0&:���>FG  8
�[k%�Y cB��$��s ��қ��z'�W Ƅ@06�? �i���N%��W���g�_� 1�ذ� p<��V$�+q����� ��`,�ٶ�? O�ƽVt맅@0:��H�ب ��������ۉ� ƀ@0l 8Q�a��}�� ��`,b�, ���n��1 ��E�q ����6��}��53�����X(6� ��8�g���9����|���ݫ�- 0B:�� � 'j��a;b�A��LzG�)��� ��q�uì@�i #F���@ �$�����j� ��� FN� ����Y�Al- ��`�L�� �O)%&�,�" 0b:��3�<[ ��L[$vQ `�t #�w ��2n]\O `�t   Ǵ@��	 ��`�ҋ,F� 'ǰ׎ز��z L'�ș6
 ��J�`�t   Ǵ7w�e� F�@0r�7�� �]JA0z:   p�8 �F���X��J�}>�����J,�?�Ob9�,�2��,"�����)�����6�R�V������ `
��)�la� p2� f�`��Y�\f N����!����� �>�,A0:��S��  N� f�`�� �ś� f�`䆛� pG�A:��Sql[9 ���Ĭc�X�`t #�$��  '.�#� Ɓ@0rI� ��G#� f�`��0t�� 8i�S� f�`�(4j `�$��
tF���`�8&� 'L%1ר fO~ F.��� 8qi��u	#� Ɓ@0I�l� ������Kt �@���� �G!ר fO~ �"
}�� ��o�5*�� �Ũ'? �+�}7_  �+
C���@0.:��H/��� p\*I3�XS �F����R�mYv"  C���@0.:����Yn~   C�f��N���D��y: �q���S 3�'@ c�9�T  �%}�0���� ��QO� �[�%*�Ա�( x�$
�J��A�'���.�u�/  <J���b�� �C��(�= p�?0s�8 �X���:t ���Pb���� �*���Y� x4�ן����N:���8I��\�/  <,�{1̑��M0:��z�B�N� �k��zb���� Ʈ���
��� ��8��(4���s �@�;�� ��E1�`t �4w �:��s�9�I �L���^�/
 `��Q`��v�t �@��=�=E���l��^&��s��q �L���KLs����t21��u �@���~��j�Nz� `�DA�Ǒq���s �B�����.{�ZK  3g�i��0���$�D�ڭ|� �-*�]�w�0���$�D驍l �GϠ� &�@0qz�cy�@�Y�k������ &�@0q�~�)��e;�  �^���IWÎs���`t F��b}qM  S��nw���:�I#���m�
�9ײ�H  S+���0��[�}���X�9�1�^����5 0�z�qG�i�7�]��>0z: ct�M/_�;bY�  �N�&�����vK�Q#�Co�����|y�) ���o7�<Z�x��Z���9�Q��f>_���C 0E��/����s�DF��`�t F��w�5֢�t�6�*b��m�ε��� ��i5<�T�\t ���sSG�Odz��J��( F�@`�^k�Z�ۺ* �LS��Nc�ȝ�Ot�\�ي7����H�^�-Vj�� �YA�U������'�DGχ�ľ ��� ��i�Vj[v� �Q*I�n�Q��蹖��� ��� �������|�+ ����jz�O����Y1ˮ ���h����b�c�  [�(�����dG�5�N ���hI[��j�X_\ @ft+U1ԩzޖ; F�@`<=�/W�0 2��6kz��Hǹe���u���9�#�dB{u�Z�~���� ���8ʙ�1�v�k�5K%��� �� �(��v����5 `�nc�n��p�2�]+H�ﺗ� F�@��V�����8� ����9�];��s�(A  0:�Li��U��\��2sx f����n��P��Z�9b�X� 2%+�4�� �1yj���T��ke;�O `t �����^��x���Ncn���+��W ƀ@�I�ե���=�XV, ����~Q�q*�ң�r�ڑ
V�� c@�Ȥ$I��zp���cY  ���i�.W�`=�+?yߵ��E�1 �d��N�Zu�Tk
 `캍CsIolxz�t�ot��n: cB�ȴvc5�������N��� �E�A�����n���� Ƅ@�i�͗��E���*��i� 0rq0(�7H�`�ھ��l`lt �v������]K�͝��[�{�  FF�w�\9h��s=r�ѩ횕��T�� �	� ��ʞ����5b�$�S���F�[���� F@��n��S/)�a�Y����y�� �	� �.:}A�"�����3�s�0��Z�8 ���Z����M�͊sm��� #@&r�\�����H���Uk�������C< �1��ڜ?�o|׵ڬ���j��Y�1"�dғ��Iε�z�%~����*��F'�� ���n���6sj���/�\�; cD��'��'�?���"/�A�9�ϩO����	� �*�{���JQ��q�դ�����) 0F:��9wgM*����a�I^s�ҏ=��>sG�K���K"��\Y*��t�o��vm17xP `�t �s�'��)���Ÿ�������j p(�7�����s}�l�^�? ƌ@�){˲�Z8�a�$I�3+QMΪ����� p\���ơ�ue�6���|������$ 0f:�L��GϏ��H?�nׂ����m 86����9��=6G��v��v�K_�, 0f:�̘/{rƖS[
F�}�B�Ǖ���� p*��4���82��sm���m��$ 0:�̸d�l�j,C�I[ܺ�J�[���  �����|�����֝k�JT%
_' 0:�L(z�����ᏣG�u��V�) �!=r�<�?#�Zw�n��^{��l� �� 2�){����o�(���z���毰���Ҵv�uG{��=��� ��� ����Ii�o&�N�T��z 3J�֮7�#����k�u� ��� �w������_<Fql�H/��}eY��)*�3��n�V��|��/~@ `Bt F��b���j'*N#��i˕�@,; �I��Բp��6�ۏ�3��� D�0Z�����7�ϑ$��i�
i����� S,����JV�|�;�����	{��u�	"�����7��^t�������Vw=�7 �Ba�]m��%#F�c��v�ڷ]��� &�@0rz�c#s��^j�?�r8ҭ�q�cI�N;_*W�F�qN:���Z�vc� ���G�)�#�K)Yp�� �0���я8�R��Ǹ�`[�閇��O�5�H�zݎW*�,�� �DY���\���IF�3εmv��'���g &�@0�B+��E��Z�#מ������~/�ő](��X�	 G���Y=8���/��D�sm�|T � :��ٌH�����Q<�����H#='��R�R�6 ���0�\>X��1j���%	���y���- G�+=�]G�FܳԑO}c�<��Ӕ�6��$���f��dI��ʭ�C��Ծng�?��֭�=����t c���p��~�rG>���/٣r�h#]��a+K!���.����j^2fq�X�{�/ �@0v���V{�H��Kv�|��U�^��Ob;_(�.�q�J��ڡ���zsmq���5��+n 0�`"6+�Z��_�>�Oݣ*��ȯ�|�wү�T*Wb�9= 6M���ʡj�֛k��sW��Q�� �At �Y�����/�t��̥{Ԗja�Wyq[�V��Fz`s^:�	����G�T�k����yߛ~� !�L�fEz׏��r�p�����ȯ���n��y��S`�;�I�G��-�gqJ�6�8wT"���� �!�L��@��r>�m��w_�_~��;����c��|߉ðT,W�������\>X��.��&��n���W_�Y �� ���ǉ���Czڻz�9[eW��(�n�U(K���l^.�%�
:�z���$�&�v����f�L �@: �lF���k��H�ʳ��s�g�?���=�N�X(ˢ�l�$
���C�(
3�����i�N�������I M�Y e3"]��@K:�P�{�nUλc���Ў�F��t �e8j�m�:�F��6_gJ�;*Q{J>;�0��)�(�\ǒ$;�l�/��=��/>M�+�%�M�P*���T�8̷V�2;j�������7?p�K># `(3�-�(��o4��������٪.=sql�a�Q�Yd4�ɚ�QsͶ�G��'-��x�|�9 #�M_���=���R�;����=��2�u��� N���B{u��AfG�5���������\�_ �`: ��<�=+]�����t|y�E��z��hz�j�B��97�c�$q�Z���Iƙ�5������~N� 0� ��0��nw�5����=���T�쬍u�����K�R9t�\( ���jkm���s͏4�cԎ��R�^�����wy`�t ��雱�{%��W���]�]���d����v�\.��%��3L��i�T��7g����ܑvX͵��%� � �E�8�`���i���ol��6d�5�g?�45W��:�s�H�f�P,F9��g��	Sj8���ie~:�f�fpGr�X�Yjs��� �d�|%/�z��Ϸ�7��t������٪.:ca�������z껞��P�I��rTR�YbY*V�@�&�o�;�i�ή����H�V>�u/�� @F� 2+�s���d�������;wj?UQ���n?(�-wԳ��KJyw���>�ݱ�\�Xb}:NN�����̐DIK.3�>�����k+�8��Z��&�7_7/���~����o�* �:�LK/����U�׋��7?(�`cǱݷ���?�;�[+c�ꌓ�����lb�>ȸ$���je֙��Q�~��Qr^�����L6��):��p��������>���@������#����svԆg��z3�>=l6�^>�E_Y�t̅f�J"��X����y��7����Gz��z��t� 2�@05jE�z��U7~k�|��Ɔ?ޝZ��ZO~���mՉ�路��yq�X
Q̧�8�o�U����]g�<�}]M��S��~�� �g�^8 �6׶��x�irƖ��L�pcS޻~$��ƃr�is�G��&�Fӵ ��V$�sMs��>�}���\Xi]{��/� d�Խ� �v�κ�c����e�jo����r�rG�q�6u���ĮP�C=���y��F�S�{��ʠם��,Li_wvn�;���� Ȩ�|! �V�Y������V���9(q����k��ǭ����.�!���˄��路�u/_ĲQ�H����ά%�/�v�^�ml�SeaJ��y���хs��	��"�L5���%{e�|I���J�l�c�{�#�z�\�wA}�Y[Ķ�I�z����P,��؜~ �˱m9�nU�����Ç?��P��ǯݳ"�BG���pU��2�W>}:�)03��� ��^�~�g���A�#���M��]�r�R[~�j�|i�CLA���8�����'�#�i����',؅b����w�F����&������$��=�EOg��l�����_���}R  �t 3#��֏]�Sv/�Ӌ����6j����~�>9g{M=�mR)�&�q�Q�-+�甼�֤}�J?JKՁS�Xv�s���sN�=�l��vխ�����M�3[gܲ6j�n����o�� S {�� �AO�Q��,������|k_C6ڮ����@K�>�N{���E=v������ ޶]����F��T�����Q��q��Sw��.8��e[�v�?�����ܫ>�ã�"���ZU�2�~�)A��Iz�곞|��ڜ��o>�)�]���o�ߒ���U=a{U&���RJl	ݳ�R;����o�r�J�<��'2���Ӌ�f�(�4Wt����޺��]�k�s�9O٥��
�צ�<�%��暣������w�K� L�l>#�&ٽP�M�?w.�7�]ݔ�f/�O߼O�׋���m����u*I�eKvU�� .�}�H�8�?�z��O�s[3ȱ-9c�-�=g��h��J���g.ʎ������`3��l������������%� �":���צ���;����h�j�ߔ�{���O?{[U���%ψPO�D�Wrμ%�.��v,�7y�1E<cF�{���Nyw��,���R�t���3����ZOL��s͏e��z������
 L �/��g��޽,_�{e8e}�t������s�#쪫���e��I%��,���=%y��=��,�|�1u�y�:k�)�Yw
UO���q5�$�����N���{W&�F��ή�<+�ˢ���'}J `�� p׶�|�6y����l�?�ܔ�'J��`c�>�){�ԥg.J�s��J�k�EEi���EO��ʽ+i�͛����cY{�n��9���l��K/�w#�Ŷ�VP����c?�mF͵�D��ϸ���� �B: E����s�n�p����lڴw=*��{W��~�rIz�rf]4�O�?kΖs��Eh�r�J_�~,��4�Ϙ��kvq{I���Ƽ�O�X��էnzP��p۴���D]Ti��o��[ �� �����p�[�_�/޹$�&m��?Η�Z���[���>����Q�Dq,E[��[.�R�Ձ���Xl����BO#?��vV�����Q�D����~�����ޑ��>-������ʇ>t�5�@ `��w5 �ql˺d��R��ms�6��X�r���tߪ<q���]����I"uO�>�����-K�Hj���1N��E��Z��Y���*V~� n�֣����$�"�H�C�^�����~4�y�_�ȵ�_. 0�̼
 �i�?y�9�������ou�vd��Qu���OJC]O�sb*�$�5�{jyQ���X�e���e�w}-f��ڲ������l�8�#����	i����P��[�Ϸ>�qTG�M�t�#����[_� 3�@���c�d��8S�_���~@�ۛ�>]��[�_�'��S�.��ZAL�c]�ۖ���Zp䩻�d��ȁv�F{(�����/��4Wtegݓ�UW��]��������,|W�Hݜ�<��A8�=t��۴Lg?���|����g��@���nw�`R��)s�����o�א�ciSG�t�ޱ�5��/���}^X*&���U͉Tl9oKQ,�"M_�j/����`3b:<���9����ֲ-�+9)8�7x�(;'
4������ᬘhD;�O�:�G[�:�9�|Ε/}z_ `F� F��-�s�zP�[��e�2��w��9;��{W���u�页�𶥚n(w�κ�N6֗&��W�JU��/�]�V�Ix���}M?:�
cF�gW����4�Ki�W\)�,�����D2�^�R����p̃�ݑ�w>�a���Apn�{�u/}�� �!���;��b���������P��k���c[O;{�<qϼ��]�r�k�>j����[�w�ǿɓ�[��I��]���r뮸��ϟ�)��j_��z*\����V�t�(KY��sr���m՜,�4�]����2��D���F����|���6~�t��Og�fE�������k^��C��w��W�����g|}����U��瞒�Z���ƺ���ƽ+�v4�:�������M���ޭyʞyٳX2~���$Ib��ϙˉ3W��=gU�=%�'v�$�r_��A�ԉ�^�S)��X>��E[��{[%G�IK����������M�9?Ҭ���O�#�Zo�������
 ̠��H`���7�/y���km���[��m5|���X?t�6����a�����:r�^jo�bn8�~�isR�g��]���~����I.��Λs������h_�+��k�(i"&�@�5TK��K��
���v���$9"\�X2��Cz����D����h�F�R�k������׼��W�� ����U�Lz��W��K�������_��TG������n�ou$��5��|��C�廖�������˙U4=���4Q�4����(���8��V��N��V �j/J�0�EI���P��w��Fx-����zd��G��z�x�k�z�\����Z#�>Ҭ���X]Zi��C�\�_ f�`��w���������}�Y��=�����:�/ٻ���w�8rI�~�������>�͗�2Mt��ǧ�^��-�%�-/e�n��^T��$�P⶟�M?�w_��^��~��~���Ǔwm�])�l�x��=+��4��8�sl�Jb��?�^��r灖ܶ�)�ڃ��YsM��_u��^��� �q:��x�^���Ho��n�F�k�������E��PS}��k��y��3�����ێzQ�KC���5������pC;��t��W9}�rZ�[\e��怕�#I#^E:�{���A�:i�u�X���r޵-����;�~��ǚ�]!�i��ӿ��mq��S��'�׏�t��Dݳ������]�	��+���8�����^}��	 �@09:�/�/�z{�#˛�!#׶�ǳ]���Yj7�{`�;�ϧ�����sPN�R�sw��̭Uɹ���>�w� ��#�zNA>'�|����5KY�+��W�m�8�=�*	�� �� Vj���a"���(Vi�+�>����輓�~ӧ�Yv��$��uޱ�k��ip���o����֧���&mɱ柧>k��>����-��@{�S�׭���b�k��ɥ��knx�eLk��� &�W_�������u���?C#���e�Y۪��Rk _�gy	���S��蠾����Z�s�X߻����������������C�ER�&�w棾;uTY���C�p�ZJ���X�)�:����~zu�G��X��X���Q|���s,K�ß[?��v�[9g8�m����_בm��m�i���,����e���{F=|����z�6<l=�u�ߵ�������u���Y�I�\Z]{�oz�	 �:���k�/{����v��:V1'3j[� Ϲh�<��Pn�wE���1�u��t������<��垰�*�/Vfjd�T� �a������!� oG���w����f�Y��#�&a�Q>��ˏ�Si����8��8�G!�ᆫ���K�O~���\KJ��0}\�>K���m������F:�]�#�z�^��Ⱥ>W��m��{��٥�E{`�{x�ȡ�pY�8����)H_\[�"��? �cp���}���eoy�%����5T� 3εm9wg}x����o��>�QuM���O�כ��/��-���Be�v��t����7�����W{���qc�cU�g��V�?��7]�� 8*�Qn��ۮ|���~}�q��dnN0������.?x�ֱ��kz���4p��_�X���p��^(GہI�S�4�r�3q���H�I��h��-���9������n �1� �s�U/\zŻ>�3p����݂G9��׎�E��DZ�p�怾���-ռ�Y,o�͗Ķ	�G���]��Joxڸv^?F����v�t/��+
 �q� ���W�{}8��?����pۥB�=F����@�Gf�جѣ�z�y}��=+������4��{��c3u�H��v��9��f?���3�G���=��3�g��/��0 �����/{����'��V��	�~T��j�mR�����v�=�iEϑsE�9W�]���z�v�0������F_V��D�����O����y��W���/� �0��>�����_���?������v)����X��x�S���w�^�lN˻N�:�J���4ؽ��O���P˗�;Ho�(��`|G�=����>�������[.�Y �@&|��^u�o��s���?��.���a���k��j�C�z��˝����'2W��u}�b5/���-�\����#6����>���#蟝�7�pr
&��~�C�^�f �4@f���+������_[�&R�
Nؑ#�&ĺ�?�Zj�v۾��ל���˞ښ���j�h�\FڳH�����4��a�/w���?�ݎe=�YW~�j��Ri���]�1j p�t ���+_�oW^��]���~��x��z�+�db��ӣ���mr8�u+U9�7�ӷE}_���]��v��f/�F/��a���F7n&h*��o��n������]}Ū  N� s����� �=�kn���=�?��[��Std�Lr��ǣ�N�o���u:�ki�ϥ�^/y2_��\)���K�������&Qᡬu�������ޛ4E��������Z_��k�� �a:����\��������_{�?���v;9FS7��̭�2tTY�����mu�����B��S�M���}��>���9B�=V��~3���"�~��� 2�͛�����$N.*���O�y�U �:�L����/z�{>w�W[���'�[^({\�o�#�F;2֕2�T�殯o?;�w+�U����0�K�+��+��^��o�4䳾Ӽ^>����"����hx��#���]��8{~4�1���ѩ[}�ɕ�����}R  ��@�y��e7���]����-g�s�ygm�d:�L����cݴ��'J���Az"Gy9���i�ӛ��[<��m����N��>JN�z���=<�]�?�����������ֱ�>m���w'`v�����I&�	!KX* ���j�Z�\�Jݪr+�,"Q�6�9g&��a��L�9�<�jY�����E�׺[[����[Y�,Yg;s���4�FdI`�y�9�����7	��?���_sh�7�F<in�V��C=�'�<~,kFx�]��o~�9o~��&��D��B�*�-���]��~�����I `F	t�-\�bE�>�S����m?a�sN8��E�S?@�2�H��z�?�f$��s��4�������Ծ�?�ɵg� 8 :�V�}�ك��Ư<����g��������Un�']�!Oá���g�n�ݏ�=�� �@���#����<_xۥ��u�1�|�)G/�]�A��g[�vf� OK�F��=�~��?��W���v (����,k�k��s>p��_~h��_>�����쫕=��G"]�w��oSw�zz憩���=|���[�� �� Ё�v��s.}O��o��w�I����^��GB�������w|�2��(����y;^�����F ��@��p��;�p�Y�\���G<��pDf��<�T��:\o}]y=?i���o����b �`�@Ǹ��V���͛����/����`�zhO�M��/��G�[��sxq��c����K��� ���@G�r��Ⱘ���>sג�o��ˊuъ�6�G<�{G��G�c�����}�< 0�:Бn��������s��ŷ<뤓������/Q�X���=oe�^���<K۷߳�����A�������p��?p�Uw.<���?kY��XP*b��ѱ�dW�g:���s���ٞ�;���Sz��O����/ R!Ё�w��s�{�~l�׿���N|�3�u�<���xt�
aZQs̣�������\����1 ��}�����q8�̵-���K�{��=�s��6�󱩓�?\�n��� $I�����r���W���՜�N���r�a��R)�ºB��0w�m�,�_����o $K�<ʕ+VL��e�^w��������O\t��"h9ˊ[8�w��W_|�W �� ��#�Ͻ5K����w.8�}�}�qs��vu y��D���;>r�ڳW Z�@x׎���o�<�����#O|���]���@�z�t�Ĺ۾�lQ���<��� -F��=���꿯����r�-�y�I'�0�["̲b���Ň�ZZ�v��#� hI`?|h��w��w��ᴯ��{���OX|��ӁY����Q�m[NX0u�GW��W��&�����>�/���K�z�=?\\}�3N�_�?G�͢|�؉�v^r�%�W mA�<W_|����G���_p���'3gA����/LL��7��O]|�9_ ��0�>���y�����s��Ɠ�;�k^OQ�3fw�����%�.}ˇV�i" �v:�ɲF�C���?���a��3N^���oN�P���0^_>w�[t��9@{� 3lO����o<�_�s�ǲC�x�P�W_>V_޻kO��Y�t �p��t���q8��͛W���{?ӽp�i'/?R�O�?�O-����M�u�+�� ����4o}��ˮ���eo=��es���L������;>���ۄ9@g� ɞ[��kg]z�%Y���sT���@�ZT�u��Y���w��� J�̂�.>�J���[���۾Y82,Zv\8ni(����7²�m�.�|�5��ݯK>; ��:�,ZX����w���4�,9>�xԒХԡ-��z��m?8b���W��ܯ ؋@H@oq:<#���?��-�B8ty8��¼�b Z_�������c�����~ �1t���<_| �m���7gYX���p���5uh-���f[��;�����]��r ��@H���x��a�;ÿ���-<&,_�8��vUR6/L֏���/�u7�u��y_���K� ��t��5o_�	���	wo��{��#�:&d�S�dB+�x訹��c��U7�~�t ��$�ZD�Ǐ��B�����?j,
��a[�5m0[v_-��q���>��� x:@��M����������ug�c�0
8��C�qd������Ͼس� ����v������_	?	�LΏ�>/��~H���̘�o�;�1w�����}χ�v��O�=' �L� m������@�cl^������|apy�_�f�Ǝ�3��%}�=-��� @�u�zxf����ƃ�{��;&�����ǿ�ǖſ�v�޽�����5׌���  �@hs�S�9}�>&����]=�]���#�<cc���������֜��  �@�t�9a<�2�yl����c���Ï����:�+�����mK�ƾ�p^�Е��v[ �Y&�:Ts'�S�m�}Lg�p���p�Xo�Q�?ƻ�h?��חf�<�wꖅs��h�{ $�w` �b>���}����L�۽�܏&煇���c.��zvߺ^�5��k��K�柞�wX�C+�6  Q��RȲ�xu[�Xx~x L��*����v��M����� ����K�;\�5v�9S_����y��!�xB=���z8��y������p�xo�gr^����0�̖��vl_�3�O�t����Ϲ) @�� 업ŉ�p�D�����}{#��DO�wj~�/ゝhn����ᰞ��b���O:����_; �t �������X:��3|ض;ط�`�obn<z��ag�rϰ�d��Wc�kW8�g<1g,����ݥRim �6"��1�`?4���_��k��Ĝp�T���ީ��{��Y!�(s�FXT�w���{&b�����% @�� Ps�z8nn��ټ���\.�=��ͯ�5U<sk������e[C����(�;ȜB)����aI<�ca,�E @'� tW^��q��#��o�������ɼ�5;�S�׻��ј3o,��ʃ��[Y���DXP����#ė�L����  �4����r�/5,�v��.���z��[��9~}�t׉�݋v�=�q��3�ZSҼ��/��Cb�/,N�E�Saaw=,��CW�� ��� $��w��Gq��=�:k���=݅��Yo��X#;5�����˻�L��E�~`t�e���м>���1��1�'C6�,  O�@��\7r��q�z��S��y��{�y��dx�����'B�1�ӅE�yW�x�8g2�[��=��X��|�k̚�W���]�q>�{�?g� ��� ����_�3��xL+.���;'^Zo��M��gL���Syq�d#�?��z롻g"/vM���tV(��k⚯)���a=�P��t�Bo���#��Kzo����w;��l� t����84������[{����P��g���؉ɩc�y8�>�L�aa#����=�Ѩ�L�����{Yw�>=ݝ����TW�
�������Bs̳�Ѝ<�P���'�Ph4�wnz*ϊ��BV�y}:���#�B}��X�^��=���Ү���1������b�
]y}�&m @k� �.?��cq�}ϑ�6�h4^�3�� �R:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @: �r�<?4 @�� @�ɲlQ�R�_.�w h hI�B��8|# @�� @Kj4��6"����e���pI �6!��V��j���R���  m@� -+��8t ڂ@ ZV�e��š��o hq Z\�^��B�P�K/l����1��  -L�@���>���:U��j�3�� Z�@��`���������<�bÆ_\�jս Z�@��e˖񾾾<�B��_�����b���[�hU Z���H�Z�>������q.��M Z�@�6������{l����F�	t h1��óB���Н����������? @� ������~T�^����ᗍ���
 �": �����s{���E���7�H}��  -@�@�q~{��N��~u\����@+� ����n�����3���q\  q ���5k�T*?̲��O�krq��{K��G $L�@����8;�3�<�P�V�����M %��MdY�� �S\�b���T�Z�)�J� � � ��x4�Q��f��y~]�R)��� $F�@�(�J?�V�ߎ��ӞH��V�e� H�@�6���1B��s���1҃H % ��'���z�Jz�R)���k $@�@������'�|V���juq�T� �e �L��W�}�)�C%F�����5�4 0K: ��y��}jlllC�;����jG�722R 0: ��/�pG�R��������h�ƍg�\�r" �A&����j��x{�N���;SSS������� D �ЪU�n�V������ׯONN~itt������	 p�t hS���(
�ݳ�!.�/��X�~�i����	 pt hSCCCߪT*7��OŲB��j���R�ts �L�@˲�� П��x�Y��sc�" �$���Ũ�5����OUO��7T*�g���K   �\�^oWW�+�t^�)���p�Z=���E4 `�	t hs�W��+�e5N���s�m�v�ƍ��5l �4�  ˲u�����������SSS_]�n�i�W��; �� ��*�J9No
̄�tuu}-�����w � � "��W������	�eY�����-�J_ �4	t �,+�<����f¡q=��R����  �� �T*��Z����̈,���H�t�V�````s ��H�@����g1�o��33"Fz1F�G�.��: �S ����ߛ����8=60��*�Jߎ;~odd� `?t �@]t�õZ�͍F�+�[�3&���������ό�^ ��: t����oT*�R�~(0�~7Fz!F�[E: �J�@+�˛�������ӛ��y��3V�X1 �It �py��;˲���3�M۷o�ݸq�W�\9 �	t �p�ryg�Z}c���P_�i�MMM�#��"�'"������R��!No�GO`��frr�����7z&��#������b��'˲�3.��k�������v�`�t �?�H�x��gǘ\�qq]����?���;�< �� ��;v�cD�����j��q�( �^: �S��_W*��fYvK<}Q�@xo�Z�R*��0 � �͝�k��o�y��x�s�ვJ���� : �8}e�X�Z<]86�_������� :�@ ����=1 _^(��~D`FeYV��'+��o��� t4� <�����U��W�y���3m^\�?����_t�E� �X xR�R�ۣ����X,�u<=40ӎ���y�e��ʚ5k
 t$� 쓡��o�_���B�ps<�̨,�N����Ӎ7�b�ʕ��#��}688��j���8�|��K'''���Y��#���R*�n]�~�oeY��x�fT\ӷW*��/�� t� ��������<�?'��+FGGo�j �ct �))��_j�,Fz�J�������](n�V��/�J? t� <e1��!F��b�!F�����yx\���ddddW ��	t �ii���V��f�Ѹ���������Ϣ� h{ x�n��=�I?:0�ΪT*_-�� �5� ̈����!��,˚�I?)0c�nZ�~�?�S �m	t `Ɣ��;k�ڋ�Fsw�f�ܸ��~���ڗ@ f������J�qzS<~+0#b�����E�� hK �q�ry����������a���Lyg�Z�r�T�D ��t ��������?���20#�<������npp�{��"��&Fz#�V�?�ayy�,��%\�n���_=��ӧ mC� \�T�X�����|U��?���y��c- �6�	 �W*����3Y����nذ��V��= �: pД����j����������S�eٜF�q��͛_�bŊ� @�� �A500�w6l���O�<��}��r�0 ��: p�5o�}q�XlF�sOY��kk���n �4� ̊���{6m�����㟎������������_�g�| Z�@ fͅ^���o|�]wݵ)��+�T=������ -K� �jϻ��]�V�ջҟ��l�*��g��� -I� I��]�ͫ�=��}Q\��8=' В: ��=�J�;N�g΅��uV�V�>��� Z�@ �R.���aÆ�4������Y��<�7m޼��ލ�z: ���k�j�ڋ��J���_���[�n� �W Z�@ �400�7�tjj�x���>+
���˯�袋 �� $k�ʕۆ��O���۔eي��Z\����q( �2: �����z�U�T~�˼�m��e���f.��w Z�@ ZB����5_��;�d����qf �%t �e�H�n�����@��x�xBq���|hh�[��	t ��~�V��,���k��H�X,^�W �'���300���/��W���-Y�x"��V�/.�J� �&���t�E�K�����gW����_ H�@ ZV��;֯_��1�o���	<��>�]�V�W*�� H�@ Z����}�]vٯwuu�e�Ӟ��o
 $K� -o͚5�����P(4#�%����6l8uժU� �$���044�=F��c�>���V���~_� $I� m��7n����ɛ����⚼yݺu��W��; �� ���+Wn��������q��[W�X<?�k �� @�Y�z��鯌1��,�^�ۻ6n����+WN �"����'�_���uK<}~`�,˖NMM5ws�D  ) h[�H��j�������qA� �� @[xp�ƍ�����Z�e�
4�hÆ��jժ $C� mo�ʕ[j��iy��m<=,���ϋ�@H�@ :������_���B�+�����,;}xx��FFF& I� @���Z���F��W1P��vh__�+��� @: �Q��R���c��B�lo  �8�r��1�eY�G��ů�u�֭;���} `�	t �#�H�p�Z=!NB�[,_�� �N� k������'��i�s�%t�$t �c���4FGG�R,o��?:P�e��iӦ�/�pG `V	t ��m�T*���o�X]:O����o���:� t�r���j���8��Й;��V� �N� D�R��J�ri�eá�į�U�Y'� �رc����^�����,=ihh�� �F� ���4n�ƍgNMM}'�.$˲�m�`	t ���\�rK�Z=;��c�f�C
�_���Y#� �T*�R�T>����� �J� <�;v����,NO
 ˲#׭[w��ի� �
� �FFFv�_��1\��)��
���A��� �8��Z�^��`O��I `Vt �'�e�`��xm��6�9t��%� �������j����c��eY���Y#� �ı�{͝w޹*�)��Z��5�P" p�	t �'q��OW*�K��3���y�<`t �}P*�n��jk�����eYvB� 8�: �>��W*�q�>��=W�� `����899Yk��:�,�  �h�ʕ�J�8-�6�
:���  �!˲O�6���-
 �
� ��S����#B{� � `?47��V�_��3B{� �D� �<��>�z[z��� �B�̒���vuu��7���P(�s��pOh_����0KV�^�5�
@�ɲ�m=~ms6o�ܽbŊ� �A%� �S�T�5���y7m�Է}�����������K� ��/�p���y֬Y 8�:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $���╈�B�    IEND�B`�PK
     �9s[���z"  "  /   images/d4c851cf-9fb5-43cd-809f-e1699313b4d2.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  �IDATx��	��yǿ���sg�ҮVZI�@Q"�����lC�rRA)!l��ep�XX!�2C�p�#�X�P��!�х�՞�;G��_��gFI�����U�_�v�{f{z��}�{�^�
uEJu SH�T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu SH�4,�|页Я4�!m��%c ����b�����=Z��vx��0�Y �<��J�N�A?o�џ@(͸�	@�0.L��r�]/�4����F�nb<\��h��ᅛ��pP�\� L5��3}<�7��?-�<�S�:F�[�X(����A�t����|�|M��;s-�i0{�vH�<�x�IeE
�e�6�xwl�4���6�I��<���T������$����֊�g	`��<�	�),O���L���>E0x��� ����,}�Yk؇��X����|�gʅP�Jni0���|��1� ���tZ�����>�"u�̪�p�ҏ�Z���j�%k�-�1 Kxi�u0��yؒ�_Ja���C9�@$�3�:q��mɺn{���;
c.0ֆ`�O��ϫR��Al{/v\��x�%��5Ky��#���Ϸ=���+�%�
5{C��Iyr�nP�|��.�^�a;E�wU�<<�%S��L춓�-oMq6��}�}�4��j�ek�D���Xa䢊���(��%E��Z��پ��)J&����㉓�uc�g��I���{L���G0��:cګ�ձpŲ������j�2�~��F�'�T��8 '4jڬ	�8�p{m�e�AL\���~��m�9cL,6:�(BJ�`p~��d�5m�om5M� �� e�"���y�WY��8��O�Z�&@�X�|Lk��� �n�1v[��3Zc�n���q%k	+ƅ�A!+���8�{]��C?�-7T���N�%5�_��Pp����m���~L ����J*��Ё����MI �N��j���B9�"�8sl,�Ⲽ�r��ML&^�(��5}_�>>A��]�Ӳ�
��3%�L���#u����C������1���u�	7����G5�@��Ko�w�]��ʸ�}
���͆q��{�Xj�)�+T�/o��MWJv�HO/�u��yފ����i���۽�:>�L�
eax�s�i��/cj�����B2��~�����V��qW�R�椪Κ�W��)�qV�@1�̋��=/�/$m�c���P�� ���6]:/c\�q�����R�@�ˮc1�/ߊ-�Z(�3�������'K��?0�?��-��5����|gA�����L��-�$�R��)�`4������ʾ}v�a�����(�@O�F�q"��k[�]��h#�P���\�{�=�p��AiL
��Oi1�S�DAw��˶W}fY��0YUd%�ti�3П�w�C���[N�Z(4 _��5�d
<��r~��!H� F%�%�����~�����,3p[�����L����FB��blk��-i��Fn-�P�]e>�fC���a�����N�����A���Z)4 IY�~䀵K)LP���h����A/�B������C�A":a$S�P#�$˰W�T`����9�
���9�^��>YG�8�.k¾Q#>�@�F?OC��i(�orG�Z�YW�ފ� !���-�N#%w�j�Ѐ8L�B^�iP��0��OE4�>�1ޣ.[�J1�B��L2�H��V���.	{[l�
�"k��C�,vtU�K�����K��I ���ˣ�e���s��z)d1��:���;��a ]�6�|��s��-�,0U��:�b�g�q�("1�m�u �cY13�5�\/���M��4-��3E�8W���@ �X �/�mL�J�#�Vu�W�ˌ�.�I��׀�"�WD���m�S4�H�0�X��'W��s=#+�eEH v�
a(F܌e��(`���V>a���n�� G*��uÎ5"�}�K���jF��`X� Cӝx�����瘆��l�|w�� @R�gm��N1Rur=�`�i��yp;~��-����y��2�`��9�ˢ�3䙔�	�]�2��T��3�0���N�W�I�g6b��w��1����H)�
�1_����u`p�.���%B�e�{cv��ݕ���[ST��3�?��a���.��R�PW\P41Ȅ*&�jaZeUƫ��t�%�h�$}�#�;O�]�<�H����|�`ڇ[��,xV�{+������͢JST]��%U31P$?Ps�>G8�kZ�AGѳ2hE	�
���P���t�@A"��ܿz��֍���[���ᘦ�x&~� � �+Y�P���޽/���1���)�B�� ڄ�X|�X����������E7AX
�'bŘA֑�j�g,�q�c��OЪ^G�r����7���iA�;#>T �� �:T������"(�!��h��7Yl��N�2�E�GK�Y���s��;mP�I���2/׶v�	��-|�,���s�/���:��H��w��qM���#%�'��T&��_�)s<P^_�ng@|��!������A���E���do�lN/@η�߆tj����;�<t���1���J�g+-�ڑ8Z�]��Zh@<ǆ��3@���5�;��s�n���;ت�#�dR�
�7K�M�A?�ǳ+�C��!,������8��G[���X���*�̟:���8%�7��K4e{便C呮Ύh̄j�sY��btϱ0ߧ�����x�����}�o�5��[�q����G����� 0]�'k�#�Gd�m�h!�4�&�h^���z���s���c�����	F�
�+l,��	�uK�L=��G�@vmZ	�b�\_2��E�M���qt�ze�/�%�()h�;C;�pǲ�4i�*�g�`dL���|��*���T9����0�T���a)\ e��o=�MO۪JK=k7��9ƌ|og�&�Ub�B9ȕ�_�GB�Nt]00��$t�>��a+ĄR`,Q����P��\OG�^��1������Ԙ�k�����B��*��eaDZ����ʍ����Z�k�QmM7���P��\[��v5�7�a�u�A�r�H<Y����K�,��cƀR�)���C�9��1����bq�)ji�ա����++�=r4U3�Msٔ/ u}��5+�d���B�!���'2��u��76�٧��I-i��"����D0�!)�<�uC���μ@��̌�ؾ�#$1��8�b�v�JxN�pGV�^�Ea�����r��	ZȗlB�!t���~��-5��;oj3���S��v�l��s��b���% =g��ؚu��(�಼'���Y倻�Qn�\���3��Z[��Ԥ�tPyxo�-Y�`J)��}�
�^�vĠ�O��|	�Th@t& S��d�"��%ʭ��i-줱X�1��۠�1gLh�F&���I(8>B�S�E_�5}/�Ha)=$�%�����
��P4�h�+0*��Ƙ�H�z�6���[��RZ���O���~��W��D����BB�KsV{��a�܎���O�ЈY��3Ʊ^��w7wó����p¨L�����֖V5�@��}��K�D�₦0N�Tyil�r�lX���:�=k��5�M��k�ܻҖ�6Wr8Q���orCE��5"���a��\:kƷ�ٷ�v��`K�Qg�Ǡ1"e�YG��9Ț����{[z �)�!��2	�%�pT����X�Eۃ��B��`��B�Ɋ�������W�q=�f�_��� �	Z~q�W�
Ȓo� �/|�̦�_�	7^z撞lnU&��wl����+��9=W�R%�<�ߕw�#���vO�����i�Al@+Qh�-a�/XC�We��;O����?nn��s��=�C�j���;�<޾�7p畧���~���<v���\ws�п�s}":����R���Q��W�c���|mӬ��Y�D����kPK�d�܏��"��}&�p�z����K>����IZϯ��x.�r�gAK�Q�I�@�c��1�d}c���;E����5�.�^5�J������y�
��>����ݻ:L��21�b�`�������A�0���XV�g�0�v�z��Ǚ�U��R��izz�s�����S�'[�w�p���؃�j0�z�fB�V���!'4�`e�_َ��4�~]�t�':YRZqGLp��A���Ն&ն����ͦv8qp1�\�� ��q0&���߹>���`�9��T�3o�&2���_í��.��O�ͅ�'�����j�k�KF�l�l���l��\/���__e~� ?�3A۰���kZϡ*�@�E����Y�.�pc0f�3��u+�Zf:��d7GK
<M�򫢎�
����a8(�@������w=��~�Ec��Qа��Au ���\Y�ݧLn��u/@$|��V��9��ic8@9^�Э�iި^��,�IQ�2�kM�� ^��]����ǡ�ˠ�A;��i0o�<���=���}�a��ˁ&���|�
���E{ �E+?XYЎ�,/����b��h#��k��?~i,�����H�����b��/�ȨA�@HT�UP�CiA��-²��5��� �
�r�JV@�|��1P�_�e&�\���B�
��K���q��~��Ҭ{��*��+ �}��j,�byJ�Q��w^� {.\w�q�Z��>P�c�"�Wa�E)�\,OD�J�d�a�C^۾�5X��Ox+Y�E-U���]��~�&w8���n�1�����gbq��W���6��"���)ݿ��i��	;�V(x|Z}��U9>?�cEH��>֕��\"�H 9�}��5<r EH]{T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu SH�T1ՁDLu ��=P��&q    IEND�B`�PK
     �9s[wJ���  ��  /   images/f9728bc6-2422-4ead-9082-90351081a874.png�PNG

   IHDR  �  �   )��   	pHYs     ��  �8IDATx���	��e}�����sN�{���  �NpILbL&���'&HLn�F�u��%��Y43sI�b���q>���I"��+��4�4��Yj뽧P�j �s����?�.h�p��_=���   8�:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @: <�6��䪹��|X�&�L.,�t~'M���L���t2�ٙ4�	�l6M�����l(uBZ�>���f��?�[NL�~2���o'� �d��L�L;�]I�<�o��;����W5 �: <��û�;>-d�K;�lX�f:K�>f'�t8��p;mW&2�b�s(>�F���7|⍍�dj���̤���X����ه�$ݒ��9�z�}���[ ��@``�n�f8��8��ɞ��U�L�|�W�E�К?j#�2O�7x��I�B.������?|V(=�p2�9����O\2��d���Ω�8�J��d�w>o�����F  9��@����[.��j�ON�:�d�x��Ei��B��4�	��!�6�������k�ۍ������U�|'w&��]��Z|u�We�� `�t ���^qB�&���3[��QI6YR�4���1�b��<�ւv.,h�p��z�D�ُg�o�إ�Z��s��ұ��^��� `�t zڍ7�X�w��gwBxq���ʵ�ݛ;$���I'�)7C�P
ݏ�������o�̵��϶r_�w�m�λm���I  
�@O��o(ݿ{�w�'���;�w�|b:ӫ�I�ۅ�Px|��5�ڹ��'��\��F�������� Ϟ@ z�7zd:+���֋�Ӹ��d�S
r�l����Cn�^5��?ټ��$��N���w���� �� Dg�������$���������ڒ4�D03������6NitW���u��Kv����3�]5��nZ< <=�@6|r�±�ɋ���/?�}��N�Ƕ����~|�\�!�^����_\�y�w
��?e�e�n����  ���!s����/,��]H~��c�v*Β��N�S�����\��͗|���ڕ��ض�n��� A�0�F7]3��=����B��zh����N>�7�W��>f��K6��F����P�|���� (���ۼys��/�v��^=��rb'c���N�^��
�l�����+���r�k6�S �#��6����c�C�?���g^���&�i=��X??��o�؟�e�U�����߾��Wo 0 : Uw����W^��4.j���f6�3�ʶ�J�ՙ��W���5�*��[FVW>zU�N �>%�8(ֿ���uJ�?�T�3��ζg8���5
�S���'�oY����'7��o_���  }F��ߴ�7ZC�׍g��2�]�L�v�=��]U_�}�%���Ul�޵񢍟	 �': �Xw��/^�(7���luE��]U���¦7}������{g����m��	t ؆��0���n��U�B{~�C��k�l�64>��㵷���\k�/�ܽ� �$���4�w�G&�ӵ�w��;i;@dZ��⩏���^�=�Z�_���� �C: O�M����K6^�]��V rIhM�گ��/[��u�+����Ƌ7> �t ��+n�bE����z���f������d:�j���L!�+k>��S�f�τ: ���y�Mo=�Z�_1V�xY7p��4����K����~h��.7����{��  � �7�����{J�^��N)@��d;��R��R㗧B�$�����k�=  "`��n�f�]�q���دw�9��J�T]�[���������y׬^�:	 �0��}`��kC[״Bkn��d���r�����k�?��~o�� b`��}��_h����Dn� ��m-m�n]{�G.}�Hk�������z �CD��� �ɡ�_W���i�	������5��O�ټ����ٗ]��v �a�����7�����?�3�o���� <�4tr�B�ōv붵������v>��$����M���=����j��I2��r�u�%�������k��� ���n]�*&�O�'�Oӎ���,�r�Ò��Mk>������o����  �H����t��Jc��
h;;<7��f���Ks�>���ѿ��5? `�t�>q�M��i_?��<9 U�K�Vgծ��Cks�МK�`:t��!ݐ�����R�u�L��i�=.R+�/h�[�^w�e�_w�;�> �A$�zؕ�\y�O���z�~x fD;�OO��K?��?d�7\���� pt����+�x_q|m'�)xf��䖍,���M���$I��^p j�ک��ֿ��e�o��h�� �#��c6|r�½��7���� h&��I�O,OUyw�:٘���KvW��w�v'����b��O&	��H�/�l^����|�-��b�; Ϛ@�!k�7�k;�=�*��8H�Z:٬v��C�����FrݏsV�?��4;;'w�wN�l?2�h�ښ�~�{6�Z��x�Q�n[��+׹7�gK���7�wƯ���/O�Խ�t����U�U�'��B��]>kY��q����ڵ��M>�~trg��nX^��ʶ%Cc7]�������Y��\� ���� �]�=��Yh��˘鲧���j�����|%7��v?��ҽ��ɶ��[�Ƕ�j��@Gi'���P�5�G����׵�����o	 p�:@�W[?���`��n?˿43�2/��8y�I����㱾ml[s�16��^�7��-�r��+.�x�;�g � �"t�7�=瞿�(���-�̄��x��4:�\)�\�>ݳ��/:��Q��%�Ƿ7ܷu W֓L{dbx�������^���^ �g� ����+V|����7�ͣmig&��m/��􀶹���ٹ��ʉ�N(��j?��ֶ��[�=0_ٝ�f'K�՗|d�1Ci���^}��  OA�Dd���_2>T���m�0�v�v'S�~������-,t?N^zr���#���jv����m�|�$���o��[��o~�o� �It�H��������7v�L8vM>�s�,��g�׷u?&ɖ}[�y���Iߗz+�Z����[���u]��  ?ŋ@�Clt�5�����&�p��M�N�油�{0Rɝ�䔡���nݿ���]�5����N�S������?c��YW���'��������G�����KӴ���V���ys�|��yG���wD�{V�{��4����������b�U����Kn��w߽��c �@8d.��������i��ݓ{���'��Y����任�o{�oC�Ql�\8,�?/���W���Wo <�p�}��M���I%@DvW�����S��;{���'4&��v��xp��fw��ߴr�����y�6�f� M�̰�}C�R��08b4�Ix|1;��9���{N���=o��J��y_�}6;i�I;�̝�ݼ~��7_{�� X^̠K?��/'˓�H�~Z������ɜ�^#T�ܩ�N:nѱ�{����T�������Y���nY�꺋�{W ` E��/@�ڰyCqof콵|�� ��]�]�?��/?m�ǔ����C���B�HC'79�X��C돾���] 8Q���O��|�=�������s�G�;�"6\ɝu�Y�G�;���G�]�S����Ӵ��,U_�f�9sk���`�t�i��}k�Ndkk�G��"w ��_|����w<����j����#�G6l���V_� �0MF7�.�7?�ʶV�!�V-�6��Pq(z@�z�峖��ZZ����7���z����R�P?3�3��oX��W�4 }O�L����^jn���%zЮ�dUqUO�2!�9f�1���,/|�o�v����J��k��W��'G7]�/�|2 ��:�A����=�6���8_�G��i����zP%?�;oŹ#�M>ֺ��ժ�ɞ����5�O+�ӛ���W���޾; з:�A4z�[N���}0�&s�����=���xxq��������߷���^�?��o1>>1�i�U/��X �/	t��d��ѳ'��ޗd�� =n�1�i&�N1Wʆ���2'.>��b���W������g+��k�J+῿�����m�}�� @�� ��^q�D���~���7Y:kiO�f�f�^|�G�C���w꽺���7����e�/{�;W�� @_� ���������ć�L{v�>����=��'�"��������}=Y�\kI5>���7���?�jO �ot�����\U�5y�T��	��/e�F�{������.�ν���ܳ�������H���r�^߸k�ޏ�n��妻���,u�9�W7�2�a �2ݳ�'���T鎭_�|t�Ѿ�7�{j{�����sܡ�d2��	�N�,^R���/Wk�Z�Mzo�Gg+���k.��[.�E����,l�䆅;�{���m-`٬�Ӗ�\)�+��G>{��C����� �@��,��m/Z�7����������#_�~Wm���V�1�|��y������~��W5 =M�<CWn�r���ޏ����U
����N�,Y��V���8w�S��6��{o0l�䞤����-f�_y�Ж�4���7j�6@�^h>o{��7o��իW��'�O� ��E�\4<��}��o���9+
�N�y7Ɵ�ǇK#�s���s[??ًgx90�M�l���������3G�;�4�27�Ň�\��&{jwH-_;�s�;�a��k =K���잏�=_?:��r��9}٩CKG~���EË
'/~~��~��K��;����=~��U�UsV��ù�������-�w�v�?�S[ޫ�ڋ�~h�;���k� �$�p��x�o��Y������S��2���x���G����=��k��P�g罍�ǂ���Q�(6{y�;h-���W�3���{w�SOC����뿵��o��w��! �s:�X���WL�����T�dNYzJy*�K��?m�����d����k�k�ڻ��j��r��y����O�[�OXt|yNyv��۾Zk��1k!M;����KG7�n�x��� �)�g�tӺWV+�ׇ>�`hA��gU�C�z�r&d2�<k�S[>3�kgwyv�z�]Q���5V�YQ<n����\��g��ZV9�E�;�~a�W��Ӑ�&�k�\z����z�Ư z�@xk޿�����������p���OXt|)�`�\){��s�?}��'�4��F������=�|p��fw��q�+�)����K�r?ԋF���ze�H'�)��4�a�=����� ���`��ˎ��j��	�g��;f�|)s�ag-^|P�ϚS��;g��C_x苓�tn����{�������[˧B��E'�G�hE��+f/<���Z�W�-�Bknfn���M׼l�ŗO �'��D����l��V�5;������sV�=T�W�%���ZZxޢ畿��;&��n�o�
���B}圕���P������=�q���*�B%{O�|}7s�U��[7o��ݑ?��S~p����r���=����KO*wCc:�����x�m���������[�omn��<j�Q�_�=��b����H�s�]�4��H��8��7N=\ ��@�){?8vu}����G��(������9+gd�~7b�\~�P�Y��S�c�n�uϨo�}�m�j=�I�UsV҃0��P[5wU��+f���+�I'�c���W��z�W7���� �� ?f�ͣ����W����R��9w������s~6�͜����O����z��G�Fy6��z�+ۿZ}`��ӗ�V�����/<��o�c��n��5�	��H���n����w �$�~�[�8a�<yU��=�����y�sW�3\Η�=�����[q���~n�V�~�������S��/<�|��cK�L����[����/�}��&b#��픪���]���_�z��� �� SF7]3<Q���TB�8l�a����!�y�y�3��6���_�?���"�}���Y+Ϊ���l�� /<��<p�dw�@�X+�Z\��M=�� @tz�D���Uy��i(�1�-���r���9+�������ƚ�ɧ�m���Ǖ����{x�t.�^|�F��E&�QGz5W=cݭ����W_���t`����N�'�} 3�7�.=�r�#������O*�7&:;�w��Ώt��߳����ɝ��54T�ٳ�B%��#~n�3�v�ښ�;���׮ߴ���^|�? �!Ё�����~y�R�����\8{�YC�g-+�u'w�}ؙC�=p��X}�������=ɿm���ӗ�Q9l��(��D���y���|~b�9m�wB���4�j�=�wm�Í � Ё���}k�6g�ߞ�NϮ�=!��g�[u�Т�E���=��:o�S[n��~�53��i�_������j�����^ ����#.��qowO2���{6�^zU�h?O�A"Ё�5����i�=��/e.Xy�pw[���sV�=��?7���?����4�+��8w��m<��D��߶��Q���ǎ}h�O�:���x1p���e�Mj�׽>텇_8<�cwJ/ZX螕�{�ݵ Ob_m_w����+�^0��'_�tߌz�����y���w�L�뿷�W�۵�{�g �TO���\����t\��=������_0ܫC����ƛcIw�4���F�g�����N����*����{�������N��v����4W/W��t͋7^|�d ����@ټys������N�Y=l�0�}�?7\��������\�Ot�|��It�L���w��7�;�,9��Fru�31�<7���n�I'�/�V���Pz���� 8d:0P>���_7+ͣC�A�_8��>z\���sV�5tۣۖ�x͡����5�I�s��Ӈz���6�sV�5������ja�G?|����� ��@������j��[��=�G\82�=98������+�����&�S�<��������y+���z�ґ��ӗ�V���✽�	��B���z�[?��׾m{ `�	t` \t�EÍ��5�|�Z)_�\�����j�t��t�Yy����1i�;O�{�{.����z��s/M4':��u_#D�{��Xe���z���'Ё�0墫k�ڂУJ�R慇_8�k�ڟ��Ë�_|R��~��i��I>������p��+�\�w��'�������F�qr����.��� 3J�}o���p�4��У
�B��V���H���]pLic,�ne�4ƚ��g��ąG��H�Ezw�ݙ���lU'���&!B�����6_�?޹��� f�@�Zwj�m���ޫ[۳�\8oչCsʳ{�����rƲӆ&�������1��t#�S�^�H�es�V�7|ۖ�LT[��Hlg��Fho�z���#Ё�����*�V����v����-,���d3�!`��嶉Z�]���#��;&_p�=w&��������?3��b���.��k/��#�!Ё�5z�[N���[z�)�N�,���P��p9*\>=��It�B\���%���~�H�Mw�]��;�3*_���j�L�v2���[F7]��/�|2 0�:з����������_:jޑ�0�����<��ʗ�}���������C_��n���=��ˋ�,8&����E7ٽ�i�/�v�c�� �N�}i�-�]6��86���+��脲$�A��/:>���{��ӽ��·爵uؙC�y��<�I�}��ɮ��v�L�X{���������� L+���+n�b�����4�2/w��3z..��	��W�����m&��3m��P�R��O\|b%��L�d�^q�Ч���x�U����NH����_m޼��W�6�`	t���˭�w��r�1�|��Q��΁�Yq��Ӈ�ݳ�~�{w}�1Rɮ������t��9�����D�F�衕k-�����S�	 L���5�_s~=_� ��\�{��������E�͋��b�]��\��];�V�������=�Z�{kA��J���b��Vn�����o�x�c�i�3�h�d8�ew;f�1�/?�2(w�?[�B���?�����1]"�I���m_���#_<����N4&:������X�={���/i�Q�����P�X�˩�� L���X����1�������9+�:�gj^e^��e�}e�W�����4����/:�#�C4�=iZmLv�N�������2�w�W���������q�\sg ��@_X�y]��o��5@*���́�}3c�T��x%��Wۗ|�o�NYr��t�\�N;o�'�~�c?|�]��i��:��1��? :��N��v�=/��r��9w��C��́g��%�/OL��#��������[�����+�8h;U����7�'�kcI����}I�5�	���=���_}�k��5 pP	t�獾g���r�7B���p�ag�r�������Y+����OOL��@D��]�]�_��*=�Yi�]�O}��v���K����}Xa��ݰy�ǮZ}U3 p�t��5g%oOB���S:~�����Z!�Ϟ���������a�[��N�闷���#_0�T�V���tj�ǚWL=�� �A#Ё�v�M�g6��sC�
��	���7b5R�-Y��՝���'�g�wS�����t�W꯾r��z��� �@z�p��{�Z�b��9{ř�aUΝ?Gͤѹg׽�G'��{w�SߺoksP΋O�vH���[��9 pPt�g��u���)������J9_�7b�I;�=[�켧��m=�I�4��^n�����5o���� <g�Y�|��ǧ���UsV��^��gi�?t���m�o<��z�]X�$ө����*�e��L�=i��ֿd�P?�Wf�U
��)�Nq�������}��w�ƚ�Cd�����n}�Ƌ7> xN:Г�#ɕi�����"�Y��Y�N<#�N���G�U��M��!N��)%��?O=\ xN:�s��t�/W�c{�׎Zpdq��BW�=C�M>ֺ��j�V�vv�\�T���7�u���yێ ��&Ё��n���yw ܉�N�X#it���7j��ok�'$�S
�ڟM=|c �Y�@OY�����G�q���*�l�'�L��T�7��qw�tv�=�R�������x�;� ����V��3�3��,,Yjk��^���ǾS�����I��Z��;�}m �Y�@��y���������K�ok���%_���ɱƘ���㪅�/_r�%�߽��c�gL�=#�t��ʽ�'-9�\̕Lm��[ڻ���4���@'����d��� Ϙ@z��{F��U�	=`nen��yGO)�$�;���Yn�j���W�^�:	 <#�	�Y��NH���.�����yR�)�_����=�=^�Cje��P��k�� xF���=��,6)���*.Z��)��o~��z��9��F��� ��1/"�����C5��k�L.s���O��GZ_�����������lZ�+���� 8`�چtCv�'��F��/<�T�W�{��}��_��A�à�T�?��N�<���&/n��ȕ���1�.~B&���~�����o`�4�׿o����k�	 �D�Ul�v�'->������I�]�]���P'�ٴ�y��õ�"Ёh]v�eG�&���]��[5wU!��������0����Kn�����_�zW* �D�]��Iw&D�E't�Y=��4��W���@hg�Y��|o��� ~&�Di��͹�
��B�����ܲYK�F��@7ο��+��c��9�V��=�$��@�tG���*���u�UK��?!��C_���!΁i�'u�,����~ �i	t J�r�������Ë�=?��~��w��9�ӺG�Z��uS� <-�Dg��F���UO
�{���\��C�������O�Yh�tC��-We�� ��@�Ӟ�yC����V��/v�|ʃ�lܳ��F x
�\2w��c�q��� OI��i[�"w��畜=����]��g)��:���@Tֿo�KƳ��!b�K���f--������������A�7�F�q�%7\2��k�= xR�JRIW��������^o�;_����N���	i!������} �I	t *�|���R��Y9g�@On��F�n�xFڥ��)	t ����_ޟ�77D��yG�2��@��}�7j�����j�'�yߚ�7��� ��@��ʶ~+D,�͇#�^l��m�-{��NxV���gr�ߝz�_ ��@��!ݐ}�㻣�޾r��b1W�����4VK�|�.ہ�$��J� OJ�Q�����s۳CĎ�����'�v��m_�L�Ĺs�9i�'n�䆅W���]�� Ё(�C�+C��V�����s�7�Vm�9�	 �Q����D�N�w ~����������'v�"vԼ�v�|Wug���8w4�b���.�~�@���>����H�3�̊��2�۝v���w��`g;p�r��F7]3����' ?"ЁC.
/[5wU!����j_{���Z�fk;pPu����/�zxk �G:pȵs�����r W���u��V ��B��A���R��FO�+B�F����+�r��������wW�4iۧ ~�@���e'���-�j���T�����켧�h��}	`�2�W�r��W_t�7 ���!��/[9gE!���D�e��� 0͚��+��� ?$ЁC�׫�>)DjAea~�8���G�^�I �n�Br~ �G:p��zϾ&��^��b�a�z�����c����h��]t�E÷\~��� �@�¬ܯ6C�2Sߖ�Z:P��I;�7�f= ̐NH�.�^��� �@�V�}f������r����p���7��Iw�3���� �'ЁCb���G�
�:l����{����|�`8`�%�4�Y$ 3M���xc��B��峗�������h��Uf\#�\�:��P I.����9�J�20�����!��Nnɲ�/�z�?����!�)$��H-Y:Pύ߳zbI��� �:ph�r��C���,�v���f��A'�� �����-'�e�Fy�y![�t'�����9�f�q�tC���Un� �@f^���!RKf-�gB&@��{{�X=�$ө�_����w�&Ё�Φg�H-^<0ϋ��h�[5��@���{�@�����.���Z4�p`��칿 "�ʶ� n`^�q��u�ζ�����Pqh ΟO6&���]� �$� �@f��ϝ�l��ґ%�e���4��ģ�K���7�����1��50/F�H�g�H-Z0ωݫ���`+ D$�ܖ�[��F� �@����C�-�����n��"= D&��wϡt``	t`F%���!B�|)3\�B�n����s Ji�sb `�Q�\�<Dh~e~~*�����f����ɠ8`�	t`�\z㕫ja�P�Ђ����޾}lG+Ma� Ћ��N�o���̘����Z�Ӽ�y���o���V����4�x�� H�3��&��e���)���@���]�v2i&=o��'� ����d�cB�*��l!���n����v�t��f�@�@fL'�Y"4�<��Wϻ{��v z�LzD P�1��Z"4o ��w�N�����v ~��$ (�̈u��U&Bm8DhNyv�����v���@��l{a P��f��P���٥�}�|��nu�$�� J�3��vN�fra�8������N��$tJ�Z�@fD'�)u��G���$�v���/	 =�����������ȥ+B�f��{{w8\'��@��:�N}w[ 0�I6]"4R��@�5���v��t�� 0�:0#�\�(DhV��}om��s����a` 	t`F��N�Sy+�J���Ƙ@zJ'$K� ���ۼys�_��
i��P��'��۵N�݈��<�SK��� 0�:0�>߸{qZH������V.��:���VρޓC` 	t`��ZQ�+ʙ�Է�����t��tBR	 H��/Ӊ2Ї���|��s�%�SZ�y]����� ����2QNp/��}���VЁޔ�z�z�-`�t`�����r����ۧ���N �A�y��$w��L�N��*�}��v=�Ёޔ43�Z�@�_.�"T��z�{�ݰz��l.�  �L�N'�@/�J}��^k����4Ӊr~	�t���K�aV�P1��g�k�t�g����(��$Ё闦��B��߁ު	t�we��Ё�#Ёi�	i!D(���{�����L1 �L�L�*�|�ࠩ�������O� OB��.M3Q>���
z�Ӷ���N6�����E3�g�i��5�l����@�f�8Q�h�M�[�s�l��%椓��?��2^���0����=3�-�~�ǒT����A�@�]'Ms��p&��.I��g �̀N�+衯Wϻ��c�Yi&�u*0p<�Ӯ��l���|*��zWR�S����vS-��m)7���=������ui?Q<	�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �  O��h��2��s�dB'_�7 }O� <�N'�U�M.:��C����Z8�� @��  O�X)T�vy_c�>7 �4�  O�2����$�V�5+ �4�  ?�М���B�J� ��@ �2�����9�k|I'� L� p 2�Lgd�T��_��i. �A&� P6�m�~lb���p��_��t�>��!Ӫ�*�\��ods�d�~�����]���5 ��@�S�f�8�ora��� },_*Lv�C�ɟ��k L�Ї�Fyb�Ĝ`.}._��F��:?��� 8�:@I�N�^�5�-��{�B�><d��\���$��D�jjSq` L�y�{�Y���C�y�~��I���� �F�Vi�g��\�5<o*γ�N���� 8X:@K��|��������L&��̟��LMl?P�_�`� =�QkTZ��-��n�/y4��F�O认O}��� <[�{w%�]������^�{k�eyw�Ƅ�!�d�K�$d杼�eN�!!���cb�:���[��p��c��wf�aBl�}1�ٖ�Œ,����.�����[����ߪ�]tI��������F�@]�ͨy� �BIdF���닅t���\uq X ��jg��Ec���xq�K{m���s�I�5�@  ��@�0���Z#F�s6�0^8�e��X�l�hF��� �t �ǧa��F�l�!2q^��N�~�  V � ���4��H�D&����j�թ�� �B���8>�.[��g
��X�6_�Z3[  +�@ �p|�]��l)[K5ʍq�� �F��%8>I�R���܂X�Qi��� �t � ǧ�EIƫ�
sb�f�Yj�Z� @�� �G����fa�8+�j7څ�bsB  �" ������l���y�8Y�QJ�X��������  �e: �ǧ?�zn�8Q�6��V��/Ԉs @O� �C���r�_0q�H,��Lm��J��
 � z��ӀQJ���Ҍ�P,��tu�8 �� ]��i�s(�
��c��b�0��\m�h��, ��t �"�O�#���D�r}�PDn�Du�֚�  =G�@�4�<�?FƋǽ���H;չ���g��  }� t��� K�8/Oe��X��f�<Լ� �  t]n$7�ʦb!s�au�:!�8 ��@  ]�-f�3�LU,d�f���+ �w:  �L1��-e+b��|u*h9 �:  �T.��+e�b��B}2hy �:  Xq�l�Z+̉���x��.
  !� ���2^�0^8!�j,6G[�ֈ  `  �7�6��Y�T��,���1 �B:  Xq������D��ڍv��؜  ,E� �eS��Ek��o���B}J  ��  �E9*(M��?Gb!�dk�i �r:  �`J��8Y<�*� S���8W ��t  pa�D��빁X(��Tu��J�8 @�  �B��xq�K{m�P�^�Du5q H  �/]/�2^K,�ڭ�q��v �!� �yɏfS�TC,�#�,����?s� H^�  �9ˍ�N�s��X�糋�u�S @�  ��d���L!Si-�:W���(-  $�  �*�r�����L���8�0+  $�  ^P:�^̍��R���d�r @��  ���L���ω�j���� �@� ����^�0^8!�jTc~�/	  �@  ���Va�x\)�b��bs�Uk�
  �@  ?�q�vq�8ck�7��R��  �  ��\�'K3�Q�X�Uk���	 ` �  �C)��s�U�X�o��F�1)  (  �u.Qa�x���@,䷂lm�6-�g
 ��"� vq�'�Ǽ�닅�v���W�s ��#� n�8^���^[,�W���-�  0�t  ��.��{�%
�ȭ�V�h�] `�  ��H�D*�j���P�չ���9 `��  �l);�)djb!i�6W]�C�  �� �����bvQ,���j�a� �!C� 0D2�L%Wʖ�B&�ks���3 �"� �l���͋�j�թ�� �!E� 0��W/�N��j�ɠ� �!F� 0�ܔ�,�g�R�rc�o�E `��  �8�[��ҌR��B�Jc�Uo�   � T�봋Ek�Ym�Z�֨  � ��tF����0/4�  �E� 0`�Raq�x�qU(j7�|�Ҙ  �ct  ���ǹ빁X�o��B�8 �4t  �N�'� �Q�J)qG�R��}�׵�A+��檫ļ�   ��@ `0hIɂ��_�M�+�v׉\��&�ͷ�c�w'�v����  � ��R�,�j���E��9<Ɂ8�{�8��}^����x�Ы��V�~��  ?B� �t�T�8o��C������n'��h�繑	y7�|�ǋB�VOTWk�]  /�@  ����S�^}�8ޝ�ֹ�;K�nb=����#�,����?s� �9� �����y],�l����H����Z�xge<  8':  I�J=���Hk��q ��!� HG�*�,����G�8O  8/:  I�HK���XJ��Q�$#  ��  $��v�b�8�G�8�
  � :  I��Wieo��Q)��  �F� `;%��q�u�r� ��  ,� ��B��\QN)
  X6  Kiё�qM�Gb�Pg�8  �"t  ,�cf�\��b�Pg�v4��  �2t  ,�l�;*�0J�&� Xa:  vѝ��勍"���|LQ�  �8  �������b�H{Q;"� �  [xb�)6���q>�D9  ��@ ��S�⩆XH�8Q�8 ��t  �͕Z�u�Q�����b~�  ��t  �ɑ�J9U���J�zL4�  �/�  �#M�v*b)�[{�)  =A� �J�q���R��8O  � �Ӣ}'�,���8�H2  z�@ ���q�ϋRZl��8γ  z�@ �wB'��k3�n!�GE	%'  �/t  z@��ܬ;�y$6
t!��  ��!� �2�N��8�A��@�  ��@ ��t�Lk%��(��8�G  �� @��8Wi� �
�F��D�hT)%  ��t  ��1眻�-�a�_�s  ,B� �*�L���F�N�S�9  V!� Xi�,�q�Eڋ�q ��t  V��TU<Uiq�8W�  �!� X)���8�������s  lF� ����R�b#�U���b�B   �"��K�`h8Ҋ�"6��\�8׼� `;^���0T:�؄k(i��� �2���q�$VFN��빑  � +Ik	�� X�;��*�,����yZ�h:~^�.���L:�峁  � +Č�~�D�9J�8��E)+W3�q>*�d��j{a��|�g4 � + ���g�|��Nƙ׶n5��8γ����2��l&��2����!�`9��v�w#�z�a�EGN�5qn��������V��u�B�wŞ� 0 t �@Li>:fF�E�	l�8��Ϭ 
A8��j�Ly�R��o �� �)����8w��ӊu��8/
�JiU�֙� �@��`vS���>�tg�vG�b�Pg%���2S�͌�|1ϔw H0 �Sڇ�J����-6
uF�zT0��0�Ly���� 	E��9�@�A�
��'�8�[b�H��v4���$3�����g�t&m�^	 �3#��,̨y�z���ʢ��(�^Ԋ�u��hԛ)s$[�K�!��L8Bm�)OU�Su��7j�xa�V�s�� 9t 8֛7e��S5�P��錜�bV���u��B�u" ,G��s�8o�>�͇�#�8��B�8oFb&��s[�Dz����r: �"���'·�#-�v�b#�U��cB��h��y�I�<�ڬ�x�m���Ͻ�o : <������v�b�8ε�s-)��lgFԳ�����E:rˡ��{nx�3rϧ � � 2q��
���1U���b��-�_;�"Z9��С�ƿ�Q|k
�IV��lyZkI��:%����[���}�>�G�n�S��:mqTg}�2�ۥ+79��{�7;�{r�%.��û���+�|�\�����'��ͷ߲��v~� � #�/�1j �W��/ҪPʷ�r�l;�T��ݷ��靯�i��? \(�P�Q��s �.�Z���#�#����>�G��^* 0�t Cǌ���q '�JOJ��fg/��w�������� �`�t�ZOy�&zC8 XI��t��w�W~�����O���g �`h,Ź��\���S-E�Y�������Փ�}�z�������� � !���q^K�!���LL���֏���}�q�k���I6�0Ht Ϝ�{r�8��Y�t�ww���G���o�w� :��W�6��S  ����ި5R���~<3��n���y�=$ 0 t �\`�M �s�(�s���SȵҲO?uۍ��ow�s�n��#�,�L �i�ڞ�0.��X�a:t���#�;* �p:���l�<� ���ly��t:��R�\�������>��s� @�� N��v��  VD��L9�������e���o�o|z��F  ���0P� t̅�  V�9�0Rl����BZ�z�?t��_��?s���"���Y�:q ]W�j���k��Y�n�V��y�K�3���"�3�c"]  ]��2GW�|F�L��տw���O���_ $�` ��9� ��]i6�ugw��k����]����ol	 $� �ر z������v��Ǿ���� 	B�H��vl��3r��ٺi܌7{�o{�/|�}��� @BpQ ��z�F���p �'fyQq�`�zt�z�q��6. �:��2�l
 �c��0�ŹB��r���z��?�W�_ H @"��-�lT$ ��2{�x)/J�SV�GZ���p��o���?- `9@�Ahvfj; X��hzf=��8N,�Cw�q����� �#�$��Z�:q 1ˍ�պ���Od�.���7������E �� �Yo�� ,d֣�z>�vD�陿��N	 X�@�fj;���̱�f-��G�-f�o��[?�{>$ `)@b0� �g��kJ��������Z:�D0�&�� �3S�ۭ��Τ��ս�mg^��������s�% `!����v3mR  �Ь7=/��rW���c�v��o�����i�Zy �����  #�re��Jy릺�Y?����U|��	 X��^ V3�$�tI $JN����"�̌���ۿ|�o1��6: k�5�Lm��j���h�%�ig|o�?�O��_ �� �ǹ��p �\�9���ʱ+ `���02u<G@�ٺa�E��?|�g��>� Kp��J�g�� 0ƙQ�|ֺ��ǂ��W��@`�u̦Bfs! 3#�Lsw]ǪQ�F��{�mox�g��� X�@`�f��� `дM/_��b������O: +p�*f��c� `��~��A��kձk����������/
 ���*����2;�缜U����)<��] �ϸ`F�`��۾��f�֢�y�o����w�Q �#�5=���n��\!g�Z�������_�w] ���`F�`8�Q�L.�v.��,�� @�� ��j�y>�!avt�m��k�x������ ��b }����s 6��k%2���� ��@�wfW_ ����t&�E�vr�W:���/�t 2�f˳-ЃL���m�s�g��ُ
 ������y��� �ab����^ʳ�\�rP}K��@�:��j�=�a�}׶@��� }B��09Z �������}�{��������� @�� ����  ~��d��֢�Go�?� z�@�7� �ہk[�W��Z�> ������  f�SF�uk�������7��?��� �!@_���  9����2��B����;�{:��"���� K̬*�e�&e�x� @�� z��� �S�i��u����^���?}�����y�!����3z �q���=Q����}� @�� z.�Y �q6��^���	 �����N�Lo <��段��y��Im� @� z*ds8 ��A�x)/K4�Vn׮]�o��% �:��
X 8���@מV�?�÷�w� �@O�)� �i�x�Z#���� z�@�3f�"�� gb�qkuin �@��^�9 �E�k��x�zS%�!���� gc�:� �n����w�Q �2@ϰ� p6f9�XD�?�J����& �e:��0g۲� p6Qd�r�z��%!�� ��'�0�jD `'�f�mo��u�2� ��� �Ud�kF��q� ��DFV]l �eۛ�-��
 � ��'l�� `/�,J�=�z!�� z�' =�5#� �scf]y�+��<���'o��c���# ]D�艈� ��䛺��Qo�_"�t��뢈�s ��뼩kW�K$�K ��@�u�� �W��z�hF�u ]F��:�: �<���ю�	�.#�t#� ���D ��@�u�e�� �gۛ��9�.#�t�� Ηm#�
� ]F�  �:ZGb�8�S ]F��>-�� Ώe�Zi^� t���"˦) p��� ��@  �ul[��:�^ �t�f�8 @�� z�@   �®�| ��@�.q'�t���*���s�����$�!d�wa@� za(/j���������J;AWān��P���5@��(�Ȳ�2 `;M>:��ӌ;  �� ����:#�*  Αm'�(e�O��"�t���6 ���w C�@�}\d ���7w`�� �����U �|Xw� � ���P;�  p�th�1k�A�:�����uy� ��0�
t ���t]E� �KV:#� z�@�u�� �܅aH::���) �Or:��C��:� ·#�Q%�� t]0M p�t��ۻ�t �@��	D)�9�  p���2:�^ ��DFi�@ ����F0�x��A���O9 ��k��V�`0z�W�z�0��8г�  �&���@�+:���}��� g����5 Ê@����#툣" �B?L�et �B���Q��M �� �sw- �u:��	�~�M� �3k7�\�Z<���+�)d �3i5[V]�2�@/Y�`��]nIk_�0Q �<�f���%�@�K:��1]Q����  ���jg�2��!$ z�@�S~��dt �i�-��� �Gt =�j�ҬC ��Y
%!�����ڭ�#�C <����m��L:��28�fݴ�  ��n���^u��sF������f��.� �g5ꍴX�(�k:��k���h�i� ��(ӁXU��9�~ ���� �j7�9���t }�4w ���s�9�~ ��Eg��XQ  �-�릷���@_t������`��M?��9f@/� ��Yk�� í^�'bz;#� z�@�7�E�W+��$ ��	Z~.B�ʗ�� ��@�W�z��)d+ :�j#/�a�@?� ���X�ā. ����k6��X��s �D��+3���� `��ꭂX�@�O:��3S�% �H�Z�ns8���7@�5��8VL��| <���0���]��3�9f@/� �P�Ԋ���  ^�R���s�t �F��B�ZO�KyO�N  ��4�����[�}���JC� ��@`�V�U̎� 0����uG�/4��`t@/� �Q]�����+JB ����l=?���:��#�X�l�Ӭ6�q�� 0pj���G��m�܈�)� ��@`�j��ɕrN|	 ``�~�m��֍��2��D�K ��@`3�ި4FX� ����X�ms�%��:��#�Xg������� {n����Lo7q�@�� �T]����9 $��jq�b����:zn�$ś� ��@`�F���J���r� H�f�Y
���-��u��pD� ��@`���Jql�8� 	��ȭ��Y�����)IU ��@`-sV�Y��ʦj H�z�>b6������w~�x,��u: �U�����S�]�d��0S��Sb��=7�*uT ��t V��HU�����  �2_)��.$�S��G ��t �3#0�B��  !��ƈY�$2q����Y��2� t� *s���ꉖ�s1# �CQ�֍��]{n�����X�G�.#�$B��Qi�fGr �Ve�2j��p2��H�T�s�κ @�� c�����3�9�E j�Z�v�m��v�BFύT�j � � Q�s呱�YQ��� Rfj{e��K]h���5 =A�H���b��� `����M�.tz��v2 z�@�8f�{*�ʻ��� `�f�16�SۗdU�� =@�H���ɵS-Q
 �o���3o��������v����� �$RER�]5�� }���-ϕ�b�厞{��z�G�. �:��2�)[��h��- ���ձ(��7<�E&Η;z^Ѕ� @�� ��Pɼz���Gf�ں9 "�i��\��t-wc�%y7wX �Gt ��zt�l�RH������! ��[A޼A*[���%Y�g�8 =C�H�+6\.f�|C~}�:U��>� @ט���g�^wnFΗ;��0�P*�?* �#:��ɍ�����a�K'.���-ΰ�; tC���c6/)2a�b��A����}� =B�H���_*���a�\���}e~�]� ��*s������X�87J�xD ��t ���2rњ���~�wݖW�ܷ��r�o�;� 	�(��Z���w]뢕�ھ$�
�
 �� �.^w�xn�Wan�d~j�u�/?q_5�" ��]k���մXl%��w/~�-��/ �C:��q�#������y:L�_��:�/{�G:K��B�M�P�/��r+�F6ʶ>��� �!@�l[�U���a4���|�����8���|�~�]��/��L����vcT� �1@�\���s�qZk5��,�d���w>� �9��03?37"�3���m����?	 �� Q֎�����9�DQ��f׌đ��{�{- ��9�|nfn���Ԍ�^w���JOMn}� @�� ����c�Hߐ_?��?<�`[  g�ŝ���=΍nĹ1���|�-� =F�H�����_wA����Җ�pmP~��n" NC���0�0��g��Xw�d��{�> �$��.��\����\4�}Tk)?y�I_  ?��5q���qޭu����Q�V�> �$B6���-�q�H�E��G�� �0#����1rޭu�KF���;�{�a�> �$�9��u��p�H�6�m4~���+,���4����^�����( �': 빎+��xE�Dzm��ϗ
u�!evk7��'������� ��@`��I.�[�� ���B1��L0\"��8�֦pKF���Go��A�>!�XM�����k�Ƒ^]���BS	 ����3s#I8J����Wc�U ��t V+dRʍt�kDQ���8�[�uB������|1)q���O��R��׽�͟�O
 ���j�fU��}�\��:�@���I|���q��Hw<7 @�Z�T�/�$!��c��&dr�o��o7 ��@�uf�#��=���A���r��?���b�Ƿj��)
�M���`��j͑�|%+	a�ۛ�=������6�>#�t���"-˙Ny`��8ҿ"?}�Ou5ҍZ����r�ˤ� I����kc�j=%	��87F����� �3@O�� ������q�K^��H�7�t8�|���U� pZ��ly��jw�
�e�S�� � ��gV"ҟ<�Wځߙ��:nW#����0�R�c� $������HR�Q[��8�D�`�+��@ �:��2��M�/���އ�W_~�v]������Rͱ�;�$�~�|b����ڗ���皒�w�f'��������.7���|��g����^͙��1l�\�g]: ۵����B%#	ӏ8w��G��o X�@�s+�G��?<G����T��Wuf]z&
�l.˺t ���S��L���D�77��ƴL?�띻v X�@�+�3�����������.d]��k��n`֥�Mqԅ� +(��l��B)i�͍~Ź+��p�~S �":��Y�H_�����E�٫~FO'�~���Z�,�
�B��t }����Oկ87���}w��� X�@�W+��v]������5z�誮_�)��Z-�Τ�S���r�<��)�F?��%���
 X�@�w�-�J-��VВ/����\o_��'W}�V�� �/���@τ� 7|���]ڗ�3΍�h�Ю��W �2: k��9�a�W���ke}�֫�W��(��b5����T&�N��2�D�Z5����Ŵ$T��܌��έ�} � �����>$�ͪ��%���Y�'���]�SA����f|�I�XQ�f�s������������#w���/ X��ϒ �+������ުɫ/�^�2��\����e?�h:�cFͫ͑��b��6_bK�;��jw���X��ϔ p�B.C���d6S9.�み�W_q����I�?;���n.�kq���(�pb!���-qn��5�����Y �Rv<[�i������H7;���ү�r��rӕ=�����	*�9F���57�y����R��M��y �� �f.���M_3]�������~Ŏ�K/֥w��0���� ʖ��%��'v��0��&�m�A�}��oz� �� �g.�L�/��t��c{e�� �_~�.�J=M�+��L6f�i�M�<:��z�>R��S�p��y.̶�\��� �� ��0����nw�:'����C^y�+��U[z:B�j6]�����y�M�� @̯�K��r.�皟��Ǩ��w��;_�s���@�� c)�Wb�w?����ˑ�#�'/�Iq�gW��֪V��S����e��1stZe�b���3�|�l��T����'��w $�}Ϣ p���)ơ�w�:_�Ǐ�錨�����#����t�d��\6�ҙt+��f Ι�^���k���nشܩ�H�Պc� $� ��
�r�ů���90�Բ���Δ�k�]�/[iO#�Dy���Z͖k��{)�'�q����NV��R�C���0���]oe:�a�z�S��u_���w�� @B� +���\��ç��=��i�Aȷ����;����:ɥs=��i�㤲���q��'��0t��f������r>B�h/���͗�Bc�u�V  At �_�m�J�J���G�����sOwFӯ��z����_u�Q�����X6%�O.����|�8�̗�(_:�FN��1���l it a��:�K��������x�����n�?>�O�ez�~Ŏ�I:����Y���\:���L�L` ���(]]�����}�������Z�W�`�;v}V  at ��-��^����C�ٳ���|�̔g��;^�7Nm��0Q��v�[>�N��\�͈:� �N�ʵR�V��,���/�E���э� H��{� 0�<�U���:�0�^�K+h-�������_�k.��n����]�������#��p��>�}��k���p�η�\� �'� ��U[��ȴ���rt�زo��'���ayɶk�����v���L:�0������y�Qo�uU��/Y-���;>�A��� 0�قz�^?rh�|���H��7�l֦�ѯ�����.����}�V��Ʒ|'�3��8�u��T����:�>����=8q�� J�%Ũ�xю�� H0�@3��_��rY5����{�QY�c:qH���+7^���t�]�w��ҩT��f��uB�5��ʺº�ֱ-�B��ٕ��/�9��}ߗ>$��D���p������Ϳz�`�S`h$� �azdJ����N����#�w/��̹��?�90���l�O�գ��:���}'�e]���l�W�j��q�j����҆l�����w�uͶkd�0������>��Lg7�ړd���_��_ H8���\O���ɚ�5�����r������%ٲj��v۵�����av�Qw�J�r��Ӈj���f�:p!�sc���5�5)�q_�������DqB��{Wd�N�%m�|�T8u�����. 0 ��, ˴ez�Z7�V�o˞#O���ū����엃��:�ޯ�t���B��"��Xz,=���b��H�H}ω'��V�R���ܦҦ�xn��v���
c�����ǿ�9�1)�8jnd���J&R `@� ��9.�.�N.Z�]�ѯ��h�Ҵ�'g��5[��[�6K�wW2#�*T޺ܺ��֗��f�`�Pt�r\/���)]�T�QXi$;�n,�/�-�M����j�K��/{��,M���g�$u��p��[��o��w �|F��flMgm����C�ȅ�bcQ̆t�����/����%Q��dnR��n{u[�^<"�O�v����*r�n6�l�VZ�[_Xޣ�/(.�+7^a����?�/+��f�%u�|�fgӗv�s�= �@0�����^t�l�ޤ���We�^^�ǝ]��O7�����H)W�$ԣ��ߓM���et��ԏˑ�Q�Y�֪cX�.N{K�
�Ң�k�jޠ��k���w��2S�$�\�3��|꽟|� ��!���GW�׽�u����<ԙ��\f��������t�m~Q�7�;Ui��N�tnZd����q9\~ZNTOH?���T���+��o(��潼��ރ?���������3u>ܷ�[f:�	�k~&ŰX[�Yu� � "���㪫��X.^��s$ۓ�����F:�Ǐ쑽���%�.�Wm�R2��5Wɝ��������X��Z8,��E��s<���&���67���L����u"/�6Q��_}�k=?�mF͍t�
6��^w���	   N��)��/�i���7�ƊM{7��z8������ŷ�͆ub��)���e��&�9Z=*��I���n�_�I�u#k3k
�s��c�Ė�-j<?����}R^��2(an���[���|�-w�P `@� �֍�U���_֏~T��=�CE�<��PvǏ{�K:��Ie�6AJZ�eSi�l�"�vE��sr�rL*����UH�Ԛ��tn:;��H�Jm����1���~���׵��e:���b�����c! 0�t 8�q�/�-�6�o�����mlvP��S�#�w��kv�s��zU�QER�R)�ֱ-��~'֏׎˱�L��CzE�S�)g*7���MeF�#^���5E��w|�<��C]����~:���o�ݟ�]�G��92����W�L��Γߑ��V��zT�f���kw�e.�b�(�2���f����j�j���b�Y?Z>*��%�JK�)Y5�J�S2���ԙ^:y ��?�Y��ȡ�];rm����j2�<������ � � �i�ȴ��*����z��2_�_��6k�M��~�Q�:�E��p��TJlfb]���c2�.��Tʭ��Ʊ>W����\g�<�B��%YU���8��sc�<���J�I-��w��=�X�޸2ann�2��T�z�|펫�^�F `� �nT��/Hy\���u�߼�u���O�w�>���bfTp�̾�m��*�j㕲ab����2����ݼl�$[ƶ�ٟ��We�Y�c�ǜc�	��3Ȧ�2Y����L�$�������+����̊Y�#Og�֙?W1,�/��v�Ϳz3�S:��[�[�#���^� &�0V;�^$[Wm��-�u��|%͔g���,�q�t�%�}ն��<O��3��Y��5��l(��+O��Ͳ�9�:V9��ͅ!#�C��)�D~\�� ��OH��J�(�m���c�և�wf��?ڵ��=̍�ε7�ֿd�n� "ɸ��hw�|�ܭ�n����'���� ��ԋ6_%�ۡx�Ay��c+>jf����o�{�'�M�K�^,�\I���
/�xyU��Bnsa�V�D�Vşo-�q��N�f�Z���*ù2���f'
2��yJ�N.�xƩq�A�wfҘS���a�|i:� �D�p}{���ڹ�1�!C�����C���;�{���7[nk`�{r��z�E/�m�	m6�z���+v4������q>�l�� ���D֍��~���DQ�$�h>�����Ƣ��Ӂ�r��[��\m.�k̇u�=q
�����d$;"#��7�O�?%y��\uN�)�{��]���07<�Ee/��;�sǽ Ch`/��烷|�{�?xݞ`�o���m5|�l*����b�|�e�P$�镞�n֩?5{�s+e��c��h�E�K�$��1Ym�7�48%��*�J�M�M�s]�k?4#��v�5W_ˍ��֪�$l6��ȸ9u`$7"�TA��b'�Sf��)��:J��-��@gm����~�a
s�ю��l��Λ��� C�@�Sw�z����7���O�m��:ҍgC}����Ïv%ԍ�fU��=���tF��Qm���%rT���({ی����#�H*�����f���_�G�v=�������F%Zl��Jk1b#��ȧ�R�$�	���)J)S�D��1n<��IfF��yB�������S[�n�;����[�[ `�� z����}ۇn��=����?�nd��N�_��2m���>�hW�\2Ǚ�}�s�g�}����MF�2HL�G�D{Z�^����
��;��N�
�aկ��v-��5��X��vM�A��(H�@nW�ݴ�ɥr��rq���x!��8��q�ɑ���%m�z��~y�ؓ&л���1�3r�=����o��� C�@�w����f"��8��C�F�3�~���������>��Z�����zgWys���m��vn�TFճ���)�+�bg�W2f�=΀��C	�fЊ�a��A+lFM�L���o�,�<�#��J�MI�Ku>g܌d���AnvO7A��o�r;���Kn�~\���0
����c{�����R�n�]�����E���|���?   @��H��7�֞`�_N0TCF��v�g�(��=��������}=�V�ܾ������[Wm�L���H�x7w°3�'�Y#�.�O����`��V��a��~d>���{a|O���#hK�ݔV�6?.���n��rt>�s$/����S�
�vMx���_^����H��7��'N�:o3~���	߸�Bhis��ޙ}b֗w{
�����as��n�#��]o��i� �@_�z�G?�oj�	��ۖ����%�|����������&�5jF���As3�!�t��'�wFW��٠.��7G~=[Kf:w�|�����9��DU|���7:#��~?���8�M�ǱG{�=~�����i/�Q���2��3��)���ک�~���?м�b��I9)e~�\'�>�R�g���I�W���LD�p��Y��}q�?5����޳�m�܌�3����-�� �Y:��3k�o��������o����}��Ҥ\�O�K�]#�-Oy�+�ԗ�s���߹��3#ꛦ6ű�n�F�/�	b�K�O��?�3�'�.vX�磟Q>���OǍ�h���mw��n� ��@`�]��u�w����{�o�ʹ1s\�9K݄�����ӏuu��a�p6#��fFi׎���q���� �Y��3Ǣ�?��̑C���=��ü��tҒ
���ް��]� ��� ��?��?p����߭���9���L?77���9����꨺aF֗����X=�J�Ol��e�0&����>8w��G�87�{�i�ϗ�2���E�t׭��  N�@`�]�ܵ��߾�棏��
5������t�K��/�٨�a�q]8ֹ}w�w;��f�����ck� �e�g�������Oˡ��2�8חc�-?���7�8�^q���  Έ++ ֹ��;gv�ڵ�[���9�f7�u������އ���1PK�ͪ<��c�����ℬ[ۙ�zt5�k�3�Ƣ<�p�3}݄y�v^?F�_�x46�Z�/���w �"�X��o4�7��}o�����/����+��y�@7GfE=�0�|]��=x�α^k��tF��ı>�tx��F�.G�f6�����f��?�a?"�\M�_���mozӛ| ���j���3/}����~.�Ô�$X�Vkn��uì�?p�@�fdSY���U�6�J�JS��㜙 ?V����L帔k�L[?;��;��k����}�e���[  �@`�O�㓯}��r׾h�[C1\���a�t
���n�K��i/݉�8���ȔL������F��W����	��c܌���@�Q~��_-�,�ۧ���+ ��B�H�?{���v�o����M���s`��L�7�F���Y#l6�2���/�ɏtb}�4�9���:.�>��?��zYfM�wn�2�y��9����Yz��ǋ�h���?��]�Q  �@��޾�����_����ߍ�Y��SG m�u�LW6�fnO}��}�rd4?�'K2Q���ℌ�%奈�2#���N����;���|_7t;��(g]���G�֖Ԧ_��ֻ8F .� Qv�e�7��u�ʣ����JS\I�'c}�E]
9���nF�ق6��渹��O�w]�����m�Q�J�r2�kq��!^��m˟��a��ʙԓG��̕w��9 \0@����;j�o��������^��r"��'��`�vs���:q���7�^��}$?"�숌ƟGr��6b�>�/�?+����#�^�J��	r3��X�j��a����J�zw�7?s�=� ��� �����/��#7��[�o����v=FS���-��#�&��Q['��z�����q�u�R������/şs�Ph�g���7Bj�ڳo�,>����0y'e1u�{<�F��mw~�ֻ�. �A�H��n�����p��,��W��_����gA���?��$���&i��/�B{"xԗ�Tn�}D@�(�&;�� vY����L�m�JD�B�E�J����V�T9�s<؋�К�K�dwv��3K�B/I��>3�����y��ln�$M����g�-[��W���Ȩi:2��<���5�}>|}��i~n1��%=K�b��z��8�v��Eq���{���4�\�陃�`�
�������c�����?w��>���ǸS�O�%y�z�s_��\�� ���@�۱y��v��9�w_����]p΅g�<���*EG���p��v:��j�ڛ��:�Gy�Bތ�޹h�	=���M�Bw{c��7c�����sc\���ͱ�}�V,v�bv�^ ��S?���L��ç�7��n�7z6��;�=�~6�O�������g�����xs>��F{D��9����'X��������� �Wh�֭k��S�Y�|r��=/:��B�W�'��#����Ճ��4#��G���pd������
�����?�k� 8!:�V�)]=r������߻�sO{ʏ�,����I�H��*�ē.א��������g�����? �0h;׾g�ߏ�c˿^���5���'�z���O����m�k�Y8�<-�K6�V�'.~�\��u�}M O�@��x6�<��9�O^�_���+�q�3��-~��Vv�5�#]�w�#OSw�zz�]�s���~��5���G '�@���#��ݕw_��[��\��5k��� p8Ď���7�Ñ���xkX�/�}Z�n��% p�t����;�v���;�;���]t�E�ȥ瑎�
���x�+����3n�ݑ�/ �t�;6�X�aˆ_���}�S.^��P=��G���w��'���!�~��e�Wg+_s�ȵ� ,�t�m�����ߘ\����}������b��.Z�Ý&��P?2ڏyx�G�O�q� �H�3����|��}�_�����ڵ���X���"����������F:ϲ��=�V��Qs�4t�c]=r��������V������c��b�R���G��c����_���١�ͱ(6
�3�3����� $C���k޶iǦ-���-�?��矶f��Ï8:|�0���\���ҵ��G+ H�@������p�;�����Y���~ړ���׻D�m�w�w������� @�:��{�u��;wn��_�˥k~梳/
��M��U�|m�����,y�5C��	 $K�eݺu3qx�Hu�y_��Kv��O<m�Z�����~ja�k�F��& �<��&K�7�a�;޿�=w��|qoo�P�כ����:�w��|�P �et��pݻw�o�Ν_���O�8c��/8��N�ԕkkoY�d�˜��z:�18t���F�Fθ�޿�i���\xޚ�B�����kU>x����%�]y����$�������qx����K��o_��9瞽����E:� ���+�;m�ڷ�6��2 ��:��P�8��qX=49�kw��S}�yO�_!ԁ����d��]k߻�];*�� ���������'._������]�ۿ�_�'̢�w���?���׾5 �V:�<�1z�{��+o���GN���g>�kq�"�̛�0/���.y�뇆� ڎ@�'��x#���^�ƶo�~���7\p��Kz�u�q[�譟Z\�ً�\�Za��:�<;�o������}�=˺�(ԁ��;�[_�ü_�t
�p�\z饳q���;w��ڭ_��╋.��l�<�E�E3k��~�����C�x�Ct����??w�{���]�j��9����>����Ƣ鵅S?�㫞�K��3	t���Щ�oknלּ���z��8�����йB�C�v��Ī��_;�� J�,�k�׼�R���=�o�{�]a���郧�B�:t�B��`c�۫z�su��?�{� �p`�����/L�����%k��9���
� �����X��������}��/ 8�@H@O���ׄ�;g�7���г�7�yڙaq�� ���3��dk�0�s�/n-�� �at���bX=�*�{C���w�����3N	�,_���%˳�tv`����_�i�e�/�t�D-͖��`��<n_�г�7��������t�6z�+��^ճ�׫�~y��M �@H\����W�����/��K�/�������cꐊ�Mߖ��XU�_x�7^z饳 ��@hY���a0�=!ܳ?��z ,�����X=�������O�^u�di���{�� <�u�ך�)aM�)aw�'�U�+|7�/�3��D+���`X~�`����ӵ� ����eKò�C#�aW|�5}w��lW��0_�n���߳�{�sK���Q]_�w��]�<� m�y쪰2��Yf��po�;យ{��=���8>ͻ<��}�W�a��wԮ�}# �	$��P1/�Ӌ��m�랙o������C�:<�,�7XQXq{_X�yǻv�U ��D���E�u^���pn�)�ý3��m��{�N��Nw�H��l�7�������? `t����
gϘ�f��۳�����v������Ŭ�/m�Y�-����� X`�C5�V�̹-��p���s׭��v����n�w__v�(���I_����= "���C�)��ᔞ�!��'�ߙ�N��Ʈ�`�A7��%5O]_�Xr`Y���,�^���zΩ �(��ɲ,,Kò��s�����w�c��]�@�7��'t��7�w-͖޼���7�._��� �����ʻ��2��^9��/<?�����	������y�l�ށ�ү��\35��� Z�@���_��Ϟ;���CaW���+ <7ׯs"u�]ai˲e���&�9����/� �t ����}y_��~f8c.��
4v�E{�Z���s���j��Z�XԌ�0X���aq|rw�T�2 @� ̛fP�a/�`�9s�����} F�����f�e����g��|�@��faE�������� �St N�ft�R<en��|K�\���+^r�1����>��ƃ�=�u�o6���'�K�kYai�aYqiX�X��� �K�p�m���8|���Ν;�o�}��y��]�v��e��f�����VVȲЛ��_�׎��_�����  O���֭[׼�܇m?����{�s�[6�T��f������.ٞ�bV��E�/�x_�/,-���-�Ǐ ��: �z�[��oqxߡ��<�����<8�����=��.L��d3E�~b4C�'���E��Z\XC|`���
]��N�X�c&�h9�����C��~�/����gg^ppf����gN����P_<�8�;�5[��w8]1���ߏ�lQXRX�dK�?/.	]��G�F܊�&�h+�_�=�?=�=���=��C^P�ן9ݘ}R=L�����0�Wo�,���=�a��^�Y^h���5���sa�sī�phk����Sh�zB!/<��q 8�: g�7&�5������nذ8�;?����������3�~�L��j6�/o䍾P�{g�=y1m�1g������Bb���sc�1W�͏�� 4�K��'p=�Y��(��,���y�P���5�f�V�*t�;�U���݅�}py6𪮬;ď��!=~<ŹHL��� �v: <�m�n���mIںu��F�񪹝<����s h)    �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �    h9y�� �f: �r�,�T*}�r��  mB� -�P(\�[ �	� ��F��� �h# hIY��*� �&: Ъ�^�V�_*�� �t �e�y>�@[� @�ʲ���5 @�� ����z^(B���za*���X� �0� -.�LOOO�T1̟_���� ��: ���K�<p�@�dy�oߺu��6n���  -J�@��������Y:T��W����^��s�; �J�@��W�������b��<��eq�# @� ��<�/jG�![c�ճ�hE �@��;�pA�pq��<����۟y�W|' @� ��)n/
4#��z��'ccc/( @�� �b��S��7��;00pC��W7�� �: ����vI��ŵy�;��
: �����ۻ��?�M�j�_�xe ��	t h�7o~�R�ܕeٙ���7c��T*�N ��	t h�=no	��<ϯ��j�2 @�: ��,�>�ÊkSl4T�V{J��G $H�@��)n��?��y��R���� H�@�6Q*��V����<�C���Z-�> @B: �����*�š��?#=�t R"���|,n�<��G�+�J�\.�A �t h#16�)F�Wb�>'�X����~�Z]Y*�� �@�6��������š#}����減 X  �̒%K�h���[cl���h�V;ull�m����  @�@�Y�~��J����3яכ����7 p�	t hC�b��h4~9x&���������HU��= N"� mh�ƍ�W��O���맦��??11�s���� 8I: ������*
�<t#4�C\�/�799y����W � ����譕J��8}Y��8�P(�M�Z��R�tc �L�@˲췃@"��g1�%F�G �@ �X�ʛc\�I��&�x��y���J���r�� N� m�^�_�����8]x\]�?V�V�X� �g �ܦM��aY��+O�[���s�����<���&��dY���\�8�xB��xff�[�l�dӦMw �' :�����J�R��O��Ӻ�������r�� �� "��W����?�ggY�Ÿ��,�J_ �	t �,��<���k�aE\Ͽ�T*����  O�@�R*��V�o��O�E�e�1�?^��.� �q� �ab��Y��?��7�E��b���u=7��  ��@�T,/���}a���O��J�߾}����7 � hÆ߫�j��h4��y�v`����l```���؛b�� #� jxx��J�R��k��c�b��Q�p�: t�r���Z�>;��D���;w�|úu�f <� .���Ȳ�qzQ`��n�޽����^;44t0 ��� ������j��1ԿC}y`�]233��� �x4 h>z훕J�5qzc�z�����7�����5� <� �)�˟����,�~/0�⺾�����1��#� x8 ���#����.����<��8� A� ?d߾}�����'�[k���8n p� ����וJ�Y��w�8��V���J�� �� ����k����y��q�?N��W*�]q�?  t ��xi�X�b�=7p"옜�����ȧ O� �htt���/.
�H?50��,+��c�J�g���� :�@ ���ȿT�՗�y�����mI\�?ݶm�s7l����%���T*��qbb��.�wW�۩�z�/��ꪟؼy���$��c2::z����%�B�Ƹ;�WY�=����O���^244t0 �q: p�FFF�\�V_��	"�Dx����������#���R*�n�����,�>�����k�˕J�o���u��"���622�������"���>11q���� C� �K�\�|��`1қG��&�gw�P�d�Z}V�T�+ �: ��H���/�������&�皸��{����C��'��'���Z��3�F�fT�M\�h^��� @�� �6<<|����='���|zs�R�B�\�� @[� ����1$��eY�9��M\����722�� @�� ��)��w�j��5���ݟ�/��z~lll�ٮGh_ �W��û*��K���q������~�����8}{ �-	t `ޕ�����^�������̗_�V�]*�> h; 8!��ǧc��R����H
̋<ϯ�������ȿ ڊ@ N��8\Q�V��r[�,���%\�?��~��K/� �� �p�Ri�V�=#���0_<qϽ�;��c- �6� 8)�����T*��'�,[x�޿u���lܸ�� @[� �IS.�?]��~&���wW�,�z���;w�|κu�f -O� '����W�n����w�<�ػwo9��9 ��: p�5O˞��x^�XlF���[��W�j�O� hi X�����ر�'8��{I�qi��޼�����s�5�%���~��}7�pë���q���׳���~5� �,� ,�C����j��M�J��m�T*�*��� �$� $�g�7���K���vq�� @K� @2=+��8�/18��כk���q�G ��t  )�r�s[�n}~�����{V��5/��|�Ν;���� �G� �i>��V�=����؜?8�޽��8n �� $ixx�ߦ��^033�ɸ���1+
�ٶmۇ7l�� @�� @��������]��߿#˲u�c��^�o��h �et  i����8�z�R�V���c���fו��; -A� -!��D�{��a���x,������) �: �2b�drr��1��8�U\�7LLLl�5 �<� �������j��y�|����)�ū��� @�: �r���oٶm�O�����,;=�h^R�V�W*�n $M� -iÆ�#���"�I�G��y�� $M� -+F��NNN�d����+���U��g�J� $K� -mdd�ޫ��ꧺ���"��s��Q�� �%����y��&&&^R(���������[�^�q��� I� @[�#��1�?c�y��fgg��7 �$���ь������������?*��/lٲedӦMw �#���244�'F�˺���7���G�*�o����t ��lڴiw�����l�e��ק���?44t0 �� ��C���������s�,[=33Ӽ��G I� @�jFz�V{Y���=�>=p�eA�$G� mmxxx����K�����e����nݺ�?mܸ�� �� @���V�]������)�0;;��8t��t �#�����
�����B�˲�ұ�����ǧ I� @��z�V{M������������i? H�@ :������T*o	߿IZ!t�7��� t�r����Y�]:X��_�e˖eͻ� �@ :R�����yq::עb���8~$ ��: б���;200�8�$t����� t������������q�?��e�O�ر����� J� mttto�Rye��cuU�<=������fq N� �\.�Z��R��E��;��l� N� D�R��J���Y���?� �@ 8d߾}�������/��܉��GGG�g `�t �C�7����z����W��i��dY�<�]�, � p��������[�<�1Fk:D�P��8l ,� p�R�tS�R�.N/"��g �@ x���xQ�^:@�ek�l�rƦM�� ,� �0���������_�S��³� ��@ x###_�V���_�P��I `At �G�e�H��xeW�6�:t��%� ����j���8�`hsY�=# �`: �c8묳���;���������j��� �t �1\z饳�J�q�����<?7`t �cP*�>Y��6���C˲�8�C ��  � �k^�T������A`t �c���s���t����.��@ 8FCCC+��G�ڔ#� G� �,�>�8���7 X �8�V������� X �84oW�V?�o�I�,� p��<���m��s ,��@fgg����j�/�I�P�F��pOh_��,��@6mڴ;���eY�z��zw��ٽnݺ� �I%� �S�T�9���yw��ѿw�������o��@ �\ �E�_�~���y6o� 8�:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $@�  @:   $����$%Gy>*    IEND�B`�PK
     �9s[	^�G�  �  /   images/9ba3df0f-d630-43f7-8169-617793654d93.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  sIDATx��	��yǿ�sfvv�ОZd����XĎ�;N�g[(���p:�w 
`'X�B�1�������#��:@ ����c��9��|_Ϭ4ZV�EB=5��������]������Z�JU ��
D0U��*�T"��@S�`�LU ��
D0U��*�T"��@S�`�LU ��
D0U��O]�f���� 8��S*V���F���!�=�J��@?��)�������w��ςfܤ��%�c"�4�w�������|~R�o�p9����ƽP	Ȣ'���y�q/����;	+��j�����ܬ	K?��`Bq�� ���}�|a��Ȗ/�p��W��i�>YB���E�h4�nmlj�'��<7���M�ŏSV<��G�Y^�O	
�YNg|.~xE���#�5X����0�~n!�����AD	�o����9t'{@���S�v^��G�1Y���eC���#<����g�����)��>���=n�lX��"!���@=��A����R�󼻗�E,Ə�Xl,�X�� Z��JG�C�����F�o{�#3�e�u �������ֲ݀cG]wh�|],(er�Ӌ��M�}��/�}7ƅ��#�
�Vl?�E���ɍ�:�������lu,�reI�p���,i˵�OK��DKy@ K)�eO^9%[���:_��
#e��>^��?��� B��N>��ke,RW[Wbb�D��=�~D�b"�����;��N��*����Y��
+���a(������ ���j����gƷ�ho��l+�2���%y���l0On�k�7���xRKJgM8���f��n�z3�$�*�riC��u[v`����=ʭ� Y�fq�-����ƹ��2|>�i�>��+��
�j�.����dw��
ZɎ��;��v6LҦ�N�k��(��4�X\�K��|=���ZR�^l_�0�-e�6Ct�Ȳ'�AF͇֡z�El��-(��S[N�u�vQ��Fˀ�s�n{5Gq[O���n�{����g'�U�P�kB����;^�c�� ���|�����;�*�P�W^�9ʶ�$ M��� Ŝ�*lR�$}z��8Y�P�]�5jB�������0@s���D�\ܾ�>o���;���:cg|MVY]�N�V�����h��I�.�-^KE���v��P����r"�*�!ޠ�l��m��S�܏�|�-/��g��������9��Zb�<eh3�t��+��֒[�f	�7�|Ic�@=�z����JZ�|(������=t-�C�~��ֆ=M
ڇsY�E��������`]��LE!�����PNE
���0v���X�!�NI�H06��dmؽѤ����(��a���O���1��~+R ���i쭉��
}Ra��q�:+�G�"3�m��޸�mK��n�cyh��`Z.n�@w�梧��}���m��^�º7v�ɟ�oy��!���S0��܊�������1�A��N �ϣ�z�K�	��s`�O�
=�V�ͩ����RwEV�u`�CA�p	�(t[0Ǖ]H8q(�"��*X��j?�7���q�F��QEր-�`gf�C` :��'%�DƲ�Hd@�?����(�
L�FKJX�����i?BQ>��3����l��,H�5��*L�TIe�����0�9� 3iN��DBwʺ�L��F���>��Y@�J��Ѝ�%��d�NʨȀP@W=� �R͜C���S�"�C�Y˕���R�`���x�$(�0o?l��X��N��;%�u5Vܷ�)4pB8�VwG���B�B�T<��A�kyI�h$
��vʵܸ$K~�9Ս�*��ɶ협1t3c�y��Z��sT��$I�U�	,1�ൌMb�6�V^H�]�c��"��D_q_��Y),���<��u\��<Y����?�ӌR�a'���AH ����%�����D/�$kpL'a����A
�ш``�ɮi���`���/���O��� ���lL��8ʵ]=��7cs�U���>�Xڲ,	�SL�X�V3��TI0H��A�4)�A�ف���P�(�8U:���R����4O�.������@���stS�讜p�R���~N�C a���}� �1TS	�� C
a����s�3˴�X"��Uv=׃���5���^��UV �uϕ8r�-&3�5�|K�1,��C�ـ�M���ޡ���S�zl�Q0�@MM�-�i!'����H��^���2���D���
�V�⺮$�Cs7P$E6A��᬴Q�P�@��_G;�ԁ���x1����ZMm���Y8�8������6&��iy�VY�Pm���]8T?	��2�d	����oC��y3r�JP�@Ё��j���/l��\x�E�۟��)��g����Wbeo��R۲�XL��r<��mnز ���bю����x�TtU�p��Vn�k9����凶�0��M��c�1M:��)�u�m��sgI�e��?�D������d�df_|`.>�:��a�w���8"B�i�f�3�K�\��?���R��Xp.�W�|	a|'�Èn\��C2U�l@PA@�K�(�i�6\���y�I$�Ӱ`����c��ޒ�(h,��M{�vWmd��qa����ވ�K�2Y��,g�i�1�塐��C~G	�RG�pe�Rd@�����EX�/�H�<��b,\������,�rP�`�A�.����0s�#������!*E�ʛ@)�k;���A��n�Ƒ�W]}}�0���.�L�2,�G�����G�i:D�%)���[ x�*��UEWt
��ذ��.Y��O���(�G
d�;A�(ad�5)�.+
�3o�=���[G�#!�����X"B��ѐN�ǰ�X�! �������u`����oow[ Ƣ�y�v.�<�j�^���!(�Ԝ�Q�����!��B
���*�`Bt3ܢ�\t�p���x-t�t2��:��K�E�1���C}�u̇`H��y���&A�Gv\�Q҃�pBm+��<���->�sC�GGa���AD���\O��gR�?�\pUd?�қۂVx����"�\D���R���m_3�Ϟ:���p\o,�;LV���'ue����$��5*�D>�K� �`��
��K�8i�{�b>�3y6�������)�;��l¸	��[2�Z�ף~%Z�/�v.������O�
��y���t�b;{v&<���4f�!�Ӻ� s�	����q�6�0�P֨��ul��Y���7���~���[a执��T�ڤ5՞9��DO��A03���
g(@�s��nA4Pb��Mz������ښl�u�vēj���_o�|���)�n�Ӽ�u<uc��aYx���nߒ��!\��^}/��ϦT�;g�ɭ��ֶu��ͩf8�����]�L�0]��`r�P2v�3<�w|'\���T$�������0�Hh5P�Po`)���*?m�a]�:���{��
(���hgY�$��5�Utk��b�����6�UAׅn)�!O�9�}���Aظ�mxi��ɂ����7��q�qjKc�J�HhQ�a�<�(��h�Sr<i{�Î��|_f_��?Qu������w�݁��&�������}��S�)�ųϹ�˻[Ͻ[���
D� L��4زwd�,�w�oc��'c�6�YBK0]�hŸ����`9&�<62�5�`8F�n#Y���~��TXs�������ƣ7<�Pd@�\~'\�����`#<��0��y��_O%S��;�*��Н���h&U1����r����h��X��s_�-�"@Vd<�O�~�t\+�������l�����Q(�"�߿����۞����Bx��o|�G+?����<���i�6ih���J
��я�acyL��(磓�7��7?�TY��z��Bz` &�8	�r�7}t?���l}����lk�Y������Q��=�vc#�Y���9�o$���� 	������%����*ҷ>����!�u����>��,gH�`�>�y�ǫ�?,��Z�F�� l>�-�	lA�<�^tf����0#��|ӏ@�}��m�����x�� ��a��O��@ ��&�v��0ض��.��	Xݴ�S���Dcz��$l)A��!ɒP˒���d߱�?��ҙ�,x�} u2���Tv #)(�kL�L������̻������0_�D�m�6��L���@���.����1����BK	09����A�T߽�@d		�T�~�9��$O�t0I� LʒMফ�`�|������a����o1�~*A�)Փ7>�����ܨ�)l�UQ@�?�
D0�@ȕ�-7rm˗/�u� �0��)꼺�����/@�X�B�N�
,�a	'x���PW#c�����F؄\�cXh��7����t�RM��n�;�K��a3:χ��a���p�hU��uPG$j7�+��=�����r+��}U<�e˖�[�`�+,��'�`����!��A�x $��(4���x�C����G�z�q�4������y��S�_��L,Y���B���yXh��H3nN�Bͬ;DZ���B�~���X^�2Ҙ�+��B��+W��k��ʭ�i�MX.��+����&�W�<.����P��xn�0(o`�ˏGؔ,�qD��B>Q��͖���J��[z��*|:��
]����@�A��.��1��;p�3�����i��װԖ�_:�}	�����)a%�c�,_.V��hHUT"��@S�`�LU ��
D0U��*�T"��@S�`�LU ��
D0U���W�cfrJ�    IEND�B`�PK
     �9s[U�p�	�  	�  /   images/42e39361-2f02-4030-a678-a3271aadd3f6.png�PNG

   IHDR  �  �   )��   	pHYs     ��  ��IDATx�����e}���}�m���N�s�	!"�UD�R)�-D5t��9�s�N�ҩ����L[�N;��g�t��3gfN;ө��V.RDQ	&$B��U.I��H�o�����jEd�<k����Y�, �F�k��z���   p�	t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t   ��@  �t x�kC��m��T:Y�YQ(dˋ���$���4)�'M;�$Kz�&I�����Wz���?ϲ��eI3�餓����]���C=��~�T����v�ggó�N�̒%#�O?��f  �@�!�B�yr��=�Ph_*��-[�BgA�Ю�J�z�6�i�`�h~��<�F�]��t�S���Vi{�Y|��L�v���]�_Z ��@`hm�z]��x��J���r���Tj�����X�]\*=8��-I�\��+���Bc����?���������fyo�Y����F�x�[����s�I� �Q'�
w�q���+��V��ˍ����B��������Q����=�}�s�5���f����j��u��ے���  ������ޫO-�����̞].���uE�>yT��ǫ�V*3K�G���=����3�<6��o]�cv6��ʦ����/��  ��@_۲�ݥn���W*��j�g�jS'�J�.�,�B{�V;p�wV���{���;Ϟ���=:=]���L��'���q�7t pDt ��C�Re����ڋ�����FF�>6M;���+���g,X�|���sk��>��o��V��,}�'�	v x�: ���������5���E��w��hQ>���PhW�����?�-����#�\���TmӾ}�.�覇 p�: �ٶmCyzz�򱱙+k����jO�Ȳ,����.����珕+û�z�=���[fg����}ڴx ��: Qز�]KK�}׍�M]Z�=tb�v��m=�}�;��.a�e���x䑟�Ɓ���t�G�<�CS �����/_�bE�����k�?�,�V���.t�;��㏿���~��g����n� : �l����ΞkE�3�5�m���7/���O���<��8p�vS�1���L �!%��s�_��p��gll����N�R�w�i��p�޵���)��C]t_/�?�v��7 2�9s�W��ti�����Tj���+��hў7��������-�ܾ}�?���� 0: Gԡ���w��=݂O�B7�"�J3��/��vٲ��<r�_<��Cg�y�ǒ���  J�pDl�|�I���?��R�� ��$��w�n��;���m�.�mϞ�zӛ>�x �#�xY�lY�����=:�詽?tW9s�T��W՗/O����o�o�ޅ���s��K �@�E˷��p���[�����Z}bu�y�-|g����ַ��Ԟ=�������3���w��v�]��~q��'ޙ�p��j����{����k_��SY��ߟy�ܫ@_� �D_��[_�l��{���,�� 2����+�������_�m��c��v�'w �#���/]qҊ��5>������ �+���K�����sE/�?�o���\p�'� �: ˦M׬^�p/�w�9M�~V�wҴ]���/�u�7�q���]�[B��y����u׆c-���ŋ�uE8�\�v�K�캬�}����-�n�>��K.�Ԟ  � ��n�z�ʕӿ�t�#W�¼`�������.ݶ���<�d�;��}�@ ��t�!�u�u�R���/Y��[�9àPhV�/�y��xy���_�������	 �0�����_����\,�.
0dJ������_\��~��w���sι� �2�0d6n���c���۵���r##S�7�?��߽w���}��� p�t�!��[�x��.^��M!dI ��^�J�~�>x�''W��ڵ� `�	t���C�T����o._�ȵΙÏ�-,^�����]��o~s��;��|� l˖+7����E3�8,�bst���^�h��[�\��k�~��  �@����Y�lپ?�Yf;;����1k�<�?��ok4V�ʙg~h* �� &��>1���S��, /K7]�d�e�恍��s����7}, �� ��;�>aժ�8:��kpD�ˍE���z袷8��"�\� }.�ޗ>����Y��w
� ̉��ȢE{�;�����_��[�k �#H������5O>��?��8�� ̋B�Y?昧��#��i���/�ŵk?�3 � ���֭W��+�|O���4^�$YV(�+v�;;��3�ڦ����^����{���g�}� x�:@�ٲ�]K.��.|�� G�t�\>$O��Y�=��t����n��d��^�k��Ph�֬y�>x�x��O.��6��x�:@ٴiݕ�V=���� GH�M���@7IBH�$Y\(���R.���1��z��}�쏷�����l��Ż.��kwl�r�?wo: /�@�۶m(��.]���z9�^s��|��T��G����	�T?��?�҃�N���wY6cy��R�^�z������/��k^��%��}���"�"��}����&�0G����N-��M��B����Qɷ�w��v��GZ��C�^�u��i�81�����������^x�c �@�X>nb�_I�N)��vw�_�ߙ&i��X.��Y���j=��t���v�m����O<����������9��xK �� �"�e˻K��#�t�S���[̱nwo7˦�IRK_�N~~�\>��9#���N��p����P���J���{�?n�v��N?��� �'� �ٴ��K������NȜ�ee�3�$9�����4]Z�=���y#��V��v��V�!���˗�����������ڵ7� �:@D6o^��ի��w�RcA�y��+������$I�եJeu�\����y���<�l��h��m�=kdd�����p���? �� �"q��W����O��|�T����}�%�C?|IRI��S���T��i�h�Z�Z!���+���V=v��-W|`��[> ��xp�m�z]}t��?]���sE��s�,keIR���i��P._T+�������֖Ơ߱^(�G֬����ח�u�i��Ul |?�p�u׆c���p�z���nȲg�I�z^oH�rR*�Q)�^S�Ϫ7�[��Σ�����%˖=��G���7�|�Ϯ[�� �@8j6o���ի���Rifq�H:���(]�w�����R����j�3{h��`��Ͽ�կn���/�ׅ��d `�	t��`ӦuW�Y���U(4�"�e;����H�e�Je]=?��j}��n�����ju�W����7���.�� �P� �l��+~qbb��G���J���y^Ρ�$�9�J�Z�|^%?��nokfY'�r��������-���ڵ7~* 0��9�G��鿞�x����(���f�������#$�X�\��Z����ln��כ���=w�O�ۯ~��5g�u� ��~��m�6�K��:>��"���.п+�C+�g�B}�l���VI�-{��������N��/ �N�?|ɖ-�j;?6:��� } ���k+!bI���W�K�״��;g;�gb�{�e�ҥ�^���/<���Wװ�0�����-Y�������Ng{��ǡ��?Sl��v�gپ��ŋw]��#wܰmۆw�~�� �P� sd��k��^��'�����H�MeY���$�/$I�xB�X<��jmm�Zw�� ����}�@�ᡇ~�ړN��F `�	t�9p���^�f͎�+���P>ͽT�@��BR*�=R,�Xj6�i�뛝 /d����=x�ܺ����y懦 M�a_���w����|Y�>u����Ї�dA�Ry�h��V����,;������������t�mW��K>�' 0�:��i��N[�zǇ�{���nwG߯>�[���+�Zw϶�_m���z��q'��}r��k�y��|. 0�:��q���{���V*5G��nwo7˦�IRKCK�RR._P-O)7�5��<۷�^�M�Y�z��k�;�?�����#���{��ԕ+��I�(��}���	}�ߕ�K
##׎���juj��>��͛7\u�7< (�eڼ��&&���b�� � �vw�C8�ơ!r��+J�Vӟ��JχO�^s>v�]�v��7� ��2|���׬Z��#�RcaIRM�l&�C��O�.-����h~6�ټ���7�&��q��7l�z��Lw�%��9?�؝�W*3K�P(&��*�ҙ�F�3S���2���y�,ke�9�0p���7T�����[���`�Uz�~�����[o����.�M� ��l��˖=������0
�W�*�7U�d���+�+j��G'�Ab��Y�l;IV�6������������L��h+��z}���zU��m�~��74 }M��H[�lX�t��V�V��y�|q�X|�Z%Y_����d��X���S.n�RͿ�k���V�3�6@nll���n�^���s�7���� /­�^R_�d�'j����X<�T�\\�c�G��$Y\�V��ff>9Տgx9<����f!�����%I�tF�PX^���y:���7�{^�ɟ���� @�� �)�ޗ>��v����J�zR.��V,�WM���R��Ƒf�K�����<ݞ��oK��J�]�I2^,M'���ώ���6��<�W[�/�}Ѷm������{ }I�����K��]X�tj�T���$��^--���v�t��v�u@�Ԛ�͍�Q(�*�g���K���0��#W���Vk�l￁�/V�xf�׾v��׾�� �;�0|�k��wɒ����$��O��������rq5��w����@�tv��G����TzM/�O�|wx�`I�r���4]�6�΄��Jϲ,������{�c�s�g }E��w�}�;V���À*V*��kI��el].�]mf�/&���./M�Mg�V��4
�S���ٕ|.A0��	�4����짧��{;I��c����M���q�y7� ��Ǹ���oX�f��	�;p��{J�sG��s*Gb X��ґ���gf����Xm���'�����7�m���J�.��i��P��k�Ѹi�_v�
�5k����o_w՛�|���0P?@��;�������Ӵ���}�,I�I�|y�X|��>+M��;������.GB���Z��íb�U�PϷ�/��z��IGF��7���y���N���[�^wřg~h* =��#�w�/[�ԟ���.�P��E���$��x*O(u�獴Z_1�}(��p/�����r����^��Q��T�3��֦�����&״�O|���7\�t��	t��_���c���jujU0���*��G�z�v�m>��t�����C���N��b��J~�"I�0����$Y�6��M�����?���G�m��{ Q� ?����������$�^4��Z,�:O����R���e&;�g�����z�uo���f�\�`�T:���>W*�Z�?ph6o���c�t�3Wmݺ��3ϼ�� �� �g˖u�NL<��0@��֋�+��1���_��?wf�/fٔ�Co��l�:��l+��W�|z~�#M7���>��x�b���ܼ���=��[ Q� �q�W��j�S�!��ս�:t�|}=IF��=��Yݑ����ُM��*#s���ޞ����b�ryme��[̵4�(����韘����B�]Y����eˆK֮�a  :�g�������I�Ь��_yU�\V�W���ב�+���%�F���w��e6&W�^VM�e}�~��5l�����T�S D�R�^>>�����= ����p���n��A
W*�]�����͏�b�r����jmi��,�ݙ���d���J�t�H?��'�x�V�vtf��Y�?�H�s���_��g��W DE�C�k_��7,�q^i(�/��JgDww{��A�����<j�;ߧ��͍N��v�ry-I����$Y�V�����0�e���g���-��_���O �!Ё��{�z���S?��I��j��	��|��e�^�Lf�.��������'+�7W�œ"����;߫��33���}Gz7]�r���~�����曟 DA�C�_�jQ���%I�oW��F9yk-M�-����RU�o�E��'�`�5�57Ow�;����~��G�V�ދ�E�ݽTj�����,{�eI��h�N�a"Ё�u�1��s�4�8��$����m�|[��
��ȕ�H��T��~X���ً�Ρ�^�C������G�7:�����o��:���x3p��w���h��熾7����"fq_�H�ե��|���� ?B��\gf�#+�+���|�rh��5߹f0�#+V<��l�r��׮�ԝ���/��_��'ML<��}w��_�j��lo'_-�#�Q�h|r�\��Z,�:����#��md���#�(#=?�b���u�u�y懦 G�@����o({��T(�GB���ޯ}�ߕ�3>4���v�!�3�Ѹm����-��8���>����J�aC���JezY���{O! p�t`��z��[�8!��Cq���o�}����\^���>��m�ֽ��{���Z?�˷��W�"��hg/,Y��[��׾�u��> pTt`hl�x��+V����wV�G���a`Tӑ������'�)�^@���V�;=��K�o}�X<��e?]m6o�u�B�{����ڰ���o� �w
��zI}͚=��TK�ZR�^ݷS����n����h|z�dw~��8D����\w��N�3��k*��k�֖F�P��]��������y'Ё��zu��+��%�O�J���6���(_Qʲ�G��;g���3���O�ғ��w�^._0�Gz��p+Dh���_��t����_ �J�o˖�߸l��W�>�$#�8�h��\�tv%��t��~�,�ݙ��W��>���$��,;0��<�Ը���޳y�Ϝ{�� �@Z>�}ٲ��_��'I!�����鲾��_�<\�R�v���eG��B<��=�C���.��U�'I)�T�V����d/ԣ;�Q(4������? �7h�������ա/%�\^׋�ե0T
�pɇ�}�.��G���'�j���ݙ�|�?�~�Ѐ���H_�x��[�\�a�ڛn ���M��v���O^�T�|Q�X<��P�z(\>��vt�B\�lWgv��S�J�ݽ������B��j�q�t�L�e�ʕ�~c���n>��M �@֊{�}�v�r��\>�R*���X���R��.���E���������v���b�r����j��d�Rifq������� ����@ں��_�׷��P��z�T:o$��pɇ�5����s�
�ۦ+��j�>��G��7�t��:�����%Kv]�q�_p�-� �)��M��Y�bŷ�A�C�B�|I���\�?��v����4ٝ���~��$c�����W����ff>r0˦"�2�MW���;�_���k����F�9$Ё�3>���
�>\�M+�����΁�sh�{��w2?k�'h��i�颴X|u_I��5`]}v�㓽(1�V�V�|�_�=�` `�t`��y��7��?u~�;ŤZ����A�-����[�33q0˦#[]$F���g�t������N~�Z�5�BaY!��ї/���7^�g\��� s�o~h�U����|;f�3���s��K�$ґ���gg?6�eѵ�ɿGfg?3U��k,��	Q�f��n����?�!y�g�L�>
�����{��� �@�W�z�?}�U�ϔJ���J��uj/V��,�Jo�5��Fw%�Ƀ�Ѹqjd���|����*zݝ��v:�u�!p��3�C���y}��%{�r�]��:��� 8�:0�kCuŊ'���BaU1��8l��Y�\�WR�<���;g��js��ʷ�g��^��!�����v�֎�nab��zO� �8�������x�#IRO*�+k�vgs��G���N��xtWR�Vkk3M'���)Gl�J~^����-���6GFG��~�=�������� �%Ё�w���^�t�ΫC_I����^�Gv6�_�߾�����d��w(�������L����$_䬇n�eS����v�m��cG{؇NL���m�6|���oh ����c����4m��uJ�ҹ#izl)�2T�J����̇�0ԭ�aif��-�##F_x��`��K����N��{{O' p�t��m�t�ً=}n�#���b�|N_}��4]R(�+�����t��4��4���F����Z�|���l��Gk�ް? pDt��-]:���t�Z�T��5;ߢxY�l��j�=�n?!�9l��g�����s�Ph�+�����_ ��������;#��r��j����
qjg�����ݍ��"u�8?r�.�}�m�]��K.�Ԟ ��&Ё��t��ik}�X<�\,���,���o��;gC�X�B�]]�j*_E�� ��&Ё��y��7��=��O�O�d,�T����y��h�1�e���,Y���7^�\��� /�@�Ҳe��z�e}�z�_�vY5�:x��f���Vk[Ӥv�S~������{����E�}g˖����=yb����J�-��jW��H���Z���3Yv�vv����{.߲嚕k�~rg �%�@�Y�d_��������ÖeS�f�3��C� �|�^?�[���8 �	t���}��o�ן<!�J%��^���v��f���١����dӦkV�w�'� �$�+˖��ՙb�R�x��퇥�5�_�m��m�/�i��`�d>��=��D�}c�����ן89�$I�埲��0t��;��-S��g͡ύ����/_�n�g ^4���˧�y�{�K��G��fj�OphK��f�� ��B�U;������ ��&Ё�p���^16����
��R��r�eY+k6o�6�ҥ��y��~��ko� ^��+�����>x�JB���ji_�����F�3S��3޼� *�f������� ���ov�a��g�uI���i�B���/ �v���?=¤��0��,y����y	Do����f\+&��y#���~��h�2�9�z��q�7����so�l �	t jY��t��[�}�T:��$c������f3��\�ðX�d��~� /�@�v����5kf��荦���*��e��fZ���*<���ןr�7> 8,�������@�|�H����ݬ���L��M��P���_�=yO �t Zw�y�	cc��"�$�
��ɥ������^���8�!�p��7o����ڵ�ŕ� �A������
L�ܡ�p�U��^���s �JͱBa�����3 �	t J�_��0>���C�
��B�x���������8X�߶p�����@8�TQ:��ɟ)g���o�7�B��}v���N�Qq|����W�G����O= ��:�ŋ��"W(�*��p��۲o�9����M-�|w�ɯ ~,�D�_|�+GG�|u�\�x�kվ���4k �B-z��,{�o$����$Ё�,Y2��+���5^CC�4��͍ ���Ƣ{����ӏ ^�7�@t��\"W.�Wq�<�v��f���� ���O�� �~,�De���o.��X"��K�4}�П=�t�����N����dll�7�|��u�>{  �#	t *L_"W,����Y6�m4n�ʲN 8i�)�\��L�� �H���؁sCĒ���J'��y~��-�Y6m�xQ��&����:�����r��E!b�♕
C�z�l~i&�� ^��у����Z��?��� �@�Q��"�$�P*�^C��~��j}�uj�K������������ ��"Ё(d���;n�z{{�pJ9IjQ_�6���ݝF�s&�/���3���#	t 
�7�s���7���J����,kf����
���9����O۲�]K׮��� ��@-�}G�X�����ˇ�5����L�����)I��ry~'� ���}�	������	+����n��V��͹s��=�os� ?D�G��w��ӯ|es4D��
'e�gY#�����޳ p��jOں����g~h* �=8�FGW���J����<�W��ZwLg�A[ہ#*���j�}[��G �#Ё��^��|{�)C�z�n?�j���
 s`ll�-A�� �U7^��V{lu�T���i:QC&���l�> �H�>yf �tਪכ��������<�Ði�6�fٴ�����Tf��u�U�9��O? �6�U���E!b��ɥ0d�lo�ݾ� �X�>{U���8j�s�ګC�
�U�$Y8t���/�dY' ̵���7 �G�G͝wn���O��z�Ba�V���G���� 0���n����e���5� Ё�h|<[���b��!�v�l~q6 ̓4�/.�Wm~,  Ё��^�:;D�PXYH��h��ͅf�F�p�90�FG��m8*�m�P�V^"��'�����j��W��]�6�,��&Ё�bjj����;�n!/�^5T������,�q�0�FF&W;�p�P��Q�5�"�$����C3�=˚Vρ�&I�����O��� ��@��ju�!R��+�굱����sਪכ� Ё��Z�>!D�PxE�[�4��@���3 ��6��R��(�?O���P��������W�<!�ޗ&���$5�̻Z����BaM�u������Z����G]�Ю~�+���{�� 0�:0�*��ׇH
���n?�ʲ)��@j�v~�@��м�Q�Μ"U(;4������ �Zm�� 0��(���ۑ�疇(��I�p(Οg��N��� "Q�� ��@���h���i�P����yMl�h�2= Ģ\�]��C�T9�?2ZC�f�C���"�����51�Z���z+ D$I���{<�� 0����(�j�ur�T��j(��w:5ChX>�S�w�s�Z�W���+C����$ɂ(��i���Vρ(���N CL��jddvU�P��*�\�Mw;���Q���0(j�7_���5����Ba�Ploo�i�� 1*���`�t`ތ�&�H
C��C���*��c7^���>�\ B�7�R�!JIH�e趷�˲,)����� ��@���H�U!BI2��P�q���`d���+Ё�$ЁyS*�&B��t�����:�Gmo�W.�� CJ��X�]"4��κݧmo�W.�W�!%Ёyq�]��҃��4]2�����lgY' ĮXl. CJ��Ph��il*����N��9����x R�i�:5D(I
�7�:��:�Ҵ]q�0�:0/���+C�����Q��)Y�̺�g�o�F�6O��"Ё�#Ёy���!B������p��+##�{�� ��@�E��\"�$����v�ہ�R(�� CH��Tj-J�a�g,�}�\� ��@�E�܌r*o��A���@_)��`	t`�]��B���Z�РOpϲ��,��@)�����;����^*F8)=�z}����c��;�R'�u�@�\�يt@\-�F�����e���'M�� 0�:0�Ҵe�;�^�W�kC���o�	 CD�s�XQNpat}�@�R�3���X "�s�bwi�P�����^�gY�|7 ��J��Or��P���+���C�Ҵ>Ё�eӽ@������ր�#Ё9���E!JՁ���t��@�*��%`�t`�
�(=I�����t�9зҴ����#Ё9W,v�B�F|���t�o�~vDy<
`.	t`�%Iw$D(M���[i��:��R�Ri��w��e� 0d:0�$+�%I%2[܁~�$�~�0w:0�z��kMq�W�ChXA�V�g�@�N�o��A��qz��|��;Ё�U(��(�4���Qnq����i�[I�}*0|��s.�3���y2�+�!�:з�A��@�A7�@O�4>[܁�%Ёa$Ё9�{�]�g٠���ZVЁ��e�������̹}�ϟw{�m���+�� s�0��O>�[�]���l�?I�[:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@�  @:   D@� ����n%˲�h~i�t+�� x �t:Ya׮沣�5��|v��ʳ��'� ^@�^�n6�����^ `�	t �c|��������c �@ �	�.��k��F�; `�t �� IB�bEe׎3+��P 0: �aH�Н��E��D�
 �0� p��Ť�bE幝;�?<�ׯ0x:� ˲�LOw���H�(��|���;ɗ-+�>�ׯ0x:��j4��]�K��P
0�j�t�^�L��?��k ��0�ff�#;w6[pp##�����G���5 �4�0@:�N:5ըu:-�x�J:�OV?�_��� 8�:��h6ۥ��F-�(��F���gG��p� G�@�sY�%SS��v��9C�X�+ʻ�k�B\���"��X��.�[ڃ���^w&&*��������5 ��Ч���f�mK-C�q^,�Q��w�+���*: /�@�3�v����gY�I��
u���B�zQ�>�lc�8��� }dv�Y��m�Ͱ��=W����<ο3$� ^����n:99[�v3�s�l��򮑑�"�e!y��r�8:@�\��0[����V+̄�q�쳍e�f� �� �r}�n��Ҟ���t��s�5���v� ��!ק1�-*�[��8"�kWc��L�� �(�ק1�za�Ѣҁ�={Z�SS��  G�@���� �z==�xq����{[�l/ 0:@\�!T����e��!R����h/ 0G:�Q��48�RIg�/���������k/ 0�:�Q����	��1���11Qy.IB"45թ���\ `�	t�y��4��RҌ9�gf:#�v�s �@�G�O��Q,�V�i�!B���ʳ�6��`�t�y��4��(�LL�<W($��F��g�N������V���[-ɒ�o�`v؆d�ea	��H�,����xϙw�L�03gNf81�I�Ֆm6�%��a��W���ޫ�k�����V�mY��ꮪ���~Nn��2������S33M� �U: tǧ�en���ض዆</�U�G��5 �* :��Ӏ�Z��T��DC�Z��ͩ0NV  t� R�Գl<F�eKj�u͖h(�rS�yp �~ @��!Sځ5�q��Xѐ��S�/�� �  t�ؘ���Zu�P�13Ӝ���M =E� ����CCvE4���f�^ ��#� @��K##βhjv�9�h� @:  �\�,��:%���|k�^� �&t  ���8�LN�����o�R	� �Ft  ��2����h�X��eH  ��  6�뚍-[�y�T��J%D  ��  6E*e6�nugC"�P��EL  ��  6̶��9�k� 3?ߚ  4F� ��,�mKϘ����z=H�ζ&  ��  ���Ql���X�����=�  �9  �Ðpjʝu��Z�33��Eb
  	@� ��8w]�%�О�nN� �$!� �zE[����i�)
��Rq�b	  	B� �u��L�g�V]4G�y�`c*�� $?�  �qsr9�&Rq����)�G  H   ���84dWDCQ$��Ls2��  �P:  8�8�K##βhh5Λ�0-  $�  �P>o��Ɯ%���\s��3 @��  ਲY�:1�,���8��  �t  pD�Y��tDS���H� �>A� ��I���Ԕ;g���Eoxy�  ��  ö��u�;�k��J^�T�G �>C� �G�q�mۖ�5M	EC岟+�1 ��  �-��`jʝ�,#�jAfa�  ��  �0$ܺ՝q���Azv�5?5 �>E� 0�V�<�2=�P���s �  � l����fK4�y�=3��Eb
  }�@ `pE[����i�)���:x��5�   � ��w�Y�.
�Ț�nN� �AB� 0�FG��B�����(7�8����  �@ `��K��NY4Eb�8��(%   �R(�ˣ�NI4��|f�9�j��  0�t  D.gV�ǝ�hjv�9�h� `@�  �LƬMN������x�f �F� ��\�ll��΋���j5�  �@ ���Rfs�Vw�0$-.z#�?$  �@ �_ٶ�t��R�+,/��  �t  ��e��m[z�4%��~�X��  <�@ ���Ql���X����� ���M  x �>b�8w���Azn�E� p:  �#1|ߏ�аLӐ���}����k4Bwf��%~j  x ��e2�R����i�ѡh�2���,k5�W~�\��ff��9  O�@ �d2aɶ�ֱ��0�0\�d����W��*�x˲N8�=/�U�G���<  �( ��s�`9���f��(����m��]��;���Wo;���Ț�nN��X  �� @��nXN��z���8���j?���SW�]=���c������ �~ ���L  *�
+�U��{��)7�Z��  p\t  �q�U�PI��H�  �� @��v�H�òh�^7���L	  X �����vlM���p�  �u#� H�[�l�$����!�7�  N� @XV�e2��y�a|��  8a:  �3���f�b�45�f��̬  �!� ИaD�J�GZ�y�edZ-3/  `�t  ��*��HEC�g��MsH  �� � �P��¢iF�h��M�^7�C  �&!� Ќ�s5rnY�/�}#U��8�� �L:  zQq�dۑ'��ܩ���: `��  h$���8o������u� �N!� Є�ˎ5DCahX��9*b�  :�@ @��S��.�"�$� �< �s���J�5�P�Y���q�[  :�@ ��l;���aE4Eb4�H�/  ��� �Gl;jd2�hJ��ǹ#  �+t  z�4�V�%��J��)  ]C� �eq�{�s�T�n��
  �* �.2�ȏ�h��k����  ��#� �È����{��  �:  ]��\�Gz(j6͜�9  =C� �qz�y�edZ-3/  ��t  :(��q^4�(y��n6�!  =G� �!*��n���!�7�z�6   � �l6*�v������M�  ��  t@:�q6ECq�;��9�9y �Ft  6Y*�'j������u猝 � �M�J�׍j��04�Z�1L  �!� �$��\7�����0�s  �F� �	'���aY4Eb�8�#�  �- �������hH�y�n�����|  4�k � �0�؄k �f�Rg����n�q�;�����T�m[�  �� �(���f�o�L��eE^&�{��)A���+�R-�N��\�� зt �$j���|3��f�| �f�g2A�0$���p�)�
�F�Ѳ=/��y�c4 �� ���<F��aDA6j獆5��FZ�w��j4=�q�l6�h: � 6@M=m�<+CF�F��y��f�a�=���Z�޴Ջ��|�3MC��  �G��	bJ������\.,�f��#�yfN0��5����;���F ��!��0�}�8W#�i9���22�g�E��Y^�3� �� �������|ɶ#O4�yf��4�KMyW#�B�)� �`: '���L&,�q����6�`�Y=j�{��f�w H( ����*�-��q�`9��h(��tj5c��%#�f��H���^:�h�W ��t 8֛�T*(�RQ]4�]����A���Ն��˹�K�!��(Xo>�R���QM4JZ�9���h��bc]: $� G�z���JE5�����S�Tq.b0�Ǵ�.}h(Ӳ,�H �� p�j�\0�l;j�nP�8�Vͱ���O��u�j�8�K �� �q>�,+l��ECQ$F�n��8j6�:/=I���~��w����~��?�z�A��!l7�L3l���EC*�k5s$G�P�ǅadd��lZ'�t��������Mo��  � �qn��FPj�mG	��C��.r�P�i��i�4Bӌ�������כ��3	;���o��q�߾󝯾��k>��>G�h��S�m�-q�y�Q&h���o娷@���]�l'.��û���ϧ=�\.W7�ƾ��w�{�)��M� }�@0�"�Q0��M��/2���T���{n��-��{�[���E�Hꦔ80��q�j�������m������ş�O� �S:����R�;##�9 �����Hߵ랳���|�o��W	 �!�@Qq^.ם H%zC8 �LI�t�P���W����5�}@ ��� �j��Q��s x��HWk���I�R�15�����O�z�?�S�>B�*Η�� ����S���W�>�>4T�j�~����2Φq �	�����W��� p,������[�,�}���?}� @� ���r��R7� 8.jw�J���~N��]?}���_�WW_���* �t }M�`�M ��:'�0�(�s��BnY�LM�����{n����{ �@зT��L ��F�e��ٔ����׭r��w�O� �@Зj��M�����M�4�(�v�Զm����_���/�� @�� �N��Y�R  ��Zm8�eD�c����O��{׻^��o��- 	�,���6�S7� �T�r�QǯY���l;0FF~���o�G8z@R� ��:�\�@
 `�EQ�{ljx8�T��u41���}��w�O�. �@:����:�PϻF �A�#]�3�w��Ʌ�_�'W\}���' �0:���vl�s �<ut�ڈSם�'���o������k���) � :��c�v �.�wv_J�J?�z��"�!�$��a�v �>�!��X�����������/~�o�� @BpS �Ԧp�J�M� �G��"���h�qcx���ȵQ�� �$��1dS8 �����^�ϧ=�жm��]/�����W $ � ������� ��� ��Ɨ��ѷn��+��~��u��xX @s:��Q#6�S�@�jӶm+Tǉf�����x��ӳ 4G�H�(��\n� ��ܨ\�k�}۶��񶷽���^��� h�@�(�j�u� ����Mz���8������ ��t ��n�8� ����t];������{�;��/���O�/ M� ��� �?]�^3M����5~J��� ԴI�����l�Fó�iG�]�'&�w������_* �!���͞�6) �D�՚�:zM�]������o���=�ڭ� nxhO�# �Ĉ��PS݇�2�Mu]v~����O_# �nzhMM�T#� H��Mu9��f&'�~���RF��@��0��z���) H�J�錎�M���Ȳ���uk��U �����8�� �K}�wø�_& ����@��1z I��qj������W_��� 4��/ -U�M�<�>�6�S3�r9W���CC?����@��vV7 @_P3��4w�2�E���˼���?o|�'�Z @: ��jLm�~���
O4�������@�n�hE��s� ��V�W�f�miu���ԃ�o{��_x��� @�� ���9 �/��{>�W�[�S(<����� =ƍ0 m0z �����L&���7'��m�s�^{KU ��t �`� �_�޲���Vk�3��i۳�Z ����F�`0�Q�l��u;}x��? �1��u��G 0 Ԏ�o�2���W���o�� =�1������s :���f$�����O	t =C��9���  J����F���c'w =E��9u6�  ��,N�@�Yo�%o~ӛ>y� @� zJ���ah `����jy���Z����|}�@��	@O�u� Hͦo��cc�� �@Ϩc�8Z ������u��o�_��M��� ]F��6� đnf2)�֢��/�t ]G���c� ��(T�@��& �:��P�9 @-u
�а,S�i�CCe��o�K����>- �E:��P	  ��3!�M��	Èo���?%�t��'�� X�fU��D'��̓ ��@�uLo �����ad贛���l����u�����( �%:��k�= <�n��;N`4��%~�F�.!�t�ڱW  XC���]�� ]D��*�S/�� �S�ܣ(���GD6;�S ��t ]��p ��Q��8v(�Y̼�W��\s}S �t ]��S/  ��ya�M��R�E��>~�7 ]@��*�	t ��xܚm/�Jt ]B�蚕ctX 82�[K���	 t	��k|�8 <� �@�5
��� @�� ���� �c�m��P�y��v箽��� @�� ���� �cQ��E#���T��O�N ��t ]�ζe�9 �X�@���Y~�� ��@���V#"  =�s�Fq��)�+ �:��`�8 ��RŉFR�� @� �B�)�  =����Ϗ׭� ��@��m� ��ʲ(Kt��չg�|����' �Kͺ2}�u=����']sͭw t��+�� p�ԋ��>}�E՗�:��"�t�� ��P/���ݼX ��t ��9 `����Q�. �a:��c �^���0�Ƙ @�� :.$� �E��Ķ�� @�� :. �.���kY�� @�� :." �.����R F�  @;����#�t\|��: `]t��aY,��y:���m ��2��@�q:   ��ۋ��E��<@ǅah��  �t �@�   �`Y� @�� �!�e�a����C��
 ���3L3�e E�^A�:�n �t�ډw��۶�	���Ʉ˂�C����� �t����M���m @wGt@:�n�& �.:�AD��C��ZL �Z��C�@7���t �( `���`� :��, �	�g��C��8�v� �O�c� �t !� X� �����t �@���&�b�" `=|�w@��>� X��
tF�t���<Ϗ=%  �8�)b �@�q�0M �.Aj茠�@ǱI `=|�{T ��o~ :�i� ��C�D3���@Wx�8�#�  p�f��ft �@��
ϋR�c� �c�{T �o~ �����lV� ���M_�{TF�t�V�� ����- pl��kU�:�n!�tE�峓; ���@,�X�"��#�t���=�4M	 ��h�h�@�-:��QŹ��  �"�Y��z(���@�4�a�� 8�z���)���7@ ]�t9CC �httF�t�V� ����ˊ�L{)�  p�VK�H���:�n"�t����<I�R�  S�{�hF�n
 �B��F#pS)�@ <N��A��F��Z��b: �H�R(�q��t ]�h�L֡ �����t����N���i�.  R�yi����猦�@�U*�8�] ��J���� ��@�u�J�w�� hS'|x��U� z�@�uLs �U�z��J��@O0� �J����t =���OL� l�f���v�t �@��	5ͽш2Ls��V������1k ��@�3�r+�4w l�r#��Q�:���T���x�2�( ����Ì�ڕ/���
���*?74d- `�,/7��F�����J��;4T �`�}�k��%�a�@/� zJMmd�8 <���� z�@�sj�c:�&�`�,/׵���� z�@�s�j����cۑ' ��W��� ��a�:��{�Y�: -,-5�nQ  }�T�kw���:�^#�h�\�;##�m�� �o�ja����[�}��&C� :�@��r�ˏ�:K �[KKu�VS�hz�Eڽ� �� �Q*�R��#�iF�  �N�ft=?���a��w �G�Іڀgy��qJ �;KK-�V;���
���<�V��j����iQ( ���lF�F����r<#�o�s	@�� ��Fї�ZC�E����Xϋ���9܊ H� :�@����j�P�\t ���s]GϏoz�
t��Q t�@K���-�E $Z���X�r���=_��Ec G��R�ڰ�M7�FC  ����|?�r��=W|�i
 t�@[����9 *�*ki���F��1k�e�#�hK����-�rfU  �S,6���:Z��.ˮ t�@k�l6;\��5 H�VK�r��;z�AzZ ��t Z��XXhOL�E $��|� �:�@I�B ��t �S#0�B��  !J%oH-S�87���Yg���
 t� �檅;
���=  my�8�n��w���4�� �0@"x�o����QgI  ښ���1܉MmW��f���zOM ��t ���TM���D�E Z^
�FK˩�ʉ��+�F�% �:�D���mߞ�7�sx ��ھ�XɈ�N4���5 ]A�H�V�3��<���ft�ڮ6�;����� �@⨩���p6�1X (��~�ھ*
� �@"�Ζ�;w7M3
 �3�z�Q/���������V�?& �:�D
�Pff��۶e� �A ��\%/���y��	����o
 t� ��t�R)5<<l� �u���� 76<�A*�7:z^��UD� �@�-.V܉��=����� �-��?\�576<�A�nU�5�� @�� -����r٬�j�� �q�z�U/���6:�}���A��!�$���Ţ����s��R�h|�% ��Q���,k��\��otj�Ej���� ��@�X�3&�ܙ��a���a�YX����� �b��TFt=�\Qa�Y���Hk߾��H �Kt �52�tu#����f*��� ����P  �jv�>�y����)��J�6uP�� �B�H$�J��Г��V˴��K�j��JaX�w� fq�5R�77��Zm���U��� ]D�H�����������.ɗ����N��-/�R���m��v%����! �E:��1KFF����L���
/�*�OT�� ���V���B9#���8W�ձ���7�B ��t �S(<Il�p�9���X6�}AT�~�*t X�f3J��.�Ds*�7sj�R�o}P�^�n"�$���E���EQdx��\>���R���  �[�%����C�9��\]����� @�� %�=E\w긇I��k��YC�|U*_j
 ���Y�?\��85e�ם�
;?�? t� QFF.^��FE��Gz�T��kK  G˴���Gt�s�q��'_���� ��@��Ըd�������}�0�:���Z�D: ��==]��@�ΕN�;_�h����w ��@�j����ݘ�y�m?-���T�����`���������y�֝+jz{�1� =@�H��J�pކߏI���H�J hS#�.'b�S��W�J'_��	 � � ���&��lʍ��t���u��2����8Wl�������az;�^!�h�0�8�/����"}y���� �ڭ}z�<B��+
Ñk z�@�����㛲ܦ�<A`�H/2u�0�߮ 6���ڭ=IqީM�V�J'�����!�hΐ���:��Ez�P�6L� @��,%�(5��;��U�����w z�@�5���ю�����j:���e�� @�ף���r>)q����j4����^��"� ���<�$~R�m�$2�c�'��H�5m�� ���rPXX(g$!:�c�Z������%om ����VF>N|�x������lݪ"����r����Y�q,�I�W�8��<-	��ӛ­
CC�-o �1@ǭ�~��锕���H�t�/�x�W*�T6�6\�i	 $\���XXh���uG��q�,-�Xz�k?�e�#�t����}��~����25���Gz��p|?0s�4�$V��Lu��hu~�&�f�+�ک��|O ��t ]��^.�$��l�֭����Ho�<+�tuV:ǰH�3���塤����q�h��SN9�M" �5@W���*�7beM�?�פ����O��{�TͰ�;�$�V���\9����Wu����g��%/y+������V�n<�%?|�l���8�S��[��=�M{�K��R�^\���0��s�w�fs�n M� �n�"�^�?��ɶm��,+��:�.=B3�uY�@;a(��l}�^o&j��ҋ8W����W�|� �&t =�y���<��-�}��D�3��f��^���g�i���q ����(=;[)$m��ҫ8C;j4v� ���g6+�[��8�đ���u�:~��Q*U2�|��y� z-i盯ի8W�����W�� �� zj�"��+��CnOw�dvt�nO���)�)� zA�6;[M�v��q���j;� �������8>�-q�D�lyA44t~W��Ԕw��Քwvy�5�F���.��K��^ƹ��p��W^y� �!�hc3�I�"_ff>���G�㿣n ;~��bc�w �{4���ᥥjJ��qE����� �nt ZٌH�o��X�S<oI��^���W�]�=/�r9��|&sX��Z-qgg+C��'n#8euIS�-,�zpϞ�>+ ������lN��5����,۶�,��|Wnh=�3���,�� 6�5/���b�����W��A`G��{D� �Q�S��� �����F�!y��e�֗E��I]uR�魖o�r�&Ǳ8Q�g�33�Ď�+�Ĺ2?�O^��[�, �)=�[�X��~�h����~����v46�̮����o���M�^�0j�������^k63A&s� 4F�К��S�/j4}#�(���;ڛ�m��ҭu�
�� ֣Ւ��\��jy�5W��o�XX���{��� ��t �S7x*�7zV�R.�$�����[/�R�Ѯ����n�ɤ87���X�bs�\�;�p��y�<�ܵ�i,� :#�$��F5�����͙��tu^z�pnWG����l���\�s� �aaa��I��k���#YZzʻ���ߺ�Wy��t ��雱�{6ez�SR��ML����ݵ���c7*�Z�q;�u��0ut��|��lz�7� �6�[�X�Uܿ���( � �}�cP7��5*A�j�u����ј��[_�Rc]�QG��J^&�I��� #��t���Z⧳+:m����Q�t���
 $� �\wL&'_,���(���7����i�������D##u}^f�ް��w����F�i �!�iz	���0�� �/���֛�57w�׮��ß H@bY�kl���hq񛲰���N�'*���F�_�Z�u45�b��\WC}u�{|��c�u��:�+RC2P� �JN��	rq�g}?�k����|���d}��g�"�$ �:�D�o���gK:�=:x����Z��r�����E���]�������X������@�5�Q:�|?�3_��|�L��%�ʅW���l Yt }!�;�ص�8��A��7����*?|����D[�� �	Mw�T�O_Z�2��Rǲšn��\X`����ZX�j��~��7@���k�Ξ�ý{o�� @�� �F*5G��hz�������J��8����ߏ���z2L�l��ǲ�RN�ͦ[������)�J��w�Y:Oi_U���\����� @��� ��0lc۶K.wZ4;�y	��-Q���<�	zJ41�����+��g�W�P���a����Uah���oٿ��* 	�w?@ @:��dN������o��-/�H��_���󢡡�{v���L}����/.���j�/㮝0�}���y?ۿ���S  ���	 (�3d���g���w⛶/Kzjm���g���hr����?ܳP_���B=�N�L�`D�*3���axV~n���(J?J�U��d��Ӟ�4�� ��@���.K:�#:x�S�y�~���/�V�OFG���=+�3�^�z�q�0�I�,��ث ��i:Eg����m��c��H�X,�)�BE����}'�V/��g?��u�K�w^ ؀Lf�q�)�Gss��Q�(un�����X��LN�^��������=�Җe���9����1�L�5~~A����,���w�0���/��d�=�����S��ۯ<$���o}l�ޛ>+ �p:��a��15���͞��~���F5������B��&r�]�i�A�>G�0'��$e����_�������);��+ƩN�e��_�CC����}��f��鶤�����?�{?�j�>���� �A���F6{J47�%)��ql�g-�r��T~ٞ�>:�L1M���E�E[SQ�m<�}�E��5��o�a�M�cR#ȧf㼬al��n=�gם4v����|�}TcR$q�\�Ն���SK� ��@0�,�5�n}��MOnSF�V����?���߉����kे�P�VK��3d���������փ��_�X?�
j��FZ��	+��ʛ�Y)��	תi��/--m�����_�����Qs%�hq�^�U� ���� �$���^�>?������M�����LOR��m21����O_�Q�q�Tj��N���_I�~w������&o�}�0�8����a����'~�j��g���G�ӟڔ%5�-�����.��e�}� }�@0����-[�/��Y���Vk~S�o�q��>=�?+WH�j�a|��g�I.w�����Z����
0gg|���a��
C���\��Ν�"��]���� I���������
 � �dv���?ZX�S�ٞ��q�T*?k�64��hl�9=�Hn���w���c�%��c���e|��,WG���a�geE�JG�p�(�§�m獓Nz͡���^}m���*̓r��єJ[�Ap��"_ �7: �a�11��dx����l��O6��FQ�T�@��*##F��ϊo�3��%��꾯���,�ԩq���x�M;�}�(@r��>=-rFFd�E���գ�\wk4;�������J������s�� }�@�#p���}�K�Z}J|3��M���F��o�w��(�.�o�Ӣ5^č�s$�9/��v�7���[G�0\ò�p�LmwD,m^+�1\w�}[����?�_�\	'*���q��H �O� �r�Sڛ�--}O���ksSޯz?��_����đ��C����9��:?���ď����p���'�g�/�,�GʣhgZd��F�#MWi�RƎ{�8б���e:����y������ �� �`�1:z����D�����g���7ڡ>4�Qg��v^t�2�>־���AԈ�v0��ټ�=��#��Ȯ��N7�&앓
��D��=R,~�cq���ُdz��o���W �9 ����~�I,�����ܗ���7�}���*�������#�3,�Z�	>%jͺm�{$A�b��8��-�=�:��3W\wg�;�k��d��0���凄a3R_��8�N��O���ZX8}zϞ~� �  �`�2��Ʈ]��Z�M�_��tv�޷Z����S#�q��s��Dg*�[������5����{,���`"��yӛr�<�m�Ɨ���k*��
�;���:�\�(W���|M7~��ȟ��\]�3��Q���Ү]�:]�N�A@��r�������gr�S�l��hy�'2?������-��n_�̎���l��D܀�q9���T���ǯ�Z�C~.��3��M:���4s��Ͷ�s}��Q�n�2���YF�j-F�65jީ���[g�X��[j�Կ?��Ͼ�)9 ���J��4ﾑ�������~�ڙ9*��>?}�6�[U�?_/��E����Y���H�L�W�V�ݶ��ڶ��h�3�����}q�OQ��m�G��e�jF���r�sG�Q�UQ�V�U{L�v�t�c��0W���V��ԧ_q�u�s� $��㮼���7�|Ź���^(��u��&������<5ZXP��}�G��T������;dh�8�/��$Q��_��gL]Ӽ J���0�(����8������*�:q��ş�*�'������6 \�䌒�
�V����������MQA�:������ࡇ.|��^w�� ��+��y߃7ݴ�9���������cYYc˖ߕ���D��w�g�o���Z�Z,�������GF�&��)�M��̈���PW�0�ϻ��f3��y�0f[�7��� +D{��v!���A9~Nďc�߹)����'w�fs���[���M�:_kP�\��tX.?g��^w� �oo��g��|����R���?�����jx��ϕ�ы:�j�z�����F�ը�:�Ͷ��� 7��<C�I���W�4���G{�P��5}_E�\�Q������R!>ҾLs"~�����W�<ٯ���ru�b��i4��5Ha���MO?�͗]v�G ������#���z[:]��HWVC}d�鑚�ډPW<oI�"��_�\��8ԟ*���kTWF���_Ċ+e*���v��R*�U���p/������]}1d#�ΰ�B|ǟ[�q8�k�=2E�#1��<�OVF�$��O::Z�Z�+*�gg��_.��#� `:���#�����WLL|��3���tŶ��F�/�T��M�:q�RR���}��Ņ��q��/�Ը��G�]���?���I�8h"۶"�5CèaX
D��Ȓ�y�H�m��R$�J�0n����W�F�е�Qdɣg���_��ըR�[����<N�h1������˽{?�? ��'���S*�''����0��ʲ�q�����?;Z^�'Z\���juf�b�/K�����Noo�����c�~��݉Ʃi���S�nY�8����d5���o� �yO��Z�">J}9ov|���?��+�w�ǿ���g�!n��8��ǌ��Jڮ�'"��Z�e{��V�u{)I�®�Gsh��?�q��  ���o��K'&��f׭ԐQJ����U���=��V����yj����y�j�{�p��rg�1��Aqh�]�$h�=?d��Q��q���Nݎ�Fh�8�[�G�f�Fߣ��a=~_�8���q�ף�����7'�҆eL�U����~��~�����Z�0��j�H�ϣ�O$��Hg�F���{:>�}��h� ����n87��o޻�CLk�Ct =�o߭��w��ǿ~[&S������3�W�1-���jGB�F��y�˩�S���'��~Z
��#AmPw(\��R���x*�V�^�������㞏��y���Rq�-Q�M�^{�~e�>�����Z�������`+g޻���oS�C���<�1n�~����Tl�������7+�D=�������>ծ��*�Ո� �<7��}����л ������&�����ߛ����ܲ#*��*۷�4�q�)�-��?��:�U*W�����c������AY?Q*�U������!jBH����P^�#����G�{�F�7��Q>��ˏD����s߸���s 8�@W^y�7�x�s��ί��Ł�C�u���俏#������NW�(o�|w�R#���)q��՞oY�J���~ԺruA��� �/?�V+��>����?t�  �@��}�|���sa}绅�|��dv�Ԇ^j���Z�QG<�J��診�F��oJ:��=������ ���J���}ҋ����x�ڰW,>�%�]v�� 8"�V����{�?O�o�;6����M�69�<QG�ukT]Qk����ۗ�����l��8�O�L�dYY�����6A��~G��ԙ�ҋ��-?�ju����g]~��
 �t ڹ���o�s��z���w16���G�U/���1gRw�畤T�^�R��Ԗ�txue2;�1b���%�"U{��
�n�~$��?�Rig�X<�IW^yˌ  ��@K/z���n{׍7����o����z�TjDl�~�Ȭ#��Ijt�ٜn_�����ը����]��7!�f���#�9T��@�A?"�x�̜�P�z�iW]�� ��@��ھ}_���[���[�|����duZ��z�Z�v�V�bYYI�Oj_�̎�q#�8n+A�`|�[|=$�ּ�b��Z�ľF�|{��~��7 p|t �۽�3/�馗�cr�Ϋ��p�8<փ �����n٫��)�(7ꮻ-J����,+��'$�8�gE�#WW��@�e�Q�~ah���şڻ�_& �u!�$�޽�M7�櫣�w}8�Yfg���BM�WVG�{�+C�����}��J�=�q���ś�M��1�9�yq��/�D�������.����]X�V+��>�_v�G��  ֍@�{�~���y��׾��JAp�֎ ��+���q�Z^�q�-j
|*5�\[�G���K�'����|{W�Vk���y/7t;��(g]���VǚKK��e���1j p�t �r���vo��{GG��۸�^'=c}�E]����W?>�VCg(J�&��ͭ<N�����߿Ԇ�j�6�[��������ڿV��+��o���ӧ��w�啷.
 ��� ��Ko��;�|��sz���ED�	Z'��`�E����U��r��U�G�3?����<���:�ϋM����o����X�j��a���E�����W}�Y"w
 `ct �u饟~��7���'�|�u۷?�2FS7���V�]���ǋ��>��-u^��w�V���8�w���s�ߗϗè��}�Ő�ǵ�u��~,L]� pù�g�}Ϟ��V  ��@�h{��z��߿����?��3��s�q��7�ڨQ�ƺ����(�Y�~$�a�H�>?���n����ee�Gęf�������:�0l�G����v5~��wI_y��w�W�Ö��g�z�����E���[?+ �MC�H��/��7��ڱZ�?:��]g�rg&:�tt��֫���t���E� =���Ê�u�}\�i�=�����N�z%]��l?>���߯�ȹ��㉢�Ʊ��G�o��_��M�zb%�ըv`��o�����V�\�s����#䌒w�z}nq���K��]uխ� �T:��p�U�Qr�-����:���y˖���]��#��ў�`"jm�iV��6�	��	�T4?�Gw���k �:���{����}��ӏ�_��i�]�w��޻�h���)��k��P�N4���������i t���\q�G�Eo��G���������'sW�e���M�v�A�C��s~s�i�{�%���& ��"��%�x��k�̛nz�_�|��ꤓ�c�f���9|�j��m�4u����ʄ�xǥ����|U  �G��k{�~���r��_���ϙ�dvP X�ã���am|32����R�r���w�[ �@�۽����n�q���Κ�bj�����h#��{r0"�|��D��S���|�E"� @w� ƾ}�]u���=3�寜}��#�;E=$�����s<����x�)�w�J��^v�e�C  =A�(W]u�ㇱ[n�}�����ɋ㶰��:�4�U���6�đ)�׾�籣�� @�� ��ݟx�{�{�SFG���s�=k2��I}����#E�ڷ�<���q�G��������\¨9 �@0������⇩�oο�S~�o۶g���P*b�qzx�kD~���H皷Eơ_�8��
��.�̥�~��
 @:���g�ǯ8p�򿞟��g�y��L��t<���K#�Թ����g�d�ޛ�#  �� �����2~������SO��۵��)�.P` �F�:�-,\�7�_~��+r�  �C���}�mo��׾����~�����OL\$�a� +�hi�I?n�����ߺ,  m� p���z�?����==��O�~��c��D:��)OYX^>��W\�
 @{: ť�����a�����c�����/tm{�P��F��/-=����kD�- �d ������������ٟ��g�o��o�^��
C��<gBP�G��Q�J��^��5K!AP
����3�ܶ���9����6�x)*xk��V���*Z_���઼_	y�d����!	��>��~k��7���f�,�?�w���ם�$irrvc˖g}r��W�Z�qv�V#����cﯾ�s���ί�p�	��pቡ�.� 0��z�w<��1�^p�'n �$��V���]qz�UW����x���?��y���i�����~�+��� @K� `ժ+�.NG\v���_���zg�>R���֭G�������}�'�!|= ��:�p��W0N���~�1���|��gwu-��A32�`|���>���=;O���0�:�?�󁋮��w\כ�.}fW�8_��ftt���m���ŋ���Oߞ @�� �$�qz[���W��˖M�~�Q�������۽{�Ķm����%ǽy�Ja��:�4�
�����-��s��>�l��K�
u`�<2��<S�t�p��Xq�d�ޱy���u�~�c©Bx<##���_�{��3��x�Ct��l��oj>��я~�˗�8ꨧ���Z ԁ�ٵk����v���ҕ��3	t�Cd���s�㪫��ޥK���^�3g���\�w�{ǎg|�3���S�� �C	t��jյ�V���喇nZ����=='�︩���(��~ʽ##���Yg}���qi+W�u ��	t�42�$���K­��
K�~7|?��!��������������w�Z��/��  ?�_� 	�����9�{&�G�(��X8�ȧ�bq~ Z��Ȃ��۟�,;�g�� <
���<�
?��3�a������?��(̛wL ZK�Q[�.۶{��8�����r �@H����p�-KÏ~�+}��Ó�</>!�s���ў��[O����Q�:眫�·�;��  �G�$�����w>+�FX��|��8��,+ y^۷�u׮'t���3ϼv2 �~� -��m;~���aɒ��󛏿o��سg�Ķm'�\(,?�mo���� �@	t�466/�s�s��91��	~',^��P,�������ؾ�����sŪU���-`�t��k��{�}��z{o�{X���!�<a�er�v�\�}Ϟ�_��>�W������<3 ��� m��(�m�N�;�w,��� ��a��;�����b�/9�[�?|�[?��!�{ ��E�����Y�ᇟ�w�����6�����< �Jv�Z<�k��GG�{�;���� �P� mnllAx��s��s��`���E��Y��:�y3ʗ��޽��y~ğ�\y�u!|? ��&�:���8��n}^����1Կ,�%��c�O�yޕo�~��ݻ��j�pD�ʕ���N9 3M�t���ly����5�����;����G���z���[��YvC���r���' @B: ab�+l����㮻1�����{k�y�QxZ�ԣ룻w/�q���ŋ���X�=!|# @�: ?'�
?;����_��Gc�����aX���0k֎ ��;�c��-�v-���X�'��|�G�h��4>>'l��zZ���C�����ϟ{��C��'�Li4f�;v�ctt�d����q��׆pG �V$��/##K��|��G�����̹#,X��;b���:Ϟ=s㟿�a׮e{
���>u�ŧ�r�?t ���k>?2r���|3|3���(̝{g��;COϽq�=~����,�⟭��Ν�����Ʊ<�a?��]�r��  mD�0m���{�{G�������1��
�������y�,�Y�_099'��ud���0:z��0��� �St ���yq<=��������J�}�̓����ŭ/�={��<4��kL�w�Fc���G�}d}t����w�1 �s	t �sι��q��O����s�o�i�]]�����vbw��K��yx��ٻ��S�oeͧ*FG{c�/��{���cc ��: 3�7~��q�|j��g>s޲��zvW��W
�O�={��ٳ�ϝ5kWW�	��c|/�{W|Ϟ�c�G󅂋B�w ��	t ����o�;N>5~��N;����My����'vw�8��k{o�ٳf������]1�{�X�����aa|��x�$��.�H �@��}�u��#S��\���<^�h��<�w=��{dy���q�[,�=g�h�qt~�;ݣ���{a��h�aS�E{�8�q 8x: m�S>�+N35է?�����1��,��ƞZ(�>�X;�P�3?��vu��*G�f��S(&
�zL\�FcV��1���������9&&z�M3ʛ_�(: �$�@�y���-N�q����o|���n+��]O˲Ʊ��c˳l��<�X�e�����Y�&fOL4fŹ{r�1��{�899�������'�
�f͚�٭��k͹�k2k4��_�b�h~mt����F��������u6Y(�l2ϋy�=29�5Z(����MN��32r�i�����5�ǻ���K� �� ��1�tҵ#q�yj$iÆGŚ?���y Z�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@ ZN�� �� ��,�W����JeW �6!���T(N��� �	� ��F��� �h# hIY���� h hUϭ�j/-��_ �: в�</�I��: в�,{��������� ��	t hqy�P*�腍y��<�z ��	t hq1��g͚:U�������c Z�@��`��=������y~���f͚{ �(� -����ɳ(t���/����P��y��V%���N�j���rQ�`1�_����� �	t hy�?��}ʆ��q6: �H�@�q~G��:\܇�<�?q饗��=�y�� Z�@����8^hF�����O�rpppw �!���(�n�{7�#����������~ � ���8�9��N�����7o�fw Z�@�60>>~swww�����j����  �� �֭[��Z�ޙe���ω{�'1��-���; @�: �����/���}�z��R�tm �D	t hY�}>�G���h4>^��f��� H�@��qC�8
�_Ҍ�<ϯ�V��J�rU ��t h�r��Z��oq����������zV*�� �� m$���b�
��0���Gb��@J: �������c���j�Z�T*� H�@�6c�1:��Ł������k����r� `�	t h3y�D�OY��1җ�J�u�2 0C: ��y��}|dddC�͞�����K�� 0: ��.�`g�Z�Tp&��z{o�q���W�^�' �!&����Z��838}�i||�s1�O���= �!$���Y���Z����<-��^166�š������� �� Ц&''��P(�a�Eh쇸e�+��>����; � m������j���|u�@](��V���\._ � � �Ʋ,�� П��8�6F�;b�, �A$���Ũ�1����5+�����*��{ $ �����{���N��y�2�9��Z�vloo�y�x �i&��ͭ]�������(�D��}��c6n��{�a`�	t � Y��o�������������O]�v�] ��@�P*�F��j%.�L�_����r���V*�� � :D�O�j����7�Ó�,�r��7���/ x�: t���<���O
L�Eq?��Z��l��  O�@�R.���j���u�i�e��韨���J�� �@�#�oc�_���"Fz1F�_�}=.���  @�@*�����<60����j�Ν;�=88� �: t�/���z���F��/�G��&����������> `	t �P�R���j���L���H/�H?C���: t�J���V��(�<�����7o>���� �8: t�<�� ˲�����v��1w�ƍo^�z��  �A�@��T*�j�ڛc�5��a��v�����1��"�x, h���j��Ƹ�>�Y�������k��3� �* ثR�|1F�fY������������c���6 �@ ~&F��c�?+������zFoo�X����< �#t ���ܹ�#�<-p0�]�׷���  � ����|��Z���e���%���=�Z�r��� �t ��4��^��_���?��g���V�[�^�U � ��_�T*m:�X,~9^86����w] ��	t �W���'�
�B3җ�U�e�8��V��S�T�5 ��: ����~T��^���bL�n����%�\�/�� @�� ��*���644�?���?��E��tbb�_|�o�[�nk �#	t `����{xx��B�p}��L�,˞����77n<y���{ G� ����﫵Z��q�� ������} �o t� �r�|����k�,�\=�i���j����J����"�������������3"���thh����/ :�@ H�R�b�x���;��&�gw�P��V���\.� � 8`1ҿ#�1�?�rI`���|R���^:88�; ��: ��4�`����h4nhFe`���|^ooo��g ڞ@ ��R�t����oM��~L`:��Z�~�R�|8 ��: 0-���C�Y�5�IF`��=�4<<������ �-� L�J�r{�^?��h4��~R`�̉�y�����|�}	t `Z�J�-�j�丼6���E�{{{/��s mI� ӮR���ݞ���cX�-0]~�V��s�\�X ��t ����2F�Ob��L�<��?<<����� ڊ@ ��8��V�����Y�	�[� ����暗�X�b2 �6: pЕ���z}k���Qa���Ľ���oO�����/H ��(�JWV�խq��,�����ذa��֬Yss �-t ���T*���뿓������X�e��ƕ�7o~�y�7 hy 8�J���6l��[1.�.^>9�D<ǎ�8�e ��	t ��k>�=44tR�XlF�s,�����gJ��M��&�����ϦM�^6::��xyj��4uo�|o``��So��E	t `�\p�;������M��]������3� �,� ̨�����V�}�Y�.n��j�z]�R�I �%	t  	�8+�yxV`��@_�n(.� �$� $c��������<,���^�ׯ���O��#���T*�/lذ᥍F�����>k~< ��M�7o~���Z�@ ��<��^���<+=6��gm۶��8_ h) HR�T�{�ƍ/�6^��g�B�/���/�� -C� �Z�z�����S{zz6eYv^`_>11�.����!���N��]�j��8_��}���q��_�Tn �� ���C18�k��;�x����q�
 �� ���W��S�7��>�>44tI�� �� @K����|�^e���c�<�B�X�8Χ �'���S*��~�%��lbb�,˖�ɵZ�r�|c  i hI^x��b��t*ҟ���<o������	t �e�H�mxx�e1Я���xTq^W��^P.�� H�@ ZZ__�}_|�+���>C�ŁG5u�� �� @�[�n�֡����B3�_�%q_޸aÆ׬Yss  I h���;b��6F��b���E����?����$	t �m4#}�ƍ�����,��[֯_߷v�ڻ �� @[Y�z�������j�8���X,�� �� @�Y�v����|�e/
<һ6n���W�� H�@ ��T�����uC�|a`�,ˎo���c��t �m5#�^��:��������A�$G� m�T*mٸq��ccc_β�遦�lذ�7֬Y�� @2: ��V�^�@�^?5����#arr�8	t��t �#�J���P(�K�\:\�e+�=888 H�@ :F__����76����:;t�E===���3�$t ���J��V�g��zIZ!t�3�@H�@ :N�R�D���Y�����������6�v �q �H1��_�Վ��R�\s������� ��� @�ڱcG_oo��婡s�-t�$t �c6����V,o���(˲�޴iS�\�3 0�: �����wT��7���c�.	�g����o/��q �x�J��Z��2.?:���	`�	t ��\.__�V�,˲��a���� ���  Sv����===/��zJ�,�=�����#� �4_�q��U���߉�G��eY�1w�0�: �#�^���Z�vV����h�B�(
��ӥ�#� ~A�\��Z��?.�"�� f�@ x;w�����}e\>#t�,ˎZ�~�1k׮�+ 0#: ���=<<���_�G����$�f�@ �����R��>��`*�? � �1dY��h4��#B��9t��%� C�T�R���g\~0��,˞ �1 �q{챗�~��kb�>3��E�z}q�J 9� �8V�X1Y�V���m.����$�f�@ ��r��z��..��X�e���[�CN� ��y�Z��+C�����  �h֬Y׌�������`�t �}�z��=�j���,�6�:���  �!˲�Cz�� f�@ ��R�;�z���\��� ���  �����Z����<=�'�0C: �~���_c��e�ǟ�7 0#:���������-����
����	��t�"�f�ڵk����h9Y��m�ǟm��͛��;�� �!%� �S�\�1N١�}7m�Գcǎ����{�1� ��@ h\p��C���[�. p�	t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H�@  �t   H��,�ST�J��    IEND�B`�PK
     �9s[񐼛�  �  /   images/a4af1710-95e2-4b5e-9600-8e4d90487313.png�PNG

   IHDR   d   }   T;�   	pHYs     ��  ~IDATx��	��yǿ�������=uK @� !a#d!@0�A�B)8��VJ>��*�\I��8���l�vbLى�KBh.��B�J{��5GOOw�|_���JZI���z�UO�3����~�]�_?�P�T��L5 ��D2ՀH��T"�j@$S�d��L5 ��D2ՀH��T"�j@$S�d��L5 �iB پ�2H�{��LP�2p�c�����Bpp]>�p̘��a����D��@�o_uu��8hZ�"J���VnA����؊�w���3�2�X�s�i%�~��6�駿A�y�K!��-�%���L��B|
-�"���"�qS������f��wu��ἁ�e�6�4Ͷ���|��9s^�%�}���Νg�%�	Ӧ�AG��+�W��Z�o� �x��(�9��A���T|����s;�j����ѳ��;Rp�ٯ���Ȼ�^	���<�A��-�3�؁�B`6��Qv!*�q>
c�!���JV#��_|�s?��gESSƙO�K��)r ۷_�0���.j�͛�QU��V[	[y|{rAQNSUu��8�ʮ���ZF03s�_�����M����لy!̚�dR�@v�x���(��d[��`�t=�e�N|6��	Q��ؠ�yY�q����-9��9h-W���O�S��ݽ�;�޽ �g�%2 [�^�������#U��Pa�p�8�8�+�
��qިp��u}fd��Pt�m��Z����//X��RK�.t_��}ɑ�E���ï�E�H&�,e��뗛��Vɶ�\bL;����6��+EM�0��4�=�`,���3p?/crэ�x� ��;;�ܜHbvw̟�"D�H�P@u]��,���EW�Gh�C�/���r��z=��En�P��޳������k��&c&#kӴO �$����8YK
��A�)���@*�2(t �7_��NrS��'o@�qeP�1�aV�Z�G�X��gr����hR}���u��XlU���}����X�A�������[[������H�B2u�A(���J3��߄�������Q�d���U�ڄe�:'DA;�3���\w�cY��c������X�qނVGY��1E���\�׺^z��"D�Ё���X��rY_��8|W�뚪��ef�����&"/ƛy�]��U��+|!���,!y_+�b���v���ܹ *�
d׮�`�ѝS�U�A���1V�����MU��V.��eۯ����*h������y�S�<]�o@0��~�R����#W�ͻ;a
���|�|����0HT��V����Qձ�o%7���z���Ӆ*�b1�<s'������ �h*����(_�2�0U����x"+9wڴ���T��u֫�B�q㵠��p�-?��?�c�W|;�(�2�����p�����S,��8Z�%�{oN�r�Rh@����t��B0rk��U�l���h[l���]~dB�%.0�d���B�˥�LB�s`��,�����J��l�:���D.��l�%�	G"Rh@��tY.i>|A�a�燺+�̩�x?!�5�F����8��(��y��Lm�J�&wD���-�;D�G�bPu�&:��� D�Ѐ`%�� whCB��-��m���H�
�U��q��"$�OF�X�R�uM����/�)t�C�>ڠ�ԥB5�G�7��y��J�R�0n�$��B ,�1���*;�s��t"��5�9���~'U,z��0w�L�@�����eٱ����͖�d�4�TJͩX�����aR:�@� a���P(�����IU'�q���թ��f=C�9��BI��u|�T6�U8����Oa��n���2c`�M��5U�KfIdX'�[�4ya�P������x&c7��d@N\�bDk�ރV�<��gvw�-��{�	�I�Þ:��RU�_�*]c�� M
 ��4ݾb��D��\�d���M������q�?��u�R,*��6G`&4�A��(�LnK�-KI�㄄A��@D,������𣆖�F��o
�!Y�9��?��z#��{�:��C���4Q����q�ױ����-5�4�C#��)�rف��|�r�[��ϱ#����U�s�0���=aXՁC��:�/z�h߅֣a��XVY��I]�Y��O��{�麳m������K��;� LE�ajj�B�13�F��i���y�q�O�>�4t�[���b�׻.�����00P�S��MP(?�����O��а�V$@�3�R(xj,c
~L������nC_@�2�+j�;hG3	����o\q���=��"X��mK!_1�'�	�B��2���ɶN���t�Z�w���ϭV�	��xB����#�x��r�)�ሠ�����H�1gͮ]6mڇe�lh�*�W^�K����	�Nj>T�yaa9t� �Es�l_Ƙ��|!�uW87��
��ŋ�\�.�U��R=62��+T���wnF �Gh@ǃ�� ���t��O���Ӕ�:���nMG�a(4 �a�2��pP�����ňdh���e�<���&�ЀX��� ���î�QG(
ǂD8�)X��x'p�[�F뺗��X�x�a�!q��7�Ԁn�K��d��`�Z��qu�)�A'1Q)ڎo	�q�sJ$��kF����;�]]eN����A���[h)�uuZ��zc����#��P:�� L�>	�'��!���DB��*Yg�X�=����Z�3��p�#Դ���.,��Z��h���@�4X�U���4<���� ���%��ٶ��aJ���R"3e��10P21�Ы�K�:�P�:��{閖p�;���jc�O�!��xl�U�Y����l4?��؞���Pu�O��$�������)ɨ�w<䪀ww�i�^5v(J���|���A��[�&4 �L�����2���
v�f�:xag]d4#���PO�|8�sjX�����/x��<��=��
�������٧��t�O���r��;&���ahNXP��K%W��Χ,�C�Ac���tzώ����/� a)T�5mZA(T�A6�-�WL�r5+F��*�i�X4V��+;R�P�,��I�QR��-&���0dZǿLGk��ܐ�E0u]k���={��+Y2y��8�b��`��6QQ]]��Ȣ�?�k��8��!A���e�qi%!�Nĺ����:�ʨ�P�&yW��>h���hIYϣB�}K!a��0u!<���55]==�����
ӜMM���9��9u�rm�u? �����q^���V����/km�ST����91��6M3����Tz]h�kcD��<O�488�[�������jU�3OB~7����8�x�~B��,�:]�����ŦC:�����0����s�0%=�
��83H˿
Z�CGG	�!h��X��L�0EiLc< ���T{���d��|W�w�ˉ���"�s	�<I��mхB�<s׷w�n��e_�����/ףK�@o�����4����\l��aL�Tu�F�Ș�>'DY룐kS��i�[���׵��W,����}aY��BP*����C��a\���>E	�&��_B�
Hw�g���%صk,X��o���ݮ[�vr�\u,�1hl\��vh���13{;1.T�l#��LU���7!�$A����M���D/%�<.HeU�O��ê��>W*�Q�s�10p�|�z�B�Y��qX��o1N��6=	�}��\.�9�HU�e�5������iY���ta'�ҲB����*cP~SUrI�A���E�"���.m���^����$���|t���e�~������w���߁�[���SO��%7���t�������>� �v�G�
VB���������ןd��|��֗!JE21�����fϞW_�WUc�f�������`)�ĹEř��򉏬��4<cX�l�v]�Q��l��6����֊�U�BԊl�ڪU���/��Ex�|��g�ԺU�	���J�Ĵs7f]�cs��`�����K�G �h�s���w����L�v���oAE>u����x ;�@�O��1�τ\n6�(c���@��#S�l��^���,�pO��RQ�s��f,�@Lb���j�f!�϶��mI$��[���o��s_��g�M7m����c)r c��+�odع41�t��W3f��]�������2�����t�칡�����x�7�9�jP�`�0��'�5̈́�k�|�6�QRV��4-�wt\�.� ƞ<ZM�͍޿�,�Vp|�R$VaR�"'u�u#��=Id�n��χ���_����>yM( 	��L��2?�S&w�=���,@F��#E�g�-ؾKO&����+�.lc-I}�_��e��͈4"I��9clB.�)�g�'���i�Y�dӄ2�j��ݎm�����	�����^f�ȧ	$����YЁ�nl�Ñ��	�!����ׄ�v�Z�c+��;�=v���6Zm�R6(�:t��!��BP�����;h]�^�C��
���A`���؜�#�.�6(��L �C�����a�9���Q��=�nV�T@H��/��
���c�/c{f��~���{!jM: �C�������/J�Wb{Z+�ȑ�я{��!P����؞cS���A��nS�z�4�5��sB�%���n�h_�??��J�
�u� �$�J�?��c9PHo��VU(,��x����'��S!)���ߧ�sBX7��� r�k�{�kx�h�HMê�L5 ��D2ՀH��T"�j@$S�d��L5 ��D2ՀH��T"�j@$��'FS��+"    IEND�B`�PK
     �9s[t���?  �?  /   images/e2e2c934-b375-45fc-834c-534243cbf361.png�PNG

   IHDR  L  	   A_*   	pHYs  \F  \F�CA  ?5IDATx���y������ϯ�i��qa�x�DI<��D��x<j�5�`��db&;;�&3�f�8��a�hČ��Q'8:*���!�A����~[U��B74PU���������#������6    �ݼ�曓�,�'���<�4dȐ�`+&    ��K�v��`+	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`�Y?��^Ql<��vd��Y{F����w��/ʳ��E�|V,>��&��;k     �����wD��w�b��E���?���������ҏK?�
_˛{-�5������u�o     PӒ&s&~wX1o�~���J��l��~����;�<�k�;,����s:     �II���=���E�,��J>��l��/ߛ3O�y�ߜ������      jNr�d���}��?d��k�,bT4fOϙ���{��?f     PS�
&3���y^���KpuN�o1�ƿ��1��_�     �f$Lf��7�<�5��K��H��>1�8�x{�     @�H"�L�xeS䅻��������s��g^Zz{C @ɧ�AQ��������TvX,   �:�D0�=��E��>/��;o������\ T����-��'Q��~�X�O���1=    �P���w\٫�;�C���б�һ� ؉�i1 ��c��!�4P��~��t|1`��ߐhl<6  ���5�[��+�������r������l�KK���IGs�3
���������>��_^ ��/���Ē6��MS��g?	 �:�o�u�std�����ڏ�~�lwuL���U������� ;X�|�b<Q��G�g�X\:�g    ԩ�&�ĉ��v���Ǉ`��?�F^�%{m�����.�^��p��   ��������}
�跳>?˳� �@�����X2d�'E[��}"V    P����رo^^�k'ɣ��A�Nȧ�AQ�� �c����gg�cm    ���&y�V�y�$�,�i�[ HK�||,��e ��&.�$V��ã=    ؤ�&Y�3ߩ� � �����1���KG�M\�->_β(    ���IG�Ya'.� �[�B��<*�m���[���U�   `��:� @=�_��#��Jo7�ј��e��7   �NL ���Gk�qo�m�M\�~vx|+    �4� jL�B�y���������a��    �K �!��qA��O�����?Y\�?    �L0��?_�<�!�(|�B%�\�7    [E0���tv�"e�e����K��D��7[z��7�E1�d���  �v$� P����Ȳ�"e}�߱��l�s�=`��#�ֵu됍��Q(   v$� ���^�߾�F��9x��ح_�   �I0ل�=���!�G�]v�b{[�-����+�     P��i���>=z��������b�+���3�     P_�we��G�<'z�6h������"/vĲ7^     �~&��u��>4��_��~*V����X�"     �� ���e�!��/k��=0��x.     �� ���*�wVS�-�D     j�`R���٥�M]�     �n�	     �<�     H�`     $O0     �'�      �L6����-��|SSS���/     ��#�lB9�l�X,     P�      y�	     �<�     H�`     $O0�@�P��}�n�|�x�g�755= �X��]    ��&Ȳ,�������c��ˈ HDG�ϯ    �#�     H�`     $O0     �'�      �L��b��/v�~     ��	&%kWE^숬�Щ��W/     �~&ey�ߞ�{�۩�Wϛ     @�L޵�7�̓��Ȳ��׶x^��73     ��!��k��?�;/?�9�C��X�"�?�@eF
     P?��Y:cj�[�8��Sѣe��!�c�~�^z�M     ��"�l`�[��M}Dc�~�w����ߎb��.��Q�[[['v�w�����.     �{�e09��S�,���7u��g��V�ѶtA��F�,�Ύn���     @���`r��g7�^���Y�}=��J���Q     �-��`���z��5k��eٞ     �E5LZ[[��^�Ȳ�      �J5LZ[[�eY�O���     `�d0imm�j����B      l��&�ƍ�v��o     ���T0immb	     ��j&��7nt��7     @7��`2nܸ?��|B�e]ڳ$�c�*��/      tJM��[�,ۣ��]�;���|     �s�>��;�����[���m�3-�ɟ     tN���P(\����tu�yY���P�|     ��Uu0;vlyfɟl����+�bP���f�_     @���`R(.��1^}s�N	&�-����      �_��1c�����m]Nk�̷㸃����r�Z�<�Y�6     ��W��������Ka[Ǚ�tu��֒8h�n�#=>��      jC����k��~57أ_
;f�Iy�r�     jCU�Q�F���1�5ޛ�WƓ���<$��uŘ����&     @m��`��ܼO�Ow����sc���ư-�=���*ˀ     ��*�ICC���=fG1����o�ғ�A}�c{x����̜     @m��`R2x{�r��_���u��>�o��[,�,��j�w     �E�L�ۺY�hr���3>�w|r�A�e۶��5�⟞����4     ��T���[�/�PyFȿ<7;^�ݢ8���c��ty���b��o�#/��a     ��U��$��i�4s���~�˕幎�w`����^=6�̼��*���ߘKV�     ��Ue0��f�[Z9
YC���=���~}zF�r<�#V�]����/ZKV�     P_��)�y%��      �	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�@�1cF��G?�ٳgGGG���m��b�رq�)��.��     �L��-X� Ə˖-��3o��fL�>=~���	'�g�qFz�    �*�j��O?ݥX�~k׮��~�r���q��Wf��g�     �D0�����-�̙3�2�䦛n�Q�FU��G�B!     �`5�S��T��~�����[�[�n]<���c���q�i�Ÿq�b���    P��qMMMq������_�%�%�=O�y�Nm��[o��7�\�P��c���:9��c���!     �`u�w��q���w��E��C=<�@��������b1�z�ʱ��Gkkke��=��3     �`	*G�/|����^��N�4iR�Y�f�ϖc˄	*ǁX	'cƌ�^�z    @��R0imm=��2&˲cK��y>��~� jV9z��K.�${���O3f��Գ��R>n���=zt�u�Y1|��     �5[&W^yeaڴig�y~y�eG��Z�� �CKKK�y晕�Y'�'O�U�Vm���˗�}��W9ޛur��'Gsss     Ԃ��SO=��iӦ�Rz{�8�xo�ɟ�ٟţ�>?�p���K�z��Y'��'�tRe��C=4     �ه������y�_�9�d���g����_��I�#�<+V���+W�\?����/�8�9�     �FŐQ�F5���ܖe��]��\q��Y'�?�x%���⋝z�7��M����y|��ߏ�;.     �͆�$kii��X|�^�zEkkk�={v%����?�e˖m��<�+�M    �} ��7�/K/_�-(�������3×544    @5ZLƎ{D��;���͋|0~�����o����
�B�s�9    P�*���+�,�����ށMhoo�)S�T��z��g+�K��C������     ըH~��_}&˲�>s�έ�$)�Q��;�t�ٖ��=zt�u�Y1|��     �f�`���eP���V�MRޠ��瞫l��Y�e�;��q�	'DϞ=    �4�;v����$m֬Y���W��Z�ti��0`@�3&�<��2dH     ԚƆ��1]�/ȁ��r������J(�:uj��}o6I9�|�ӟ�ҟ%    P��<?6�����kq�����ɓcժU]zv�Сq�i�Ÿq���    P����,��],�	&Ĝ9s�X,n�����W��^�z�����~z�1"     �My�w@[�bE\x�1o޼n����&9��c�]v	    �z՘e���6eʔn�%�0r�'V�&9��     ��@�ʳI�8�8�S�w��    ��j�ȑ#cРA[5�d��w����ʲ[���    R%�@�+/�u�wtz�������L�c�=6�1     �oJ�0 ��o     [G0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&�-\�0�y�X�x�V=?p��9rd���'     ��`l�����K.��˗o�8C��;�#���     �F06�n��XR��oƝw��^zi     T�ج9s�t�X3g�    �j$� ���y��U,    �	&     @���ƍ�]v�f������_    �Z � ]֣G��u�]7{Oc�?^    ���o4    ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	ԉU�VŒ%Kb�=��,�    ��L��u�]q�7ƺu�b�}��뮻.�     t�`5�׿�u�p���y��Y�fŵ�^7�|s     �9�	Ը�^zi},y��	&t��k׮��ܜ9s�����s,    �Z!�@�kkk���]�˴i�*    @�L     ��	&P㚛��V��w    �"�@�;�â��1��ۣ�s�1    P��qÆ��|�;q����;�ըW�^q�y�Ÿq�    �	&PN:�ʱ|����<�M�>}���!     ��`u���%     �:�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O062��X�hQ�}Ϟ=c�������     �W�	��ڵk�+��������5�\#F�    �z$� ��y�Œ�ķ����4i��&    @]L��^|���V^�k�ܹ1lذ     �7�	�^[[�6]    �U�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     P�����+ؾ�\0    �jU��#�`{+&      �	     �<�     H�`     $O0�khhئ�     �J0�>|xL�:u�ך��c�С    P�`�/~�`2cƌ��ݻw\y����     �H0��u�]c	1}��X�hQ�\Ϟ=�������    @�L��ѣG�1"     R"�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @��y�ǓO>��̜93֬Yө��o߾��~��ȑ#c�����а~�_����#��+����N���wjܦ���s�=㤓N���??z��     �J0�:���W]uU%ll�r�={v����[o�5����e�]���b���[5f[[[̚5+n���ʸ?��c��    P��7�t�Vǒ͝;7.���ѣG,_��[�,�x��+��n�B�     �F0��p�¸뮻�u��r^�]ҫ�^~��xꩧbԨQ    Pm�qS�N���";��O?-�     UI0�W�a��,����|��/���k��/������k���?���f�1eʔ��ۂ    �	&P���cC�`r�%�ti���;����M^;�s��_�z444tz�9s�lL6�]    ��`T�w�yq��V6}�]w�5.��.�    �Z#� ������C�F�=    ��	&�z奼6T(    ��	&     @�      y�	 Uo���Wf��>�>�ڶ�X���y   v�<L ��mKz�)����b��پ�-֬�{  �'���У���Y� �OG���I�Ʀ����y   v�����<`us�9��Ӿ��j���}��  `�$     �`      �      &�z�{o��n�^�    ��	&�zGydL�<��:�     �w�	�^kkk̝;7��(�1v��8���    ��	&�zY��W��ո��+?
�     H�`lD(    R#�      �L������s��[�l{�G��    T�j�'?��J Y�x��s��zj�l\pA<���f͚�����q�y�    @5L�ƕg���?�c�v�m�p��J@9��sw�׊�Ç�]w��&M������    �j$�@:th\}��Qm��k���    P�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     ժP�B����v��	     T�����M�;�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L     ��	&     @��˖-���;�~��8��c���Q/^�<�H���ǉ'��
    �j$�@�[�zu\x�������>�gώ/}�K;�{-Z�(>���Ƃ*?�~��q�wİa�    ��&P�L��>����;.�(
�B�,�/�Œ�+VT���W_     �F0�7���έZ���LW�~�bg�;wn��    T�j\��Q+j�    iL     ��	&     @�      y�	     �<�     H�`     $O0     �'�      �L��eY������3�Z�j�s    P��q}�����'�|2�>����,Y/���F�w�}�     �F�	Ը�~���<����ҥK�s��\���s�}�Y�f�UW]��&���    �	&P�>��QG�>��Η���[��.�(N;��$ּy����o����g��ѱ�����hmm    �j$�@��W��?��&�-�?~\s�5q�]wU����?����l�TB�<�֭����=��hii	    �j$�@8蠃����v\}��zϜ9s���f|���}-?��m��e˖ń	�{�5k�l��}�K_
    �j%�@�8��Sc���q�7nr��{^}�ո�����D%�>�K��r����\9�﷤<�����F�=    �Z	&PG.���1bD\w�u���/o��g�y�����'��Ǐ���o���,��'Vf��7�ߒ���8��+q�W�^    P��3���{�L�2%n�馘9s��[,cҤI��c��g>�8��bȐ!�����C=����.���766Vf��7�8p`     ����ȑ#��c��ɓ'�-��o��և�[ެ�'?�Ie?����/�@���G[[�?�P(�)��R٫d��    P��c�1f̘8�����[o�u��D�<�3fT��ʲ�f��Tb    @-L �e��<��J<)�")�CR^jk[q�q饗�     �L0������=�β^����3�	��.� !���� fť�d-��(-�h圥�ǶDT��Cת�T��9�Ğ��p"��B�.nB�T@��p5W��o߽KN���f������{��;1����<����>���Ї>T�k�ܹ�v��m���������#�    �V �@�����s���:����?���)9ꨣ꟫�    Z�`�c�=��/�s�=7n���뮻b�����K/E___�=:&O�\�d���1eʔ     hE�	�Ǐ��|�#�     G�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0��v�����Q�FE�R	    �V'� �lٲX�pa,^�8{�X�~}�x-���q��������P    ��$�@�-Z�^{m,]�t���j<�������7&M�g�yf�v�i1lذ     h�	d��&ɕW^��w�6}���~����r�Yg�駟.�     -��(�WSJ��Z(��7�<����g�����1w���'�	    ���SJ.��hIEQ�w����w��ܩ�^�r�p    ��ڐ\O�`-�6�ȭ��W_}u<��#�LWWW�|����އ���W��U���7�1�\w�uq�9�Dwww���    h�!��O)@K��Q�p���%˗/�gj�����SN9e�7Dj�M����ƽ�����Y�bE\z��9Nj��9s�p    4�Z0�=�tf M��&ȗ�����;t�ĉ�2lT*�8餓�ˢE�⪫�z���k��K.�����/})�8B�    [{[[ۂj�ڟRj�i�b��g��>��[^[%�3t�q�W_~�����������׆�:��bΜ9��W     U{oo����*�O�)�_�>.�����%���?������~���__~��_���<��������_\�4�vX     4��Z��!�@Ӻ�k��~��{�w=�����P(��	'�P_js���Ƀ>��������.����!�     M=�̟?��������Tjo�\��[=7a�%��v�N%�{�{�S_���ַ���x�裏��V���    �h^?y�g���mJiT Mc�ҥ�z��-�|��q�W��ѣ�{9���o�\~����I6W�K0    �?����?:s��O����4�|�ɭ?���5�lTr볟�l�r�-�r��M��&�    hD��$,X���f͚�R�@S�ɵ5x`�Z4�=�`�f͚     hD������ݽ���o�hJ�rΒ�ho��?/QE     4����?�WgΜ�XJ�;�{ M窫��h�|��     h�otb��?>�S�loo�FJ�_��M��lm�u     ����N�t�M,Wg̘1�J���)�Y�     ��p�7��\�5{��O�[�nZJ�r�Т(&�ۣv��5��     `�P0�h޼y����ז]�����r�_     `lS0��ĉ#���zhժU�aÆ     h�	���s�FWWא=���D,Y�$     ��`     dO0�&W�T���`��p`C9D    ��L�����[�s�=cԨQ1���o���8    Јhr'�pBL�6-n���~ggg\t�E1�>�������>�l}̘1q��    @#L��Ն���׾�/�U�VőG���P[��^{ŏ~�����[�Z��{���7n\     4"�Z@mn�c�=6MWWW|��    �F'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {������{��{�1v��lo��j56�Uc�Kk�����g^.��     h����J��=���IcG�����W�?��Z��x�O/     ��2�EQM)��g��>��	1���bܨ����G�}|}y왗�ǋ�Ǌ�     м2���������=����W��gʞ]��ǂ�=�<��z     h>L���˕Je��{��w�ON?�Mv�J%E��o��cG��_?U�     �NC�����v�����5�c��������-���â	     4��&EQ<���9bX{|�}��X��a����G���x      ͣ!���G��ҥK�/7��{��ĸ�4כ���I�Њ⑕/     �2�̙3������r�C;�~O�~�1R��>vJ|e���     M�!��k�N
&3��7�^��G0!�z�      _���������.O)ۑ�L�0:�?*۴C&
&     �$6���'?yn֬Y?+7Oۑ����
���Ǝ��^X     @ck�`RS�T�Q���'����wL     �	4t0�������r����|�n�b���*�'t�_W     ��:��T��RJw�K۶~vϮ�1����-     �����d���̚5�r����Q�;b(��    ��i�`R�aÆ�>�������am�J��C�|     ``�"�,\�pMww��)7�ˈ�~.UR�����     ��4E0��?��===�U��)�a     ��4M0�����yOO���j�{)%�      ;ES����������V���R      ;��IM�M�3f���v}���      �MLjn����Ϟ=��u��}��=/�T	     ��д��f޼y��էzzz�)�����     ���:�l��ۻ�\����sR�Z��r�T��     ��d��������rʄ���٣�w|��?2      �DK��n��g�����u���m�|�}X���h�{վ�����e[����(�6v���Α��3     �-Lv��c9!*����bՒ��+/��*���7\����E���	     �4�������[��s��1qڙ����ņ�V     �:�׌�x�ƒ�R{G�ylO���E�?     �� ��f�w3���G���o{g�~��      Z�`RJ�J��_?|�~�	     ���T6""�_�6|d      �C0�نX�]�     M0     �'�      �L     ��	&     @���T��X�z�����cĈ�:::֗�@&:��    ��`���(b͚5[���l�`2u�ԗ�Շ �}��    v�     Ȟ`     dO0     �'�      �L6�R�O𾹎��      Z�`��J��ƍ      �	     �=�     Ȟ`     dO0     �'����r     ��	&��+���u     ���T���+/��ac����{*     ��!����G��SO}���7��5O�>     ��!�����7FL:(F�3�/*�Xu�Ϣ��      Z�`�QQ�3��1��=����69ݿ~M���X��      Z�`�:��LjQ�ewǈIFǨ�Q��^x:�>�HT�^	     ��&[�꟟��z.  xs�   h	�	  ۭ��-=�   �f'� ��*������_�����L��t������_�{�h����˗   �`@�K�����fAqw,�ߋM�����ѿ��tt�]@(8�#�  � L �����bI���_.��D���o���Ԙ    l� �L��%����q��������k.
    L0�&��և�:�ܜ)Fmv���ܨ��dP#   ��L �I���Œ�Qn�P.]���O�=�^񩔢    �)� �X�w���(��rw�f�ϋ%1��-�]�V��   �7����-R1���aP ���Q��X�J�S��Ǧ'��ƨh/��Yij�    lUK�"�u����SZ 0�1���8)����G��MOƿ.(�,n��iZ�    �������K��{~�x. `������]1-��r�m���Y1:���M����u   �&Z:�D%-��g2�� �tl,+�ɑ�r��ӧFG�/�ķ���_.w�#��    hQ-L��q��]يib�� Y:&���r�M��dL/�Nߦ����/K�45�   ������I�aI��'G�0 `�c��bI�\n�~��7�1Q�_�[�   @j�`RI麢(=�E<>��/��� �������Ҙո��}�N�后sIf*��Qm;#  Z��#>y�:�j������Y�����˃A���d������| R���6�#��K �ڼ#Ž1=6���D*�m��_$���W��y �V�x�%��(��ɱS>��#�����$͙S}�G�]Z��/�E�����oۄ� �����ruj�$��\���E_��L���   ТZ>��L9�?\>�+�>EL��L꙳6 �����P�z(    �B��64ֲ������W[��KVĵ����    @�"��t�E\>�YEQܒ"���(����vç     h*���f�G�]zZ��?FJ�w潋��E��'�3g}      M%�`R��s�c�.}Oq}��Νs�����#/8h��     @��.��L��7�>���~��ξ��R|�<4l;o�hJ�?N����     д�&5�|�sk�Յ�\w���T��*���m���jW�����S�;��      �Z��d�?���,W,���??~��'Eqr��H�ۋH��s���K�,E������>���     h���^{S��-     @F      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`     dO0     �'�      �L     ��	&     @�      {�	     �=�     Ȟ`    �PQ�SJ��x* ����}�
Y�    IEND�B`�PK
     �9s[e���  �  /   images/6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.png�PNG

   IHDR   d   0   ��ߵ   	pHYs  \F  \F�CA  �IDATx��{LGǿ��w��AN+Py\0!���hB������jL�6��h������Ķ�i�O����i+MK�6��FKm5)6& ����X�x���3{�	��=�N:������w�7��E'dnݺ5��9���T߾@�I��ڕ������D����	�\���`pA.H��I0��\�����O�&p.� 3�`,(Z'��Duz �v����%HFk0��G�s
49�&�6O�����LJ{f�낈4w�C٠iڛ�o��nĈ�	������W
����,���������x^^.T5�����;&Ռ6�",H�&����$�y��f
rV�oP<��b�D���^�Iϫ��?5��������)�#G��X��.UB�%�~�+�S/�Xh´��R�>��Ȳ��E���"�H%Z潷D7b���3#��P�A�[��}�w���L��R�$�:��ϜGEަ�����9^Mo�#�{ox��*!�Z��l�BOk��p���\HNIa"%@GD�#���6�(P����@��59�꼼�:1�K7�����Y|
oF�&�-��]��J�G��Oh�մxz)#b��>�������������ے	�]��wpbd����F�����?H,����?zoch܁��Q�>c)I�.��(��μ�}u[�}�����T�yj%�C{?/^��f������L�#�ʩ�YF�DBK|p�"��斖���������b�	�Z$����|jkk������!�.$k7L&�����ގ��.444$`o��#"A�ks:����@__233��א��$���鍺�n�#|�7pZ)�Q/kԙ(gϞEii)o�ç�Z5�����!����v���.N�|@�����a�?::�'N�b������N�yͅ�Ҩi����>W�~�F+U"�!�E#++K_�ĺ��,����	�j��(�`Â���F�c������E�����t�jCX&���\��{Y��.56��F}��K?����7�����ڵk��ƍ�	=�ߩ������l�cǐ����%|>+z���^��� V�^=o��:L���~ϡ�$����Ass�>u��ۋ]�v�� �}�-��(ӒN�4Ҭ�X�V466"99Y�h�b��ˢ�,X�������dJ���|}{��ˉ� .��gKs�?U�C�]B�c��]��hL�px�^4�N�<�Ʌ��e;��G�r���C}�1�F��hLVp�Ejmm��-������%w��(/\�����@]k,"�)�:+�Nё�i��#Q/��s�9,'`x�^C�|��:�C3)=g��&-�[6c̻�4j*-a"C� �9�/f�
Ց�Y!��<f�@_�D��2�&���^J��!�����P���]�� D�P4U?��<9QN�p�(nTVV"xߊY/�_��!l)�p\��['��̾�7������7m�2`0!�P�{&G3�(²W[��]m�)�#}l��wLL�®_���To=MK�iĘ�����>�����9BުU�<)�twq�`|�7�4o�k�9�:��a�FR��:�F�.�}k��oDF�3�L}�N�I��Ĥ��Yw#��N�q��V�V��T"� K�9��$\���`pA.HdL���{��X��aT��Z�    IEND�B`�PK
     �9s[F���Q� Q� /   images/028dc4b4-5e34-49e4-81aa-ecc68ea503ed.png�PNG

   IHDR  �  �   ���   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{�$Y]��߉8'ND�8Y�U=W��8"8�e����˂�<�a�6��(}����]�v _�/p��+ �E�gĕqaD�2�=�0�׺�-�?����������y�^��ꪬ8߮��ʎ��/D        c�e�C{y��H�, NV�:��r�        �8t        �ι��e٢1�"�^���Й ����}��gc�(����͏�       �L�        ��9w���(��pX�����رc�80��(��{�H��<\���6n���,p.       �kLp      �1˲�c�ڥ��+��1�_EQd677?20���_{��Un��X+����Ϳ�       ��      `����h�Z_������������	�W�,��;��^n���v���        @��       cU�G����9��$Ir�Խ���'��CUU}�(���Tn��؈H�����d�       D��       c�e�e���Z�q_l]ײ�������GN*0o�sc������n��vW��?�\       ��E�       ���Z��l�v�;'�{�QU������Yk�J��k�)���$IR�e�s��       �+&�      �8�.p�}k7�����n9r����HoLр�b������i�&{����ͣl�+       `gL      �1����Zn����v�}@D�1��J������o�Zn��V��Ƒ       pzLp      ��k/--�a�9�}�G:t��a.`n�y�D���0Ɯ󰟍��Çj�2       �̘�       #�����ED�4m-..�KG�y����{����ED�4](���Q�       ��      `�ʥ����[����v�����Y^^��(��:��/9����z$����<x���ől       pVLp      �*���*���$I�Xk�>˲��j���rν�(����ED�$�E�ԑm       pFLp      ���;��1km<�������������t��f�ʲ���zj�~�����w<x��7       ���d      �y��]���Ǳ�(��1�"��^��w�X�RqQ.����(����q�R��v�_�       ���       �a��$1�\d8�kkk/=v���ƹ0%���.��J�������<x�X       0�       F�9����ƽ�RJc��J����ƽ�`yY�_(��q��ED�8�qrss�kc_       ��      ���N��b�M&��p8�����[^^�aRk�j�Z_����I.���q�СCw��       0o��       `�E�+�,���DQ$EQ������\�9wA�պe��vk�EQ<b��      �<a�;       ������4��u]����Mǎ�t�����Y�}>�2*����?>|��P�      ��c�;       ���/&I��."����(�WU�9a�/fX�$��y�!��""i�^�h�       0˘�       �N����4M�n����}�ȑ#��^�,�(eY�y����V��""���v�#G��       f�|       �eY����F��ED�<���n�,t`T�<BQٔr��H��߳��p��9       `Qp      �s���+լe�i���nKDBgΗs�'�s�7�4�xFE��zW�       0��C      ��Yk#��k�܏�iZ�α�4M����"rI�,������E�fcL��"9.I����#t�dYv�s���      ���@      0E���t:G�,{h�,�.I��4mz�vI��N疢(�:�Wι����8�CG9�(�$�����1��4�!˲�[k�8t       �A�      �I��Skm�����Ox��TD�й�QQO�ֶC�8km�e��eY���Y��*����_hr�}���k�U�ṣ4M�^ŗZ���45ƘKCg      0�     �)a�}QݹK/�"���H��9���m�h�{�h:c���ߔ����8������aZ_ǧ��Q�sFeY��y���,����q�j�8      ���=�       $��u�Ǭ���j}�{�1�b�k�c�4�:�^h�#����sׇ������TUտ��r��4M�e�e�s̃4M������W�iz��J���      `��k/1      0��1撝>q|�����y���6o�,{�pED�8V���z�_:p
��\QWJ�βgJ)e�e��x�4M��s����O���~؄s      :       ��˲�Z�L��.I���~��g�;�C"�2�xs#˲��i��� �")��FY\^^~y�<��TUU}�9wi� �#M�:�.\]]�v�,��Z{����y�_~����8��D�      ��3      �!c���f��RJ��x`��9�{��͕$I�>��۷SJ�s�o
��(�}UU}m���""Q�$I�:ǌ�y���{���(�Zn��~����	d      0F�w�O      `�����4ݷ���������G�>\D��)��p���{��i/�o��ZVVV>������Y0�,��Z��<�}�,�2����}���w��2�$��Z�?�s���9w}}���~ؘ�      ���8      �6���^�(�"q�]s|��Ϗ#�<�����Rn91��G˲��0�$ɽ�,��,��E���C�r�9�ڲ,?��s�]DDk}�r      ���9      �(k�c�1�\@��j��o�e��sQ"I�|_�e��cԎ���WU�9a1& ˲�{��.M�4t�q������B�FƘ��eykY�/N���i��}g��       L,      ���־�|�E�Eq���ҷ������5O�,{Wǡc��s�ޭV�f1��`vYkW�ǭ�:t�q��X�e���9�������V�o��ا��]PB)%qs�      `�q�Y      ������4MG6��kY__�ucc���4��Ϊ4M/���8�g~����w:t����΂��{N��>W����`x�m��"�:K�i�����s��-�o��������6      `���      4[n��F�A���y~����܍���,�־k��""i��k����v�,�Y���9��y(����q�e���s4\�{�����.�b��vc�U#�       ������      ��r��xUU�?����~�p8��ر��k�i圻�9�M��\�K�v�k������F�,�nιWE�8�CG���S�s���i��?�{��ը���;v�ڕ��/�m       c�w      ���8�a��?>���4M�\ś�}�'�����."�$IE�W���W�,�^EQ��{?w�v�;��{��:G��Y����n��sn��v��Kƺ       ����3      �4�t:���bR뭯��v�?�����I��`����ۍ1s����VVV������Y0UT���/��	Q4�������w��\D���������(ޟe�w�}���恃�m"�      ��ݳ      4_�3�r��H�e�(��(�w����]��{��y.���cb��My�?>tL��(����j���""Z�,�7��X���v���y�O��."b��hb�      ��޻      4�s�!
�q��,���tgY�Љh�*M�ǆ�Z��{���sBgA�Y��g���'Ydn�4M�*":t��,��V���,D���(�˲���/      �Qp      Jk����[k}UU������$!�LZQo2ư���8����-��_��U�e�EQ\K������{���9&�U�G˲�y�g!�8~a��      �3�2      �����$��CDdsssuuu���e����QcL:H��u-+++�Z^^���Y�(��蜻 t�&��z��o�݊�0t�q˲��i��-˲4t�n�{�;���      `o�@      4P�e�cQn�ֺV����(�LD�k�s�M�}gJ)qν�{��BgA3�y~Q������3��,_:ǘ-E�,�ݔr���1f��K/�B�       �7�     ��Z��Rͺ cER��c��y����I�eٳB�h�(��(���� t�e��k���<o���ti�����Uu�4�񅅅o�e��8nֹAJ)������s       �
�      @EQ���N'I������e�)q��R��7&I�C�h:��E�,o�-��̌1�u��Y�1{��IY�7��1Jι���l����,˒�yNG)u}�       ��      @u:���ք�q6���ݍ���Z]]}G�,#`:�Ί���E�&ZYY��c��#"��Y0i��`QM��Y����m�~��i�����s�4��4MBP��_��w�S��      `���      4L�$ߟ$I���""���{�����^D|�<��9�k����(�{�Z�[DĆ΂�˲�i���Qn�;c�����s��<�/���,�7LC�]D$�c眻0t       �G�      hk틕���/FQ$ιk:��!��χ�s��4M�5{py��maaဈ0%y�eY��EQ��1fz������Αʲ�Ei�~�{mM��%��$I��9       ����      �����3�k����fY�_���y�"��'I���1Ͳ,[l��ߔ)��;y��ǲ,_o�T\\���$I�����9�"M�˽�_���u�2��TQ]:      ��c�
      �,���R��r>z��`}}�WVVV~#t�]�����4M]� ����n�z��?z��-��`4�<��,_0MS������q��p�������Uk�T�����w�m�%�s       ؝��!	      ̚,�����r���1&���z��:�e��B�9���Yk)��H�$���Kι��΂��<oUU��G(I�y�g���eY~��j��i/����qlZ���B�       �;S�S      �%Z�)5^TJI��E�ιC�9k����ySXkM��SţBg�9������,���1zI�4���y�+EQ|�(�+f�Ć��       `wfj�$      0�1�Cg5cLT��K[�֭i�^:�vy����և�1��1q��Ͳ��Bg��%�����?r�
΍a��EQ�0t��$��,�.��W�$��;>��
�      ����J      `�i��R��p|���eY�\��H#FB[k_�t���ZGeY��{���Y�k�,�/Eq�e������y������+���Y=��s�p\      �
q�        ����<Z��E�J��Ƙ�q�g�^�PY��xZ��Ϣ�;^Q)c��R�n�{S�<8�����\�e<.�Ok���7���߆�`��OQ���?*�㙾�՝?ԟ�v�_�      �����J      `��e��(:Ǥ���zuu�ͫ������o�Z��y�8�u�U]ײ����^����Y��<�5�2:�<���8|�Сv�������'�1�cmm�G���߳      ����      4D��>��i+t�I[__?����ص���LjMk��>EѤ���������j�؁�V������ʳ�;��I�g���s��Y���mR��=r�w,��      ��8z      4Cn���r��H�e��O{��XD&2J8˲7Qn����CG�i�[ѹI�$y݄�J�,{[����<���."b��.���,t       g�      ��<zǡcǱx���t�i�/ǹV��?�e�E�\�6�Xvn
c�bQO�Z�G�Z��Z�ֳ���yD���R+++?:      �3��      4����Bghk�k�Z)�����o��ܛ��&��Xk_?��gιw������OD)���       �w      ��1���)�(��,���x$��'�r�y�?0˲��r��,��V�$�e��Qn3M�n�Z��e�d��(7=Ռ1��      ��Qp      �kc\�M�$IZU�ʲ������c���(b�h(L	v��c�G��<��?*��y�{N^8��:[\\�8t       �Ǒ       0����t�3��E�N�s�9����VQߟe�գʆ��h�\�7�%IrqUU�9�mdYv�����V��bj�����_�      ��q�      ,������t���{�����^D��l#��wr"AXLpNO)%q��9~yUş�e��,˲��Aq?!t       ���      ��������
�c�c�7t�iE�8�Y\\<轿a/_k���4M�W6`�1����w����^�&M�g.,,�V���q<�h3Ek}Y�s�:�^���T�     ���     ��$�y�߼��p ��'��3�,���چ�1M�$1ι7�e�Y��פi�?�c�{sQpo��h�߶˛����XUU�Ȳ��#{Ǳ����s̉%��[:��rY����z�H	     ����     ��(ʕR�e�%UU�oqqq�(�_��c��~q��n��(��(�^\\��s��t�,�.���R� �|�izEY�9�m��n�o+��Q��sn�(:����$I�������mUU=�Zk�RR�u't6      4G�      �]���RJ�$)ʲ���������'".`�����Cg�fI��eY���j�S���t��;�֌�n &�g���(�v��^ž�(���j�-M�d��fIǏ�aYkW��-_���7Ɯ��7��Ce     ����     ��(2;}<I�{�}�����\Q��t�Y���3L;���y~�s�s��S>��e�Ã�s��������<ϟ�$Ɂ�,�Ǖ?Ο�z�p�lTl�e/k�ZG>T�����p8�x��      0��q     ���g���Z9�������<ϟ8�l�(I�k�$9���g��ʲ|i��:���""EQ�w��7ܛK)&ME�(��)"✻�{���,ߐ��'�a�(���zR�Ӭ(�}ι�t:��V���<�˳�|E��     �)F�      'DQ���S(�$˲K��z_��9��w¾�=�־�R�h��~IY�7E�,�~8t& 8I���{��4Mx�ej��EQ�����1�~eY~:˲oWU�k������Ҙ�     `p�      '\p�u��~�n�����G+++?#"��M6��9˲KC�Uu]3��a�=*�^/t�,KI�$t������zGo���V�SBeY�cI��&Mӻ�������>|�	#�     �ø      lIΧD�$IR��3��۷\U�gʲ�z��fQ���8t�YF)�y��*<���ֺZZZ*B�h8�e��Z�֑����;�r���R�a6      �(:       �E�Nk����_����������}`�fJ����Z3�@#P��<RJI�����:t��q�] "�K���I��Q=G(��H6     ���4      ��H��we�1�"ɲ쒪����t�E�D��G~�c�)�b�0�@=#t�&1����,?������z��vd��㘘     ����      ���qlW)%�ڲ,����t�˲|���q�5M���Cg  `�c�:CDY�=�,�[����E�c�X��SJe��.      fw      ���R���^�Zk��xʾ}���������q��P�1�:0iLp�4Z��j]:G i�e/k�ZG��zOQW��x/���JǺ       fw      ���R��I���Vι,,,ܼ��p ��'Lj�&Ȳ��h��2 ΅R<%a��B� �䜻�9�����r��ze��>�&v�0��B      �^�      ""����I�����    IDATE�dYvIUUh��G�s/��m ��Bg B`�{sQp�<���_��0	Ƙx�?�e�7��zz��zҏ�(��D     �T��      ��jm���iZUU��N������Py��s���(Qh"c��Bg�(˲�TU��v�����$IB>�k     `JPp     ��V� ""�Z���}���������ЙF�c��!����\�|�yǱ���@�#V�i�˭V�HUU�r�]��/�����$      Ί)	      �(�����Z+���,�ycc��n�g���>:��*��YM(� ����E"�W�s��<�/RJ��Z�dk�n��+�     ��D     ���(���vE��y~YUU�n��8�^&"S����'Bg Ba�{s5�L��z����@������֪����i���""��P6t      4w      l�B8���iZUU��N������й��sm� p*N>���Z/���@eY������n�?�p�$�k��bqq�:      ���;      DDD)55�4���{��}��������{Bgڥ�1&�u�5q�30IQ��,�:�.�4M��j���]ι��xz���~���      �l:t       4�RʄΰWZk��~@�e_����F��}���ڇB�:��(^E̜  ���8�AD�:���y~�R�Fk퓭�zZOL��	�      8#��     @DD�RS;!�"������>�n��8�~QD7�Tk����P���l�Z�FIk}��vb�y�����y~�����i:��v��E�3      ��(�     @DD�-���4M���^��tֽ�o:���ա3  ��i����B:�qQ�eO���������N�dz[���uM�      g4�-     0J���Wd�5���,---�e�Ik�U!�iz��:	� v2͓��QRJI]�/��y��V��\Uջ�s��q�.Js^�8� t      4�L�     �9��Zp4ƨ�(�j�n���k�cB��Z�h��笮�� ଢ(zj�u�4�"��?j�ۇ��zy�����n��z1t      4�       �eY�8��-q�s�<��lsssycc��kkk�YD�X_k��I� {5����^c���zJ�����J�d^���      �l�9�      {��U�3L�RJ�4�UU�Z��Y+��D���Z��ƽ�dLpo.���8�����2Q�eO���@�������sTn���_w     `�Qp     ��u}E����kmR��3����e�Ik�X��y�����4܁�i�_:�M�y����j�TU�.��%q�i�F�      ��8�      �Z_:CH�e�yH�e7oll|ccc�777?2���q�b
��wL	o.����EQ��Qn/M�+�(zU��O���y�)���      �l�      u]_:C�q,ι˲,�p��]���x����+Edp>��Z���" �1ՉƘ�i�[��%I2߭�m�RY�      h�(t       4¾��$�"I��WU��Ng�9�v��qs����Q��Q��i����8�[�֣���M���WUu��n�{�`��'SJ��      �l�      QuBgh"��Xk�������t�{��4M/��6�4}�֚�p  L�ԋ��%e��h�ZG[��[�s��q<�l3 	       ͦC      @#��t�a�QƘ�������olllܰ����]|��3��:t��Q�]i����Yk����ui�>�Z�x:�(�L�      h6
�      �(����E�✻,˲?���<����굵�W��`��k�>�  �<�q�#"��>��~d�e�����$Ih���'     pF\      ""y� �&�"ɲ����7W�s�M�:	?1ƴC���	� �IE����O�p����eY���t��������N)��      �f��      QJe�3L+��$Ib���ɥ�������iz��HQ�i�)� 0��(����Vy����ji�Zo-���8��}��R�6     �q	@      ��$��c�2��_��~���Й��������N=�ퟫ�z��l_�����}7�ζ���o���ۭ|۷���;�nR�;�Z��9��Zkc��x�������Y      �L�     �,--mcl� f��B�֟^�'�nWD�Z^?�$��m�ó��V���?Q���Ԣ��������>w����$��ey��\ ص����>|��s      ����      QJ���]l����w���S�z'Z���f8�X�to�P\߭��=]�}��(�����ޞz1����u�
�      �.      J�ݷ&L������Ϩg\s�m�O�����Nex��������I�������^�	 �S��R�      h.
�      �(�h+3�������)P�K�דn�d�Y�u����f������SK�['�i�۷���Ǳ��IS�)�8���3      ��(�       ��ZV�i{55�,����E��%uc�c����'K�������b��e{
��|�����      �\�     �\UU�P4�c��UZ'MbFa{I}k�(��g���{�'��l��	�      8-
�      s���_:0��
�ۧ�o�LR�B��S�{��I���h�? fC]׋�3      ��(�     �9���Cg f��海�y+��ۿ��tW,�i���[ Se!t       4w     �9���$t`�m/�����V]�2DD�����R�D���;�|J�V�      h.
�      sn0\:0-v�ȾUh����ي�QIE�:       ���;     ��SJ-�� 4�֤��e��p:0r�<��L��������,/�&QJ��      �\�     �\E�3 ��Zbg*����D�l��2N������[ ����Bg      @sQp     �sJ�*t`��
����  �ݓ]�O{�>�}��w �N)���      ���     0��.Bg �e{�}k*;�������v�Nz����;�J�$t      4w     �9Ǳ�������h�梘�wg�����;��)�L�      h.
�      HC ���"�N�`�N-�+�N���1' ��      ���     0�RI��n���'J�L�du]�8	g��	��1ϔR�     pZ�     �\E�#B�l/�RhƋ���l=��z=����EQ���d(�x      p�      4�V�s��v�NP �j�sߖ�ޣ(��$�����K����     ���     0�"��" 
� ����Wl�^x�c�I��X]]]�o��     ���     ������z���߼���Y	�i�1cW׵���2��4m�»��Ąw`Z�C
�cf��Jk}C�ORJ��ѣG�:     �nPp     �����Z{��<�,����z+�^����wVVV�'"��g���q�^hgB;8���w��I�����i��b�3h1��c~\k}�1&�z^��ظ9p6     �]��     g8���""Q��������y�׽^�`�߿���߸���I�5y�Z����΀ٱU�����`꺖~�/�~_D�,�k�%�"�Z3��6/�a�y�?&��k�y�1��z�ÿu]�p6     �sF�     4�Rj�t��Z+����\W��uιA�߿�����`0x�����	F�z�����0��>Qh�*W ©�Zz����lnn�(�o��)��I�R���0�bc��$y�1��Ƙ�֊�6     �5�    @�(�6vy;I�$N��2y^]�����������߲���&96޴�M)uY��.��u���Y@1rvm޷J�q�(�s�#4��R�� M�+�R7c�d���GQ��m��ZDx�    ��A�     4Q]����WJ)��&��kD�F����^o���}���~}}��"�K�)��L�M]�'
���R;�	?7@3'��o/��V��b�M䜻`8>5I�gk��5�ؽ�OU�5�     S�=�     ���p8�q|^M�(��Z[Xk���~�}��������������QީU�����<�~�Ĥv�� 0����$�tw�:@C�,���s�11�T�>�d0tG�A     �1��     ��뾈$�ܦ�Zi�E人��s������~�O��o����:����R� o��Uj0_(3C����Q�(��q:f�R�:C ��$I�g�y�1�B���s1�    �T��     ��람�ྜྷRJ�$��$�LD�7���y������yuu��Ddy\�7E�LΜS���D�}0�� h��p(��Pz��(�N����`R�4�R)u�1�IƘ��$�&|rg0    ��H     �H�'�OLEb�M��׈�k�����z+�^ﳽ^����? 38�P)U�΀��*���}��:t�~ހ�u��~�R�=�"��(t<L1�T:ø�y~�R�iZ�g�q|�$I������    �T��     ���#���k�~�_E�������>��v���}:d�Q����UJ���	 8?���""qK�b��	O������w��h��5��Ok]�q:�v&t      ����     �i%)c�2�\$"����{�^���}���GD^�������E�Y�=J� v�i�o1]���v�E�h�OLw�F)eCg8Y�珎���Ƙ�c*��y�u8�R<(    �Ti�     0��(��nd���twm��ZD^>_�e�J����`0���������9w���4t�����[Eú�CGN��$0��át�]���5�T:��Ƙ$I�|c̣�1j�U��r��p��     `�(�    ����8���9��xὰ����ι������7�z������+�ι�(�L�87�� Muj�=�c�Z����)��:4M�+�R7c�d���O�	��7��    �|��     k8����~*���Z/��uu]_����^��~��'�^ﵛ��7�θ����V�}�� @��C������S5�u~Q���S�$�^k}�1����iO��     8`    �&니�|(��c.������z�n���J������D�P�|QQvi���e0�(�3��()�BG�9u�;e����
�:�eY��8��k�y�1��z&����;     �23��     ̆��{�3�ZEb�M��׈�+�����z+�^ﳃ��wWWW�'"�ʣh66��R{��8o���T��ݍ1��椋9�uhl�y`�$�3�<�s��z�_��?     �$
�     �����0n�v���w�ս^�`�߿���v}}�"2����f�^j� ���P677essS�8>Qv�lSJ��/�8��7��6�5�4�R)u�1�IƘ+�1�<]1��kQJ��9      ����     ���|��VZ�E����늢�z�[�������766n�Z���9�7�V�}0�p8��t h~�i��QJIǢ��8��Y�QkkkK"�O�ڞs�By����q�;I�d�
��}�����w/��ey~�k�s΍ȪruvUwQݶ�a�mu7Ƙ�,���� &`��G �ŀ�b� &H� &H�0�%du˸����̪̈{��{=Dܨ̬��x�{���|>�Q�x���}������   6G�   8[9��Z�k-���b��O����G���~g]ץ�����������ED|���_������Z�Zc]W�v��	���{u��]�}���4M��q�z�ߍ�+���ӧ��4M��~��k���ۦ��Dkm�9   �"wx   ���{���9縹�9����VD��o}�[g]�g������ٳg�]D�o�凜~�����zﯦ��RF����l�=���.�����`���{�W�=y��_�����n����n���~� �.A�}�u   l��;   p�Zke2��^޿yss����|�A_������������)"�tlr���/��j�ź�QJ1�8;��lMk-�e�eY^Mu7�{�Zk���������t8���~�������v��{כ齗�   l�   �Y뽯q3:��v�������7��o�R��SJ��K)���t�������?3&��k�E�5�u����8 p�j�Qk��ҫ��}�ےR�����'O~5�����w����~��r�#�m^J���`   `���    �]`�RJq8�����#�wz￳,�RJ��R������2"�7:�%齿*��ZGǁ����!�ޣ����9�*�+E�����G��=}��o�����~k��?�)%;>   �Mr~   pv����o�4�zDDk�������Z��V�����{j�ź�QJQ�/�,K�N��1x��n|���� �v�=��u]K�yg�����Z�'w�^��������L    o�=   ଙ��0�i�I�蝙�\�����r�Z��9瘦)����3���U>�Z���   ��r�   8wSk�眵�δvx7�^��Zk���Mu�Z��W:   ��r�   8{���s6m�!Lk��a�;ע��L��   �$w   `ֈPp�Q�� ��S�w�ݫ\��R����    �:   �����\�R�i���0�^<��R"���!v���6/�d�&   �Y
�   �(��z�QJ�eYLk���
؂�{��˲�4Mq8"�<:�����   ��Rp   ����ej�Ų,Q�= �w�J)�s��~o�;��{o��   l��;   p��6�����X�5j��� �)�Zk��T��n����g��f�&   �i
�   ��K)��{Wt�}�֢��F�}t�*�怭�Ǻ�QJ�i�b���4��y��.9��1    ޙ�;   �	�ֺ����୵�bY���*� ����(�D�9��}���ѱ�sz�kDh�   �eQ   ؄�{	�2x��W�V �[k-�y�eY�p8(�s6RJ5�  ��(   l��)�OF���MU]�5Zk�� ������y����9�y��~����C��[   l��;   ��p�����g\���c�i���9���    6M�   ؄���2?���ƺ���  D�O6�����}�v��x���!    l��i   �V�+��WRxw:��j�Qk��sEw\k��O   `��E   6!��[k=笉w��a�z�# �Z���)�WEwLx��5g{�  �mSp   6��Vs��g\�RJ�����Q  �Y�=�y�eYb���~�Wt�^��׈�F�    x�  ��xY�p?㊔RbY�h��� poz�,˫���pPt�^��j(�   gA   ،�{����{5�]��a)��x�ƺ���܋�   � 
�   �f(�_�eY������>:��[�5J)���b��G�yt$6��)%�   ���   lFJIC�B��˲(� W���j��n������k���0�   �<w   `3RJ�=F�`��� �\�R^MtWt�M����    ;   �)��Z�9gm��Sl���k��)��Zk��   �(�   �Rk-9�����v �w����I)���   \ 78   �M齗�Ppߘu]c]�h��� �i�����4M��|N･�+   `��  ��Y#�����eYb]W�Δ"$lS��sE���_�DJ�n   �"(�   ��{��3��z�Qk�eYLl""lrx ���i�����_   �"��   lJ�Yc���R� �]ѽ���>�����i���    ;   �)9�<:?���<+�l�,\�u]����!v����+�{_|�  �K��   lJ�=�֚FA{�    IDAT��y��Ʋ,Qk ��z�1�s,�777��Y�t��5i�   ��,   `sZkU�}��Z,����Q�3�{�j���t:E���Dw.V����    ��],   `sz�k(oq7T��2�ס����~ss�4���=K)�Q   \w   `sZk�Տ���ƺ��1 lTk-��cL�777�P��b�   �nt    [TG������<ϊ��;����Z���6v�]E��k����"   p1�  ���9����]��5�n �KTJ�RJ�������w�+   ��(�   ��R�z�R�"��b��ՠ|�K�y���k�Z�p8�ng�pkZk�)�   �%q�
   آ�Zk�4iqܣ�Z,�� 	 pmZkq:�"�7771M��H��5"\   C�   ؤ�{�����b]ט�yt���GG �-���x<�4Mqss&�oBw   ��(�   ��{_C�����˲(� �9��8�����p8DJit$���   pi�  �Mz9��w�Z�y���::
 �(D_���F)%�C���ёx���5_   ࢸ�   lR�]3���cY�X�ut�J8!`�z�1�s��7771M��H�T_�X�c	   �(
�   �&�:���u�eY�M x'��8����������g����8    �F�   ؤ�s�+ռ�Zk�����Q 8#�C�wUJ�RJ�������{Wp   .��;   �U��֦iʣ����{�����Q  �@˲D)%nnnb���q����   �EQp   6��^"�0:ǹ�G)%�y z�# ��Zkq<c����͍i��;   pa�  ��j�����9w�v�R  S)%j����c��+�?��   \ w   �G��������/�������R�^���nnn~��ٳ2:ߥ齯�3���Z,����Q ��H���_�Lzss�d��C����~t�tx����K)n����i��jD��i��\D���|��>:    \:w   �G�4��'O~="�jD�;/�ǭ�x��Io����g��Rk��������R��v��N�?�G��f�� 研��it��r���i���x��n7776�<�Z�kǷw��|g]��O����4�����i�~%��ݜ�r�Os�i���9�ooocLl   �.
�   p�RJ���?W��9�-���8D�Ͼ|������[k�{�o}�[�ֺ��n[k������{���3��{�O��?�c�����Z��z-  ��RJ�Z�p8�~o��}뽯�~M�O�<y���_��v!��/��~m��_�9?��͜�᮸����ש�.��   �8�  �~�Z���n���֧iJ���/��?���������Z{�Z�8"��������=���[k�,�F���|��Q�y�ↂk1�s��:: v�ϟ����<�QJ�����.��Zk�4M�c<��O�<�~D�j������rο1M��SJ?�s�f��pW\�ϳ�ڧ���   ���   �����m�o�3%�����xQ��+�����[���G�5Zk��v,��(��Z��Z���w{�?X��E���k�u��]M����<G�}t  xc��8��������/��U��K���p8���)뿕R��i��bJ���?|Y^��c��!�^n��3   ��;   ܳ�s5U<�)��2��|����DĿ��|�����?]��#�wK)����������!o��e�:�Rk-�y�Z��( oņ ���c]�(�ē'O⊦�?��s���ly�_�9��4�RD�b��gr�L�4�M]?�y)�R:��5   \w   �g)�\J9��������W��!"������P�ﭵS�����WJ������Z����?���r{{��QoO�D�E��,���t  �E��s��ϵ�|�RJyp������v�_N)�VD���n�˽����v?�s~�sNwS׷�q�?O)�G�   �k��   ��vgYp_(��x�<�%����]	��O�>��Sk�Yk��Z�0"��������_���$"�}��˂�E2�����!pJ)Qk���������/�Hy���>���~��ߘ�����~����n���ϖ�_^7^��{7�   ��;   <�i�������l	~��}��s�/&3ޕ�?����{�k��z�?������{��/���{����t:�QD�U���~���u]cY�x�[�.�� �*��W�:��ŗ��Kkm}�W�y���/�R~a����4M%"~m��_�9�|���)�'�R^�>��   ��  �a�R��~���� #�f�����F�_���������7��[kk~!��[D��%�/&��/�?.I�5�y�����e  �w��onnb����uZk�\�xq�_N�)�<Mӿ���9��]q]g��#�0:   \w�   ���ޏq��7��rE��^�{����T���z�����ٖ�ޣ�bj; �f�ϝ�����t�i��ɓ'�O}���!�|�R�+���Ưs8���_���r���9   ��(�  ��9�_.��w�/K)^�8">S��*S� �'j����󸹹��^��u��w�#(�<�9�i   ��;   <�Z���8_����9�ǣr;p��J���2�����   �)�  �ò�k�Z�x<ƺ���  ���s3��ZKJ�0:   \#w   x@)�}�������ǲ,&Q0\Jit�7��#F��>�   ���;   <�Z���8��8��,��( ���>: �����QJ�+�R�   ��F   �+`Q�X�5�eQ� ��t:�b������������Z���~t   �V��   ��9Oň���{����<+�pVRJ�# ��Zk�G��y��OGg   �k��   ����lt_)%�?���Q  �����t:��t���{�{�d   �    �AJ�������<ϦID(��J)Qk�'O��4M��q��cJ�'   d�;   <���Tk]F���R���V�  Q�=��c��ls���|t   �v
�   �Hj��Fg�a�N�8�N
5 lBJit�{��k��h�!Z���{7�   �Sp  �G�RJ�ϗ��fj;  ���Z��X�ut6f]��)%k�   0��s   x$)�\J9����2!���������	K����    @�nt    �&��ۈx2:����)j��� �;I)�� ��J)Qk�'O��4M��p�z�-��   0�   �n�K�5�7�������  ���8�1ϳi�|�u]�E��_   p�  ���s�Ց��{�y��x<*� �!�/8���x����(����<:   ���;   <��������Z��X�ut  ������6J)��pFj�%�t�   xA�   Y�y�Z3�vC�u���[��()�� �9�N1ϳ�F���Z��   ��Pp  �ǗJ)�G�����c��g'��+�A �պ�q<md%RJ��  �3��   c�F૵��x<ƺ�9  ��j����m�RFGa�Z�R:��   ���;   �s��Z���^)�$G .^Jit��q:��t:9y�
��>�   �<w   ���|t>���<+�  �����Z    `,w   $缎��O���t:ź�� �A ���ϟ?�R��(<�u]�)���   ��)�  � )�]њ8������Z��( �hRJ�# �����<۬u�z�NV  �3��   ��,��,K�N'�  �s�u������Qx ���R�F�    ~��;   �R2�}��{��X�et  �L�Z�x<:���RnSJ��  ��`  ��RJ�R���#k����
�s: ��ns캮��p�z﷣3    ���   ��֞��pMJ)q<�.�j)�� 6g��8�N�cpz�-��   x=w   ,�ܕ��]!��  x�����uM�q�>���   �L)�  �xS����{���뺎�pU�� �D������Z��(����<:   ���  ��Z���p��O  ��f�v�ZKJ�0:   ���  �䜧֚1�������a ����� a��8�ȵ%��OGg    ���;   ���R��jEܓ�����r;  �J)q{{��c#RJet   �)�  ��h�ݎ�p	z�q:�b]��Q ��� ע����Qk��Pk]RJ��9   ����   gb���k���Z�G� �)�� .�Ͷ篵���   ��Sp  ��J)����Zk��h���  \��{���<��   �Y
�   pFZk�������)�8/�/p��u���8:����1���   �z
�   pF�i�5#���<���  �ٹ;eʵ�y�?�   x3
�   pfJ)��@�=��c��::
 lNJit��Pk���ۨ���r�z�=�4��   �w   83)�et�s�Z���$  ���{�N�(���r�J)�)%k�   �.�  �̤�v���/Qk������Q ���� �,ܕ��y�*��oGg    ޜ�;   ��Z���Ѻ�q<&�=��FG �J���trM�z�-��   xs
�   p�r�ή��eYL;  6�������u}vv  ��(�  �J)�J)����t:Ų,�c �� ��j�N�z<vJ  ��(�  ��j�=����(�@{  ಴����6Zk��\�Zk�9F�    ގ�;   ���s��i~we�Z��( pqRJ�# /N;��������Z?�   x{
�   p��Z�U��Z���h�!  pN�S��::��I)�9    ��   g���|t��Vk����<��R�^ on������ j�KJ�0:   ���  �����5�k�q:�"����FG �5�u�y�]݃Rʳ�   �w��   g,��K)��9ò,&�  Wo]�8�N�cl^���%   l��;   ������m��X�et �MK �nj�q{{����zL)�F�    ލ�;   ��i��~�����뺎�  pVZkN�zG���3    �N�   �_*�G��o��8�NQJ �NJit �@k-noo��6:�f��{Ji�   xw
�   ����+�+�  |��{�G%�7TJ�M)Y  �sa   0M��.��pWΨ����뽏�  �uԛ�ߎ�    �w   ؆TJ��"}k-N��R �R���{w��轷��~t   ��(�  �F����އ��   ��侮��(gi]�ga   l��;   lDJiW7�o����m��GG  ؼy�cY��1�Ѧ7�   /(�  ���Z����j��� W��~ x8˲(�F����s    �O�   6$缩s�k�q<G�  � �4: �`Y��gC�#"j����    �w   ؖ])���&��  ޺�&�GDJ���    �w   ؘZ���N�5N��� �{ �µOr��.)���   ��Pp  ��I)���J)%N��R# ����� ܳu]�v�q)��7�   oN�   6&�<�R����RJ���  0�݆�k�sv
   D�   6���|t�/2�  `�k+���zJ)�F�    ;   lPJ鬊��V� �͜�s \�kڀ�{6:   p��  `�RJ��z�r�v ؞��� <�RJ��|�%��{O)M�s    ��Qm   p����O��Rʭ�1�>c]ט�yt   ^��777����RSJO#�G��Er����   �F(�  ��{O>�������q7=.��2�g~���Rz9I/��4�Kw����0Mc��)��u.yb, lE)%z������Q��~���ּ�~�H)}�g��kꗿ�_�֋�_\���W�}�w��?����>���=F���V  ����m�   ��^�K)�ޟ�ޟ朿�s�ٜ��"�{���䜿�R�f��Ϥ���ޟ��>H)�SJ���眧��RJq��+�_�d��*���t�3��'������ַ�u�?� �y��.�<y2:�f�޿��#���K������)"N��~��~��?I)}�Z�k��RzVk�8�tL)�^�?z��   p�Lp  ����>MӇ)��M)}7������9��D�ϼ,���~�~�R�E��uE��GDD��+��E��   �SJ�y����ft�M��}�/�QD�_>""�����]I��/�����|k�Fĩ�>ǋ�����m��YD|�{�qJ���ڟ�Z�a���R�)��q���s>����0"�  �&(�  p~n���b���n��Fk��/K�?�s�^k�/���L���D�)�"���"�>��K))����B   ۳�kD�������|�=�[kw���{o���kkm�Li�6"��֞���{�qD������Q��j��)���n�O���?~��   ���;   ���?�onnn����]�e�j�1��Er �*�/ �<)�_�/ޛ����E�����ZkQJ��x<~��R  ��Sp  ��k�N�Y1��Z�t:)+���!�)��.>s����   xP�v  �^�Z?�����  py�u�y�S��,��I��0:   �M�  �{�s>�R��sp���xW�; ��)��6Zk=�\F�   ��)�  poz��l�����QA .LJit �Ⱥ�����l@���1��  ��Sp  �ޤ�v˲�xt�_k-N���   <�y����J��%���  ���  ���9��Z��w�{7�  �������18S��E�c`   x
�   ܫ�RZ���9x7�� ��% �=J�κ���oF�   �z(�  p�v�ݾ�2���۹+�� �-%�Wx��{�����Q8�Ů�et   ���;   ����ɭ��{����  p�\�Y���RJ��9   �.
�   <���~]�OF�����C�� ��	_DD�ZK�   0��Q   LJ�6��go��(��� <���� l�]�ݦ��Uk�(��S   ��s1
  ��I)�u]?��/��  ��Qr�^�>�9ߌ�  �uRp  �AMӴ��.�s�Ӗe�u]G�   �����t:���#�/v4G�   �z)�  ��Zk�����RbY�; ���
 ��֪�~E�u�8���  ���  ��K)�ey6:/�Zc���1 �ARJ�# �A�גW��V�   L�  �G�s^�Q���M��   �m���4�WJ�(��G   �P.L  x,Ӻ��q�z���   ��eY��2:��r�9F�    w   M�9�R��9��r; ��s��J)�� �������1�G���?�   "�  x\�����!��]�]�   ��pw��Z�{���RJ��9    B�  �G�sޯ�z;:�51Y  ��椰��{o9g�   8
�   <�����f�,����1 �B�n p�Zkq<=�oܺ�?��it   ���  ���9O����q��u�eYF�  �LJit .Hk-N�����Z�s>��   ���  �9�Tk��s\�Zk��<:   W�5�v��>�   �H�  �QR����!.��y   <�u]c]��1x˲�8���   �H�  �ar��R�qt�K�{������Q �r���WJit .Բ,ᰶmh����   gI�  ��z�
p����Z  �+�t;J)?��it   xw   �J)��u������<   F���xt����.9���   �e�  .�ԛ�n�eY�X�ut xE� ���$w?��Z�#"��   _F�  ��RJi]׏G�تZk,�2: �)���\���eY>�9F�   ����  �Y��iWJ�G�ؚ�Z�N��1   ৬�괱3�{�)%�   8{
�   ������/s��8��|  �l�����1��u]?N)�F�   ����  ��H)��u�dt��8�N�� �-�Q�+�4: W�t:Ekmt��Vk-9g�    6�,   g%�T�Uﯵ,�	x   lB�=N���W���QD��  �����    IDAT&(�  pVRJy]׏G�8g��X�et   xc�5%�A�u}�s��   ޔ�;   gg��]�U��5j�
 lB�}t ��ذ��^�Lv�   ކ�;   g��������<�� l\Jit �ز,Qk�j���qJi?:   �w   �RJi����9��<��Z   ���tr��#h��dg   ��  ��J)-݊wD�(��RF�   ���{���8:��+�|��  �)�  pΦeY>b�RJ��:: �{�Η� 砵��it��UJ9��s   ��Pp  �MӔK)W��n��<ϣc   �����a�ޣ��|t   xW
�   ���Z�����N'p  �X˲D�ut�����RJ��9   �])�  p�r��u]oG�xl�<Gkmt x'6h o��ns�=꽷��w&   ���  �&��O���Y�]��1� ��H)��  ��{�y�GǸ�~�R�   `�\�  �	9穔��9Ck��>   W��˲���i��9��   ޗ�;   ��sN��::�C;�N�#   ��[�%j�����Z�tt   �
�   lIj�}<:�C:�N�Z �[�}t�DJit �R�����`Y�ORJ��  p�  ؔ��r��!�R��2:   �{�y�G�ؔ�Z�9��s   �}Qp  `sz﷗6ͭ�j   ���eYF�،R�#b7:   �w   6'��[��ǣsܧy����� ��eY��::��+��9g�v   .��;   ��Rj��6:�}8�N��E�) ���FG �7r:�l����E�'w   .��;   ��Rʥ��G�x_�F)et   8;����yt���,˧9���   p��  جi�v�nv��B=   |�RJ��::������2:   <w   ���V�+?�N�# ����s�5H)��  om��h���qV�e�(���   ��;����݄Z���A�x眵V���荍4B."x�	jC1bP�jG�(�}A;6�M��ӈ�-���A��bK�^�V��]k��~�ac��gԮ]�j�9ޏ߯w�0��n���� ��E�n�׭s|����4M�c   �"���y��d���뺮u   x,
�   ,^DLeA�ܦiJ}�q   �T���'�4�L)��  ��Rp  `�""��u�OQkMwww�c ��2] x�0l�6�a���s   �cRp  `��ۍ�8�Qn��Q� h&°W ����n��է���u   xl
�   �F��M�3�cǱu   X�-ߌ6�ˈط�   �M�  �Ո��0o[���Zk:��c   ��MӔ�ah㢦i��U,   l��;   �}��]�[�B���7_zq ���x�Ԛc���
�   l��;   k��}��u����>M��:   ����]�1��m�y�:   \��;   ��u]�ql�#��J)��6   .a���?s�ZS��]�   pI
�   �Q�Z�i"��]� )%�} ����TJi����*"Lo  `S�  X����p�2�0i���  �'"ZG ��;��#<�RJ�o  �9
�   �V������ �����o��   �)�4��|�_G�3}   6��0   ��s�a���w��ݥZY  �K�!�RZ�8�i��9�}�   Ђ�;   ��u]�q��w�}��Cu �\^򚯈h E�5���1Φ��u   hE�  ���i�^]��J)i�K}   p2M�*������  �Y
�   �^�u�an/�]www��  @#K�U��Zs��o�  �Pp  `+n�x��Ct   X�Zk���k���q|�Rڵ�   -)�  �	������R�*�A�sp��|ED� ����>����   l��;   �]}����xT�  ��X�sz)�69�   W�  �N�k����.��#"?���q�4M���   ����ݥ����1>��p���R~�����RʘRSJ�j�  �Pp  `�"���w��."��w�/�����x����Xڴ�-��	 �`��4�c��s,���:"rJ�s>(�  �5�y�  ���w9�|�&�OX��   ���1u]�藼>��>�J�CRz  `�  ��8Mc�M����O�   ����kWWW����J�9缯�^��m�|��^�  �Pp  `""v�2{7�2����ݵ�    ��q�4M���Q�J�Z�UJJ�   ,��;   ��m�=��;�.�����_ |����Zښ ��x<������~���R���*�  0[
�   <����p�\JI�0��   |����áu�Y��w   fK�  �s��RN)u�C�Ք�?���u   �3Ðv�]�9��2K?UzO)�RʔRk�C��  �G��  ����v�?q8���~��t]�G����[9�!�bx |̩���D ���t<���u�(�qZ;D�u��Ү�z�RJ��[�u3��SJ�����K���O)F  `E�d  �1����(����v���?�u�׻�.�X�������= �777i��1�������[� ������ngܹ�ZS)%M�t7��M��������Rr   �m{m   ~�����wr�F��Î�c��u �=��Rp����Ϟ=kc��iz_z��i���S���I)ݶ�  ��i(   l�ׇ��O���?����P�uW]׵�5[��tss�: ,���|)����~��<y�:��|��^J�_�q�˷��=���u6   �C�  `�~y}}�����g�����6M��: ,»w��n��ӧO�n�k ���t}}�rέ�l^)%�ЗR��4Mc�����毦�~�:   m(�  �������]��ie���!���1 `1��K� ~��t}}�:p*������4���8�������   x|
�   ����?�s�gr��T�u<�������󪵦���Tkm C�}��������6.�J�-��W߾}����  �y)�  ,����@�����.�c�c���K�8�� �����TJi�x��Yr� �FD�gϞ�������7�i�/SJ�ٻw��v�l   <�&  ��\__����������ݮ3���J)���u X��Rp�;�p8�����R�8�S)�e)����R������o�  �O��  �V��/~��F�?�u���u�/v�]��>���i���1 `q��K� ~,"�ӧO�������a�q�O���j���۷o�r�\   |�'t  ��~��_�����;�l����1��ݵ� ���>_
� �a��.]]]�����ǿ��ŋ�n�  �s�=  @c9�:�M��F�5���1 `�j��#�L����-nq<_��   ��)�  �)��8�C� ��Q1   6����xd}߿�n�:   ��  0�k��K)F�5fz;   l�4Mi��1x$�0��K�   �<w  �����4M/K)F�7�� _�M(��# ���X��͉�t�"   3��  0#���y�[UJ1�   6�֚�ah�3*��Z��Џ   Xp   3�s>à�ހ)m   ��xt#�J�Z�4M���]�,   |:w  ���}��/[�ؒi��4M�c    3��}���0�#b�:   �G�  `�r�y���sl��k 8�N�-"ZG �E�!�RZ����"�|h�  �ϧ�  0o�4M��!�nG��  ���2�r�}�*"v�s   �0
�   3Qk};M��:�Z�Z���   ����L�0��Y  `�<�  �߮��R[Y�aR��i  �3�}Y�i�SJ}J)Zg  ���   "��8>W�>�aZG �U�^��=/ �\�4�qt���R�i��F�  ��y�  X���a���u�5��^	   �(/��_)�N��*�ܵ�  ��Sp  X����x<��u�5���f   �Y���[�5���<"v��   p
�   �u]�����9���5 xnG���h �K��5���u   �G�  `�r�e���9�����   |2{	����˜�u   �K�  `���z7�������tY   ��`?aF�ax�s�y   X!{   �����RZgY�RJ���u ����� `�Lq��i��RJ�c   ���;  ��E�n��_W��>��� ��� k����4Mc��&"�   V�  ��E�~��s,A)%���:   �P����}��Uk���W)��u   ��;  �
�}�+���   ��2Ž�Zk��yD�[g  �q)�  �D�y�����9���v ��Zk����h V��6�ax�s>��  ��Sp  X��s��]�sd�   p.�.�x<�:�lr;  �F(�  �K���i�����֭c    +a��r���u]�:   ���  �2�ַ�4M��̅k�  �s�!�Z[�X�qos���   6F�  `��Z���5�Z�8��c �fX~�WD��  �RJ�����iSJ����B   6D�  `���0<�zɬ�{E;   �Q�wx��7)��u   .O�  `�r·a���ъIj   �crs���Z�4M/"b�:   m(�  �\�y�����9Z��5 �0����# �*�}�:ª��<"�s   Ў�;  ��s���[�$�   �K���aZ�X����"��  �q
�   �s.�8޵�q)}ߛ    \����������v�s   О�;  �vD��v�M���� �}�: �V)�^���&�lR   )%w  �M��\k}]J)��<�aLo�F� [e���L�ԧ��)%o�  �RRp  ؜��M�����}��}�   ��LӔ�ijcQJ)S)�MD�.   �-�   �a�����q49   h��OWk��4���]�,   ̋�;  �F����E���  ���|ED� �z�8�RJ��WkM�0<��}�,   ̏�;  ��u]������9��U�   @k^��y�8>�9Z�   `��  6.�\�ax�:�98@   Z���6q<_��  ��(�  )�a���u�/QJI�8�� 0[�: l�=���]�u%   |��;   )"b����4M��<��� 0�� ����u�L�tL)��  �g)�  �RJ)�ܕR^�Rw�Zk5   �{�WJ�J)oÕ2   |w   ��q�/m��0��   �ⶹ{��:M�ˈص�  �2(�  �=9��0�[���`>�t6_��e�R�4M�c4UkM�0<��}�,   ,��;   ?�s��Ǘ�s|�q�   �Y��K��0<�9Z�   `Y�  ����r��oZ��9[?(   �k��;����˜���   |6w   ~R�y��u���o �O�# ���Z7�r~��or��   <�J   >&RJ7�4���|H���#  ?��	�  ?e�M���i��n�{I   ,��;   ?�+������A��֚��Y)   0o[��n����zSk�E   ��<T  �"b?��:�qc[��   X�-�c�{�RJ]�,   ,��;   �$"�0�h��=��`�f�>?�# �fMӔJ���xgUkM�0<O)�[g  `��  �d9��J�k?   �g�S܏����u   �A�  �����i�a��   �:�u?���_�v;��  8w   >[ι�p��k�i��_ �h�: l��J��0��9w�s   �.
�   <D����8����qS���_ |"��  ?m���f�ۈ(�s   �>
�   <HD�Z�R�Eǩ�m�   ��4�R��	��iL)ݦ�!   pV
�   <XD�izY/4�u-��   �v-}�{���R^����Y   X'w   �HD�k������  �a�* ��0�B�E�u��}�   ���;   _,"�Z룷χax�  ����Z  �RkM�4��� ��1"�   xT<  8���>��r;   �K��(�L�J   .@�  ��������%�   |�4M����Tno  ��Pp  ���K��4�R�7 �ђJZ[�� 󳔗�k��Z  �KRp  ��j�����6��>
   `�Pp?��:   �E)�  pv���\���   �M�5M�ٶOCM)M)%��  �(w   ũ�����q��� lR�^ �ќ����XD   pq
�   <���~�5֦��rx) ��L�4�5�i?G�  �&�  x�R��E�={*�   kUkM�4���#�#�K��Ew   .J�  �s�)��t�Ň���   ���y�#�}���:   ۰k   �e��')��9
�?4ù? xD����	��T �d��Tk����)[��������SJ�   ���;   �-"vq�c����n   �s���q�~�o�u]������ZJ)w)%S
   8w   >ɩ���Tn��bs��   ���VpO�~�{D���Zk*�����6u   �"
�   |LDē������Rp 8�/� ��4MS*���s�(��]JiW��Zkm�  ��Qp  �C9�'�ѩj)%M����/�� �p�8����:��{��Ҿ�ZJ)�i�;   |w   RJ)E�.��$�k=���v   `k�Rp����]�]���J)S)�RZ�  `��  �-眯"b�[�ߡ�   lM)%�RR��]ι�9?���R�x��n  �Qp  ؞��C���;1}� ,O��u~�e >b�S�("R�u��Ү�RSJC)�.�d1	  @JI�  `3"�p*�w��|�4M�#    4��}��s��q���Zk��  ��)�  �XDt)����n)S;�ah   ��i�R�us��DD:�4x�R�*�L��cJ�F  �)�  �O䜯RJ���:�'���RJ�  ���5! l�8�i�߷��Tι�9?=���ֻ�Ҷ��  l��;  �JDē�8�s�,ez; ,[��u ��Sp���H]��RJ_�RjJi(�ܥ�,<  VL�  `�"bWѭa*�4�   l�4M�����9GJ��Zk�����c�\   ���;  ���ON��՜t�Z�   �}�}�s��!�""���RJW���4�}l  �3�D  �Or·5�ڿk�A���Z[G�'�t		 �5���'�9w9�g��XJ9��LQ   X0O�   �v�9r�]� �M�   �^)%�Z�����>�/�Ԕ�p���-L  ��Qp  ����RJW9��V1k�i��   H�7{%��?L�9RJ��8�ZK����[�  ��x  ����*�����ڿC� �qmp�	 �7������9�t�R�*�L���   �Xn   `þ*��;]�}���~�-��S�?� ����: �jp~9�n��=����W�����W_�v�L   ��&�   対��_�����'O�����{��B ����m��u>���*��1 ��t}}���kc�J)i�7���y��_O)�n�	   w  ���ꫯ���������;��ީ�wLӔnoo[�  �@�}�����~�o �L��>=y�u�M(��������͛?���A  �F�  ������v�ɓ'��~���C��O}߷� ����MG=�9Rp�e�9��O����9�4��������o����W��   l�v  �y=����p8�������9��3{777���: p
��� ���ٳdpB;}���8���������W�<   [�)  ��={�/��=�u��>Q)%��ܴ� ����|)��r=y�����R�0����+o޼��)���3  ���  ����������>N`�t<[�  �D�}��>}�v�]� ��v�tuu�:�QJ�}���8������aJ���  �&
�   ���������p�Ӈ�����2wwwJp �"�޽K�4���(���={�,ه��q����l:	�    IDAT�0�ݻw�m�<   k�	  ���gϞ�O�<���<y��8L<�Zkz��]� �)�ϗ�; ,���u꺮u>�֚����q�"�_y�����:  �Rie   ���������w��?���r�<k3MS���m 8#��Rp�e����ɓ'�c��J)i��}���7o��ٔ��֙   �D�  �;������p��ß<׭���xL�0�� ��۷oS)�u>�ٳg������ӧO[��J)������Ͽ~��?J)�֙   �N�   ���_���v��q8���J�p{{k�+ ����|)���=}�4���%��K�^��O[g  �3O�   ������4Mc� [PkUn   �^$\��~؛��c��   ̝�;  �ID�j�o�ax�:��)� \�[� `��,�4Me���Ε:   �@�  �;��x<_�βfd`�j��#  ��8�xp��q<�Z_EĮu  ��Pp  ����r��ϫ�֣Pp   �<�V/.L���SJ�)%��  >��;  �O�9�i��h<�Y�ZS)�u �M��� �304`j��x<��9ה��  �gRp  ��]���07�����X X/E �9�7MS��E�u��Y   �J�  �gDD���x<�l�e�   ƾʼ��x�����v  �/��  �����}�?/�M�L   x�Z���L�}�:�t�R�Zg  X:w  �ϐs�O��b�&-����Z�  pi�: p&�����Zk:�/r�5�d�  p
�   �)"���7�8޴β4&��zy� �2܎7�4M�8��n�:  ��(�  <@D��p<_�β$
�    _��y��XJy��   g��  ����}�?/�Y�	�   |�Z��s;��SJw�!   ���-  �/�s�O��b2��g�' ���h 83{,m�R��x|�u�7   ��;  �Dľ��zǛ�Y���+ ��)�  �c����q��q|�uݮu  ��Sp  8�ӕ���x|�:�9x   8�,�5�m��uιk�  `�  ά����y)���p�
 �FD��  �Y)�:r<����4�  ��   �r��i�^LZ���O �` pY���V��Z��㋮3�  ���  ID�K)��a�k��5�    �e����q��e�u��Y   �H�  �ED����x��u���   �����1�m��m���v  �F�  .��t<_�Zk�,-8p h'"ZG  ����;��DDP   M)�  \H�u�q_�R6w��� �o��� 4UJiaj��x<��:C�  �@�  ��"b_J�f�c�,�RkUx   x�
|�q�a^v]�k�  �{
�   �ץ�n���:�%�$ �VD��  <�._f��Z�ۜ���   3��  �F�k���n䱙$ ��� ��Sp����*"��6   ��(�  4�s��Zǔ�jaZ   ��SJ9v]��  0S
�   �E)e����	��   �x�|�ZJMm  �7w  �8��Z���n9d hK ���˧���ZkQn  �?w  ������3��k�`;j��#  l����+�L)%V  ��Pp  ��(��i�n
�    ����ǕRFC�  �e�:    ?Qk�RJ9"�r�	b  �)t��)�X�7��  ��,�$  �����{J�� �Q��/� X,{0?RRJE�  `��  ��2���j�W   .��o�R���K  �ESp  X�����ܝ#   \����^T�u4�  `��  ""�ֺ�	TV �A� �o��0���1�d�  �
�   �)�Rk�Z�9�4�� �-�< �U�r���ZRJ%)�  ���;  �B�R��>F�   �2J)�܋���)����   +��  �P�C�Y2� `"3�-�R������n�  �B
�   ��ֱ��s�� �G� ��RJ�q�Sn  X1w  �勔R����s+�    s����Zk�����  VM�  `=j)el"���ij   `S־Skӷ�  X3w  ����C��A# �|Dp
 [����Z��r�E  �F(�  ����{�qV[� ����  �����5�iK�  `c�  V(��t�Zk����;   �孩�^k-Q�r;  ��(�  �[=Ms�엮�0 `���} �`-Cj�c�v�;   [��  �r�C��X�u�    K��{��}��z   ��  ���1����s�v �&k  ���&�)%�v   �  ��4ɽ�Zu���'�   ,�R�eN�U%)�  ��  ���R�ǚ��Ia  ��' [��}���.1;   �C�  `�N������N
 ��B @{Kڗ���Z���  ��  6*"�4���m4�6   �v��7sڏSJ��   ���;  ���&d�Z���{M�t�� �E�m���Z�R*I�  ����  @J)�R�����	a ��  ��9�k�_��  ��)�  �R�����%�9�   l�_<���dj;   �@�  �oED�������9�   l�4M�#|ϩ�>%�v   >��;   �s*�O����n�; ��ܿ� lŜ���%,H   ���   ������j��  �,�   ~��Tz[    �d�;   ?��r{J�m    �����|*�  �'1�  ��ҷ���P 6/�A�. Vk�� "��$wH   |�	�   �t?�����   ��\�Ľ."t   �I&�  l�� �l��j�
� �Q�   ��Y�&������  pY
�   ��S��   �R(����0��N��   0
�   �c}�\�� ز�w��YJ�=�o�+����%e  �q(�  l�c��s� �e  0/DХ�jJi�    _N�  `�""�Zs\hl�N   Ve�/ �����R���p  ؠ�:    �"���K�� �'�A ئ%ܿ#N�Z�   l�	�   ���ef�   �aM�4���j�S�,   \�	�   +]�r{J�� <�u  ���m�v���   ��   �/���Zۡ)   ���q�&�)�  �ܮu    �4�=Z�xo���  K1��" pakޫ��ENWk-)����   �f  ��y?�}Vm�5� g  @����   �E�  `Y��ቝR   ��le�&"R��;�   `v�   ��� �3|7 ����S�͚'"�z�����   �
�   ��8����t`
   �[ݯ9�u)�ZkUt  X w  ����R�}����� ��  ���E��R�`  Xw  �YZ��=�6   �y�_���b�|���  �e�?�  �B���r;  �u*u ���#]Dt�C   ��Lp  h("�����Y  ̏5ڇEDWJ�   ��)�  4p���4�o���   ̋����s��Rʱ�zl�  ��Sp  ����U��I���� `�N/V d���""�����>)���Z�֙   ���  p!9�CD\��    �BDD��YJ�L��.�TZg  �:w  �G���uD��Y��` �m�  ,�iE��v_�R�Rʻ֙   �L�  ��DD��뜳g/    .�K��s�E�/k��R�]�<   [�d  pf��OO��۷�r)L ��6 �3DD��'q(���Z�֙   �D�  ��"�I�uORJ�D �fx� `�J))��:�bEDt]��ܻM)��3  l��;  �D�>�|���   �Z�{�J)S)�&�TZg ����{W�$�����#bg5}��/�"��%P0��A�x^^ �p�fNuw����ήʪ�KD�G����Mv�u�]J�Z�/�#p  x��(9�7q�UX�  }:��K �U�KD|}�^���/��  8*w  ����󛜳s    ]��`y�J)�<������z�~ߺ&  ���   x���M�yl] @/�  8��Hq������/)���5  ��;  �EĔs�""Z���6   ���٬/"���UJ�zww��ҵuM   {'�  �Q#�M�Y� �]q7 `}��ʥ���y��^�n]  ��	�  |Z�9��9�օ��&0 ��  �.��~YƷ�<�^߶�	  `��  >9盜�к�=�    ~�>�>E�x�^����C�   �D�  ����%�<��cOll �ˈ pn�6mED�Rn���t�^�>�tۺ&  �=p  H)��u)囐     ����z�ޥ��n]  @�r�   Z�կ~�W���o������	� ��͠  �e9�2Mӿ����[J�Һ  �^��  ��7�|�j��e��,��:m    �49���͛6M��{�������7�k  ��  �����������o޼����E�}>C �~�Y �O����W_���~���|�����u=   =p  N��o���7o��󜳤    �����p���_���������o�����  �Am]   �ھ��;�㿯�^Z�rD� ��r��g��?|��/���� ��y�e?�q�����^J������O��߶�	  �w  ��~��_��i��e�� ���Һ��<�_"8����@����\ܗ�s����'o߾�_)�ߴ�  �w  �辽^�����n���  ��ß�z�p������ ؆�������z���VQ  �ܜ�  �Û�9��~�����s~Sk����HJ ^f!| `�lp߇��:����1�r�9�t׺&  ��� ���9����?���#�Z�к&    X�Kt}��9�����r���   �p  N'"jJ�/?��õ�����H��M`    �<����_�׿ln  x@�  8��s��������G!헳	    �������?�]J魭�   �p  N-"��2�����<����     �3�s��9Eĭ%  >ϡ	   �%�4��|;[�    ,D�  �yj�   :)��<���лg�� �G   �#}�v��  ^�w  ���<����ں���   ����   ^G�  �3""���?�&0    xG  ���  � "�    �G�om�  ��j�   ��~����?    �ӿZ�Þ��  �2lp  x!+    8�y��  V"�  �
Y    ���u�  �K�  `g��   pd���3�   �"�  �����   8����Rn  ؊�;  �
�    h-g��ך��r  ��9�  ��~����   p��4Zb  �Fm]   �Q�ow��	�   ����h  ��   9�6w    ��v  �~��  ��������(rv   ��l  �  @#�g    ��H��0ϳ�  @��  2H   `�   �Um]   ��e�x�?   �Q��   �W6�  �j�    }ѯ  `��  :4�s����   �/�5��  ���;  @��6��[�    G�_�3   �+w  ���aӔa!   @_�k   �+w  ���#{��       Kp  ؉�C��   p&g������b   �O�  �E�eh
   �g��D�i��   g!�  �s�l�2H   �^   {%�  �s�E���   �5��  `}�   �C���    xק9b��&   >&�  p@-�Y0   �A�  �=p  8�CL�S   �>��   �g�   ��6��1   z�O  ��9�  �Í][��       ^B�  �D�|��f0   �>�Oc!   �ϩ  ����   ���ԧ�S�   lC�  ��ܒ���`    G�G  ��9�  �\Dx
       肀;   �=m;   @{��h�y�`  �'��T  @^:p\*(   ���؟��.�  �O�   |��޶�   ���   {�d  �bl�   hK  ��p  `1�    m��   �w�   ,��    m�RZ�    �"y   �bl   hK  ��p  `Q��   ��7  ��9�  �([�    ڈ�   vO�  �E�RZ�    pJ��   ��;   �2H   hC_  �#p  `Q9;j   ��/  �8�  �(�T   �6�e   8�[   ��   h@O  �#p  `q��    ۳�  �#p�  `q��    ��   G!q   ��S   �%�  �Q�  ��RJ�    Nŋz   �.   �3P   ؖ~   G�  ��<�   �-w   ��	  ��E��*   ���b   8
'\   Va�
   ����   �!m   �*U   �!�  ���  ��RJ�    N�Kz   �S.   �0X   ؆>   G�  �*<�   �w   ��)  �UD��*   ��`   8�\   VSJi]   ��Y2   ��8�  ��U   �u�   p4N�   �ƀ   `]^�  �h$   X�+   ��,   �h�t  X�!+   �z�^   8']   Ve�
   ��   ��I  �U�   ���Һ   X��  @#Ѻ�M�   �C����қ  �#w   Ve�
   �/�ND�  t�i  ���   ,O�eB�   }q�  ���V���[   �z.:[�  �gN�   ���Һ   �Cn  �j�   �����   ��߲���<ύ+  87W�  Vv�p{J�6��    �#ྞ���  hH�  `%a���l   ���oC  `{�   +0����+   �2,؆  @N�   3�z��;   �2�Y���  �-w  ��t}��+   �2�Y���  �w  �t}��   ^O������  ؀d  �����   �ur�zQ���  �%�  �
�6=��;   ��x!�z�   �q�  x!C��p   x��~�  �C�  ��D�-c    � ��/<  ,O�   ��V�V/g   �2��K�  `9N�   lJ�   �e�U�'�  �z�u   {`0��X   ���W�"  �2lp  ���eyJ   �ej��n"�_   <�D  ��eC�u�   <O�Y`  �S�(   xDDx�yE6�   <�~�>ED��u   ��  �����Zm   x/��WD�  <��;  �ϲp�vl   x�R���N�  �i�	   RJ�N�2N�P   �ir���1ϳ�H  �/��  @Ji��_�������   ��V�����5��#"�  x�S0  ���甒��JJ))"��   ��Y�_h   <_n]   �^��,��0�Y   �/��h�  ��  �Da����   >��<��a��  ���  <ӇC*������.   �k�'����.�  �w  �W2�z����6   �gx�?6�  �K�   `%6�?�-d    ��9[И  ����  V`O �   �8}��lj  ؞�;  ����,��s   xD)�u	�aQ  @?�  00�%��    ~)"�7d  @?�  x803<��   �C�%   ���;  @c����
�   �̋w   ���;   �ED��    �w�w   �Jz   �sg��nh   �N)�u	   Ќ�;  @�"�u	�p   xG�  �3p  ء#��#��   8���   �Sp  ءy�[��
�[   ��r·\n    O%�  @7�  ����u	   Д�;  ��u�{D�RJ�2    ��  ���  h��X�   gUJ�u_   9��    IDAT� �  @W<�   �U��u	��  pO�  �zFD��q   8�3��yn]   ��   8������   gSJ�v!   lI�  ��y[   pN�!   ���;   �����_[��TJ���   �rĀ���   ���;   �z8��^��ݏ8�   xL)�0a��Z,N   `��  ����<��z�n�=k���   |�0�Kx��� 
�  �w   ��>t��V��H�����    ���Kv�<[P   ���  x����5����p   ����x����v   �&�  �""b�f)�0   ���pb  `K�   ,f�0zD�b�   ��J)���"   ؒ�;   ]p   ���*<   p  �k�����+   p<.�  ��$   �a/   p49�TJi]   tG�  ��	�   G3C�   �K�   t�F3   �h�:   �q�   �-�   �Q�ZS���   �'f   v���   �Q��   �&�  �n�   {��Һ   薀;   �a�;   �w����   �n	�  ������,   �_.�  ��I   �b��ƱZ��   `)G��ߢ'  �y���  ���`�
   ���   �e�   �H��yD�RJ��   �Rq���,!   `�   <[��mg   ��-�~�u�  ��p  �YzZ�Rlq   vŅ}   xw   ���p���n=   ����r>�x>"��  �o�=A  ph�0�   �`{;   <��;   _��.[�  ��E�iz=��   �w   >�����g   @��ֿ�uQ   �!�  �n�S)�u    �����  ��  ��=l�2$   zUk�E   z"�  ��   �r1   �O�  ��3,   zSJI9�  �s9M  �{�0��   tŅ|   xw   v/"R��u    )�w��RJ�2   `��  8�q[�    �R��   ���;   �`3   ЋaZ�    �%�  �aL�Ժ   ��lo  ��p  �0rζ�   �DDǱu   �k�   �'�  �Vj���  �+	�  p(�֔��.   �=�  ��L�  8�d   `k���  `N�   ���  ����غ   8w   '"lq   6�sN���e   �!�  pH�   �Vlo  ���  pHa�   �.�j���   ��p  �lq   ��=   ,K�  �Ê!w   `5��  ���  8�qSD�.   8 �  `y�   ZDؤ   ,N�   �!�  ����   ,M�   �!�  ��ED*��.   8�����   �w   Na�&[�   �Eà�    +p  �"�f5   ���   `]�   ��0�K    v��v   X��;   ��sr   ^,��ql]   ��;   �2��-k   ���8   �p  �T""�Z[�   쌞   lC�  ���8   �\�4y   6 �  ��D�'�  �'�9��   p  ���q�u   x��  �v�  8��0�   ���v   ؖ�;   �UkM9;   �6MS�   �TL�  8��H�0�.   �T)%�RZ�   �"�  ���ZSD�.   ��8��K   ��p  ��"�S�   �Gj���  @�   �^�5��   ���  @#��   ��-�   �O�ap   q"  ��R)ų�   @��4C�2   ��  ���"�u   @C�8�   @C�   �m   pn9�Tkm]   ���;   <0�-m   pR��  @{�   �@D�q[�   l��b{;   t@�   >PkM9;2  ��L�Ժ    	�  �Glq  �s��ew   �:  @c�<�y�[��j���Һ   `.���>  @��  ����=��>L����   p,�����  ��   z,�~��l'�j���    V���f   �!�  �#������5MS���   ����}z���k�   �aB  �S�C�ǆw����u	   ��J)��Һ�@�  �|�  ȐoY�0x  ��DD�\.���	��   �G�   �`��%    ��x   �)w   x�RJ��u   �+圝�  �c�   |��'��y>����8��   ;�|�������G   �^m]    �z8����!����qL��}�R   ����Z��_���zD   ���  �gylXy?�<� s�t{{����Z�   <CD�i�Z��k�<��8E  �vr�   ؿ����>��Ԟ2  ��q���/�s|~   lA�  �U|z��>��W�ϙ  ��8���͇�av   Zp  ���C�=���qL9;V  �������{��   p|&�   4�jϡ��H�4�.   ��aR)�u�f  `��  �ʞB凜4C�2   �O8���(��   �^�  нǆ��<����|@�s   ��Q���}����_   �+w   v�>X~�սE����   `�j���ں�W{��x����   ��O�   ������y���5����������   ��EDǱu�����   ���   �C`[�  ��4���5b  �w�u�  ���U�{�   GTJI�z�   �J�   2�c*��.   Nmϯ���   �   ����Һ   8�i�R���   �gN�   ޖ��""����   �)��aZ��j��  pv�   ��qS)�u   p*�4�.a1B�   ���;   ��j |�\�|_   8�i�R���   pN�   V�mgq��q   ЫRJ��u   �B�  8����!�RZ�   �v�W�z�m   @�   ����  ��4:~�?   |��;   ����7"�4M��   ��)��aZ�   ,L�  �Ù�u	�0C*��.   �L�#����   �6w   �ס��r�.   أi�R��w�v�   �t�?   4t��r   ��aR��u   �J�  8��7��Z�  �rΧ�@��u   �w   a/C���r�'�  `Ig�  �٘�  ��.��n�   ЋqS)�uM�'   p�   ��ކ�9�4�c�2   `7J)����   �%�   �p��s   ��.�K�2   ���  �k{�Z6MӮ�  �-8?��  ��	�  @#9�4MS�2   �[�0�Zk�2   �	�  �[G�VVkM�0�.   ��b��E�!z#   �!w   hlǔ�#:   ܋�t�\Z�   4`z   ��  �/��t��  p4:   �����9�  @J�֚�ah]�n��ܺ   X��;   t�֚j���   �f\ ��-    w   v��C�i�<�  �)E�p��_  ����  @G�  8+��  ���  ؑ�l#�;   gSkM���e��Y�&   ��;   t�֚�ah]   ��Eo   �!w   v�[��q�4;   �i���e��'   �)9   t*"��͍�4   �5�c*��.�P�   �;w   ���F�g�  8�a�0��    :#�  @��yn]Bs�ϵ  p(��4�c�2���   �?w   �f ��0��ں   x��s��əe>_   �J�  �.E�A�.�K��Q  ����4M��-   �I�   ti���%t�r��  �[�4�RJ�2NC  �=p  �K���9���Һ   x�Zk���.   蜀;   ]���/(��q[�   OVJI�4�.��Y   �w   ءq=�  �.DD�\.����  �w   �2�s�v�r����  �p;   �\��   t#"��!"��͍�  �nM��2   �Y�  `�l�  �W�8�Zk�2xO�   ��p  ���/WJI�8�.   ~��'��  ��   p �0   Ѕ�s���i]�0�s�   ��  h��ex�  ��"B��s��  �;w   �2P]��rI9;�  ���H���Y   xo   8���a   67MS*��.�'�;   �W�   4c���   ��8���ں   � �  ��J)i���e   p��4�c�2   ��p  ��0   `m��t�\Z��y�  �	�  Є�6�qL�0�.  ��9��   �p  `s�ۚ�)�Z[�  ��DD�\.��   ���  ؔ�w��%�RZ�  �A\.���q�Q��   �   8	�   ��5   �&Sm   6cX[��  ൦iJ���e��   z!�   '�sN�˥u   ��8�i��e�"!w   z �  �&H�QJr  �Yj�i��e    ' �   'TkM�4�.  �(�8C   �p  `u���iO�  �Y9�tss�l"��  hM�   Nl��Tkm] ���u�md[��*I������u��#G�CC�X�9F4����`��j	 X�9n   x$�;   <���(r  �7)%��  �E�  �8QJYz   ���   X��   ��"w  ��6���R2   ��J    W��Q�   �RJ�  ��ye   �2�  �9���p8��   �8W�  ��̑{Ji�   � ��!��Yz    w   �D�   �C�   ���   xS�9�ǣ�  `Ǻ���m�^   ���   xW)%�����   �t]]�-�   ���  �?*���tZz   ܑ�   X+�;   �W"w  ���   k&p  ��j���e���=���R   �Gmۊ�  �U�  �e9�<��l��V��c��7?��?��+���x�  lP۶q8�^w���O����[�   Kk�^    ��H���>�9o}�����拵�8�4M���Ϛ?>�/��e�����"8  �F����Nw��z���|��y�5�ۏ����w   �Fw   v��)����?�Ӆ��mJ�z!z��sΑs��b��y��������R�p8ď?�^
   !n��������9�8�9�����o�%L��k   ��   �	�/Z�)���5�������{/�_�w�4�I�   �S�4����;�������#~��c�����  `��>�   X�g��-a��  X�g<g[��3   �qw   �K�`BD   �m��>nw
   �$p  �Z�E����k[  �3���    �H�   �ֈ�$w  ��=���[�A  `�   �ݔR�*�   X���rr��   �E�   �U)%N����   x*m�F�uK/   ���   �ݕR����=  �x���   �>	�  �o�s���$r  �F]י�   ��   �6"w  ��s8����y'   ��   6"����"w  ��;Ѷ���    �;�;   ����=g/E   |EJ)�ǣ�   �-W�  ���#�R��K  ج��M�,�   �o#p   &�$r  �Χ�.���   �;�  ���"��xe   |��   x&w   ���8�mۥ�  �j9�xyy��]����m  �g�U   `1��!��[z   ��s���$��$_/   ضf�    ���]�EJ)����K  X�RJ�N���   �p&�   �k�6�����   X��i�#   OK�   +�����1�  xz��g:   �%p   V��///B  �)�8K/c�W  �v	�  �U�9���K��e  �9���x<F۶K/   `q�   ��R�������  �渽i���   �
w   X�g����  �;�{   �K�   +��q�l�ܻ�[z)   w�s���9�d�]�[  �6�   �^�u�R�����R   �����i�e    ���   ؄�m��{�u��   ���i�x<.�   ��r�;   `3��m� �-�N��`�  `{�   ���R�t:E�^�   ��x<F�uK/�)��  `[\	  �I)���9�xyy��i�^
  �����    |��   �, �5+���ˋ;P   |�WR   �M�.�ǣ��  ��4M�\eE�=   �v�   �yM�DJ)~���֥�  <����m
   ���   �B)%^^^"g/w   �H)��x�   |�+�   �n��u)�xyy��q�:  �r�q:���    |��   ؝��m�.�  �I�R�x<�����X   ��   X���p8��x\z  ��5M#n   �#��    ��4M���M  ��K)]7�ڴ   p?��   ��s����h�f�   ;�s���m�.�>)�dC   ���   ���c��8K/  ظRJ�N�(�,�   �]2�   xm�FJ)��s�Z�^  �1M���p�Q   �	�  ���4M��Ǐ1M���  6 �]�E۶K/   `���    x��s���D���  �YJ)�ǣ�}gL�  ���  �BRJ.�/�x<F�uK/  X�RJ���D)e�    <c�   ���u]�R�|>�4MK/  X���l�   X�	�   ��+���t2�  ��R�N'q;   �B�    !b  l~}6)���    ��Yz    k�u]�R�ǏQk]z9  ���m]׉�   f�;   ,@0�n��xyy1�  ��|7����\   `�   �`��m�#��m�^
  �Mr�6�>9��   �>��    X�����8��Qk]z9  ��t]m�
�����=   X�;   �_4M�����G���r  �/H)��p��q�   `���    ؂�R�N��n�   �����I�   �b^�   ��������  ���:V   6�w   �O*���ˋ��  ����G���^   ��\�  �r�|?RJq<���8��K/  xC�4q<�^    � p  ���S۶QJ�?~�4MK/  ����]�    6(/�    ���9��t���^
  <�RJ������4�  `��   p)��.J)q>�Ms �t]g�)   �ƙ�   `
��(���t2-  �]�    �ÕV   �;K)��x�a�|>G�u�% �n5M��q�e    p'w   �o�4M�R�|>�0K/  ve�XZJYz)��|6�  `9w   �f��q���4�?~,�  ؅�i�p88�   ء��    �A�4����tI  ��y��x��<�   `9w   �F.�s+���ɤI  ���8�N�4nR����.�   xZ^�   x��m��?~��i��^  �ZJ)����m�^
O$�$r  ���   �s������>.��p  ��4�;    <�;   ���i���9�q\z9  �
)�8�4.g   <�  �70]���9��t�a�ǏK/  ej���Z}} ��n[   � �;   �j�c���=�M���������i�  <��R��(�,��՛�)rο}l��J   �s�   Wk�ZkL�t0�i��M�D���8c��FJ�4w  ��������I���1�i���ǧ�"���X   `Iw   �ފ�oC���o1�������~�L�4�����%�aXz9  �-Lm�7�=�S�>M�����N   ,E�   |���N����������k����s�q<����\.�� `ڶ����2��7#ߺ=�߾���~o�g�ـ   ܇�   �N������m�p;���:��mM���|6� ���9��p0�����ߛ�^k�q��O�9����ߝ�"�    IDATC�-�  �c	�  `�n�����m��zJ���Vb�g��SJq<c�8�����  [�u]�m�4���i��uJ�zNy{n9�������_�,缹   ��;   �џn��n�������8�v}ۉ���RJ�N��!.��j�  ��4Ma�m�\�o���4�v�!�  �g"p  ����^'��v��{���z��R��m�������  �I�9����qY����y��;��>g���lyS   l�-�   pG��������c���z9�8�Nq<=.  X��m���E��M����s��)�o�   �ūI   p'9��L���?�u�]��g5M���\.����� ����x<F�fm}'q�������  ���  �������k|=I)��p��i�r��8�K/	 �'�R���mۥ��RJ"�o�   �!p   ؑRJ�N��!��� ��h�&��    �/�   �Ukм�i�(���r���^  ;�s�������   �N�  ����YJ)�C�m��9�q\zI  �DJ)����m�^
    ;#p   ع�s�N���>.�K�Z�^  ֶmt]g��
���   �#p   xm�F۶q�\��{!  �RJ��뢔��R    �1�;   �I�E����i�8��1���� `�r��͒    ���   �&�ZE�_�s����0��r�i��^  +�u]t]��2x��2   {$p   6I�~M�D)%�q���,�  "~'��+�Rr   ��   �ɥ�����r�aD2  O����!r�K/   �'%p    "~���!ڶ���  <��st]M��!    ��
    ��9��x�q�r��8�K/	 �o�R���)���    w    �VJ����0��|�Z��K �NRJ�4Mt]'l߸��cu   `W�    �Q�4�4M\.��\.K/ �/j�&���}'��   ���  ���,��h�6.�K� � ؘRJt]�������   ��   �K)��p����|>�0K/	 ���9��p�   �	w   `sj���/,���1�i�Nt `]r��u]4�K�    l�W�   ����G�9��c����%�q\zI  Oo�뎰   �-�    _VJ����8��|�i��^ ��I)]'���\RJQk]z    w!p   6E��n��xyy�a�r�� �m������   {"p   6��*�ـ�i�i���>.��� ��t]m�:F~r&�   {"p   �۴mM��0�����  wҶm�m9祗    w%p   6�d��I)	� �D�   ��	�   x�; ��I)E)%���   �{w   `Sj���o�� �c��|FJ)j�K/   ���   ������u�~�\9  !l��8�   �B�   ��Lt ��m�h�V�Χ��   ��   �U�C��m�݅� �3�=r�"���   ��;   �b���4M4M�8��r�q�^ ���a{�uK/�0�   ��;    �UJ����8F��1��K ���Rt]M����݈�  ���   �Qk =�RJ�Rb���\.Bw `�J)�4M�m��R�!�  ���   �!n'���1�i�Nt�  kWJ��m�i\�   ���*    ��s���]�E������ X�yZ{)e��$Lq   �@�   l���%�]�E۶1C�}�4-�, ��5M]�E�y��d��   ��  �M����yWJ)ڶ�-t�q�e O��x�q+K1�   ��;    ��4M4M�4��r�a�^ �c9�h�6���   ��  �M�Y9�8�Qk���Y �RJ���    ��x�   �]K)��p������!�iZzY �F�mm�F�y�    �.	�   x
)��.���q��; ��䜯���Y��K)�s   �iw    �N)%J)1M�5t ��R�a;l��Z   `�   ���9��p���b���>�iZzY ��RJ�4Mt]gZ;�d�;   �uw    �^J)ڶ��mc���\.1��� (�]י�    �
   �z&g�H9�8�Qk���cS�`�RJQJ��m����r    ��   ��RJ�u]t]�8^cw `�r�Ѷm4Mc3%    ���   X�Z���E�R���4�8�q�\�ֺ�� �O0�    �A�   �ZJIH�j䜯_Mu�m0�    �E�   ������ �^��   �v	�  �U��W�5�a���]�-����>C��8��`��h�ƴ���\.�����}�   �ew   ����8�1�c��"�)�H)�4MK/ow�n���}�8.�, ص��uZ{�y���I���8����y���'n   �L�   �Z��$�O��i��A{)e�e=�y
i�41MS�}�� �N�����mz}lt���P��(�D)�y�'��   l�W�   �U���4M1�c�Z�Q�G�v��c䜣���:�}��� ��s��m�iǉO�6x�ẁs��   �>	�   6��z�f�R���6O���a�q�^ ��3�m�[��s���Yk��g���   �~�   V���8�8��R���]�vA�rRJѶm�m{�����i��^ ��-7MM�r�u{<<M��9)%�   6�+�    +4�cL��4]'U�o��z�?�s��q�<� �������3n'���ҵ��cJ�   �w   ���)�q�Z�u�y}��䜣��.�q�abW ������=���0�4M�s���c   �u^)   X�{A�#'K����}�g�6z8b���>�aXzY p9�k��X�9=r����Z��n9)�]���>   ���  ���S�Tk�qc�kH�蠝�c���Nu�7H �V䜣i�h��1������K)�M�2Ǌ   �V	�   ����Zc��k����&�oO�4�4��16� �Fs��4�n�a�cM��m�>M���*�����   l��   �N�q�i�b���&��-j�%xٮ9�z�����J)�4ͮ&ask>^�}�������]u��   l��   �M�t���f�A�kk��8�; K��g���a�ZsΛ:�   �
�;   ��Zc�k0|;���u�>MS���c �j��7�펇�����nh��F��Qk�~�   ���   ���Hj��=�c��v�o5,�cn�����[�>M���`c��y#|�^�Co��c���k���R���   x^}   �1�cL��4]��yB��]�K�9�����8�a�q= x��A�|L���5����>�[�Z�����k   ��   X�Z�C�i��q���=j���DI�s,F�u����yJ{)�X�����.:9��9?�c�	   �}�   ��]�u�5�a������ͱ{�5�i����4-�4 �ټ�o����x�q����}�_�Kl(   �E�   �Z�5�q�q#�9gA��ym�n�qMwؙyz��ã�,�����YJ�   <;�;   �:_�����4]�-�����u�{D\����W��vS�46��
�އa�~��-   �L�   ���S?��������/�]�E�u���\���I�$h؞���yo���Y��L��   [#p   6g�3�P�6l��t�q��� ��)�D��:�ؗ�U>�1�1   �5^�   V�H�6޸�}Q;��<Mt6�]a�;�7��X�4ͧ�9�`�;   �Ww   `�ދځm�9G�9ڶ������w >G�Ξ���S�   �D�   ����v�{�����w��J)E���眗^�1Ω   �-�   <1�KI)E�4�4�^�|���
<���� A;    ���    �*�Nx���O��8�8��w`wn���il<�x�   ��;    �Js�޶m�Z����V�lIJ�?��<�i��^    +&p   xb�:�"���	��4��O�$zV�6f����    �ww   �'7MS䜗^|��6ͯ�9��}��� �0�즳��ِ   ���   ��x��Z��緢:�+RJ��Ub��|��b    �D�   ��F�YJ�	����Ͽ�q�} �k�ocv��    ���    x*oM[��������6b����j�    ��   <9�����RJ�R�mۈ����緾g`��)������     �!p   xrb]x�m�zk��>G�����`}RJ�Md���    X/�;    �'̱lD�6�}��>��'��o��}�>5�֩���   �w	�   �� �.�tlo��_���y�;�qs{;��6l��s     "p    �&�An)�:�="~����}��l��_���~�~   �O�     �'P�R��{s�>�&��'s�:G뷓�_�    ��#p    X���5����L~���_���s��:`�?     ��   <91,l�����������x������p]�    �=�   ����60�[�V?�������X���Ϗ)�:     � p    x2�C�R�?�v��_���X��(��Ƈ��x?w    ��;     ��$����G�u2���{����}޾���LX    `O�    ��p��a0��=B������oߦ��Կ��ޮ｀~��>�up�������s��>�8��    ,@�   ��D[�Uk�a"��4�����`�^�� �6C䜣�m��YtG��    ���    �`�����s'��m��)"~ݕa޼�s�RʒKۼ�k    �qd    ��a�r�D�5rο���4�8�� �����н���9��_he    �&�   <9��?��z��R��ߟ#aJ) lO���ߛ'�ϑ{�4��>�O_[    ��   ?C#a��M�}�G)�� vl����ω�y7�i��m�?nz�'�;    #p   ���1�i���uj�G�m  ���S�����4M1�c�?}�     �b�    1M��KX�Zk�}���ˁ�0w\ �r\4O~�\.���W�&�   �7&�   ��y�j��H��ׅ\ ����J�?gL͑{�4��    $p   @��8�0�s�{�&h����{���a�i��mۻ��    �Gw    ���圣��-������ ��0��禔���4]7�5�s^��Ǆ|    ��9_9   �7�6���z�RJ	��q���="���.�K���m�o��   ���   x����>RJ��l� `�9]|����Zk�mk�9    ��   �'0�c����i�o���=2n�5o��!j�QJ�R���    k��    �v�x��q>���9�E#�R��� ��y3�R�x��8�����bk   �%��   ���Zk�?C�5M@��iU� ~�q5���:.�K���iw�   �i�   �E05MS�}������i# ���r�y3�ab��h���1    �+�;    �6_9��L]}��9  ��k5ߕf��q�=�q<   �߬��:    fk��k���}\.���Ui�RJ1���  ^�q�%|HJ)RJQk���}�/�$    �;�   ��$�Z�5�����f x���W���Ƚi���?    �[�    ��8�1C�7n	�`}�||1�}���)ڶ]��m���   �1�    �64�C��s�R�^�]��69% �j��]</�����4]76ͺ.NӴ�    ؀��o    �a�4U��}�G����@�/RJ1����  ��������r=�   ��X��    �����є�*���q\�DU xV{���m�R��i�]ӦJ    ��U4    5�cL�)��Mk�^#: آgx^����a�Zk�R����u�   ���b   ����}��y�SSߓsx�
���T�!��Zk\.��a�%   ��   x�Zk�}}�GJi�ɡk!(����3Ou�\.���C6���   �G4K/    �u��I��8�0�s~�)�"� �`݇a�Zk�m�x   �E	�   ���	��a�i�"������"��y>�%�)��]f�   ��;    q����z�RJש��.�t�����Q����kRk���9�h��.�w�1   ���   p����>"B��A�8�Z}#�u~�}/��7Op����   ��	�   ����>��u�H�s�55���C�����Y�G�������:Q1���0�4MѶ��>    ���   �2N9g��?+��|'��19M��+�7�0\7��}���4m��t��R�RJL��0D�9���F    �˕G    "�c���xx�(+l���R���2v���kl7�9�0�
��^��9稵��|v��;��>ÿ��o/��owN   ��r   ����).��5�ݏ���j�q�\�}l��lM��o�<+��0�;��s���#�t�}m   �*�;    ���*���=L�������f�;�%�����R2͝U�C�q�|>�   �g��    `}���Z�5T���R�^�&M��װ���l��r��s�<�=����c�GJ)J)�=W7Ms�=    ���   ?c�����H)	�hǥ��)����w�9�:����z��/��i���3?�/�K�}��j    �
W)   �J)��� ���L����7_�:k7o2��9���Ϲ����9�   �#�    ���}�8~����kVk�R��R�Zk��g�_��   `��    ��9J������*p�j����+����_�H     |?�;    ,,�$D|�=����s�i�����ý79����a�^    �w    X��/������X�{Mom�����/�    X?�;    ��1������j|wp=��    [!p   ��9?ux8��Nm��R2�X�����^�i�?���    ���*   �:���ܞ5:�����aJ��`q��94�����)���    ��   �JLӴ��S�_K)E���o������[1��S�K�a���9秜��1�3��   �D�    +�D且%����R[?�01M���[Pk�a��{���3Ns�f*    ��<�3    X����#�%����R�>H����v�9.���+�V���s��sL����A��_��`���ɾ�w��d�U|�a){?�   �E�    +���pS��"��^s�{��w�X�?��n�m[[�(��_ q.z�&�cKE.�s��[�5�3|X��<��'��6�ϵl�����{b    �#�N   �$6��F|�G���QJI��F�}�LkMpz�Z�_����+����F��>��+    �J�    �D��6�R��Z���	�WJ��;\p��l�E���.�R"�:�}��W    ]�]%    ����S��e	;��#����������4��W�G�@ؤ�D�;{�w�����Z��>    �    .fY��/��Zk����p��y����9�!ڞ<X��D�QOS�G��>��1    �;L    L�a�u��v��R����t��t�[kԃ�t�u�y���o��k��3r�i�    @|���   ��~��i����kg�������?�$�=@k�4���$��|���i�5�M\^O�Y   �i�   A�0���Ҵ,�ٗ�mj�O��HLq����TJy�5�sO�Y)���w�O��������rο>�{�,��    :��J*    (z�>��v��s�u�5���Y�WJ��>�R�_���������^#��   �*�    �SF������q뺾e2rkM���Z���I���eY����QJi��z�    ���VS   ` )�p��S�?WoY�����    IDAT�����o0�>Zko�,��x�|/�S9^�R�RJ�<�ᾷ�u�`    �Ϊ    �R
D�<��#Sܿ���<�s��y~�Ͽ�R�[��v !��U4�No�h��4���    �4��*    t*�T�Lm�(��>�R��Z;�����y>$��9O뺊���J��h��#\    �<�;    �+Mm�(�|�(��$�#:��6��Z�S�SJSk͡��2���(�ܯt0��A   �G�[U   �!���rΧ��u��y����q�P�_�<��ZH)�?�Z;�;T���+�9{������   ��	�    ����Z�e't��.�nJ)��rο\�m���?�������t:o���    �/+�    غ���9�������&���|o��QuJ����Ξ�    ���Un    �T�S��"�|��=J(�i�v�W��P�l������9�=��    �g��   @`9�M�m����-���Man�M��=\��R�ܽxFk-�d��t��Ͼ��y����ܗe�    ��C    ��;B�RJ�i�Q�/39|;�p��ξ�O�/;�;�a��n�ۥ�[k-콈��ܯ���(��'   �Gؽ   �����Lm�U&��֦RJظ}�E��+��v8�
�e)��냎��    �G�   �&v�i�P����K)�y��kW����e������s�J)C��Lo�������     >g�    �K)�������n�e4�N˲t�ڸ�T��ֺ��G�ܷ�Z���4�W��e��    �3�   �?�Lm�ϫ"Z����}�s��y>�2N�kL�M������t��ξ��圧u]|�h��    \�]-    ���ӎMm�_Ji���[`���c��h��c�m
�h�)���i�w    ��    :�L�\J��e1��M�=lQ)ej�u���jA�(Oe�&u����~���i!�    puV�    ��L_����v�c�:ݳR�p��k�C<xDkm��֔��Z��}Uk�=ͣ�ܗeq����]   \��    :�U�gj��z��F= �s��y>�2�PMϑ{���yd��՞�     ���   �'�|�^X�u����M䎬�)�@�n�/����<�=�>�z���:���i�    @��\	   �}[�����+���ތ:����Ұ�k�uظ�w)��"���%�[�䜧eY�x���.�   �+��    Y�eZ��W�,�<Gι�w�ߟ��vw �;�������M�����پ�i�=>Y    ��uv5    ` ��iY�K��Lk�rq�4�s���8�QW��s���~?�2�t�C�圧u]�}z    \ѵv6    �s��˅�Q���Nq�jܾ��na�ͳ�����c��
���� 6p   ��Yy    ���Ykm*�L����K9UJ���ε����m"��     �!p   � l"�9O�ֳ/�u]M��M����u]����圧RJ��G)��4     ��.    ��L	_�uZ�Et��m�w�j���o"F�     ���    ���/�"n����6�Rξ����l
�'���هJLo    x/+�     /:3�݂_��ߥ�N��UJ�!�4�Z�eYN�S�    ��*9    ��rΧ�����&n@�5|��K�����i�9     ��*,    ���mK)SJI�����4��ٗ�Z�������Z�j�����I     �@�    ��#����,�����6�Rξ�O��l2���Z�# <q   �X�   �!� �;"p/��l_�R��u=�2�����v�㈃�^7     ��b    ��wOq7�}��0��D��H)�5r7�    �8Vc    v���}�g��Nr·L��Nkm��:�����4��[~��     Ǳ    ����1lkm������E��K)���r���~��g.��>    Ȋ,    ���
�[k�<���v�����i�����s��v�����2     �9��     ;�9O���~Fkm*���߬���z�YQ��䜧y�_����=9��   �]��    �,����u]�Z��� 9��&�?��6�Z���a�Um������v    ���    x��Nq��v�q����yvp�@�D    ���,   ЕW��)��t4�,���$)�i]׷����v�����r�S����kz;    �9�     �IJ��9[�kr�yj�o;H�ޞ+�4�Z��4    8��Y    �7yt�{)ej�	�O�s~z��#ZkS�u���sr�Ӻ�E    �G�    �F�Mq/�L)%q{��K)�����:p����t�]O    8�Z    �7�j��<����RJӺ���,q{L_E��    �˪:    ��}6�]�[���i�˲�t5�m;X���Ik͡    ���=    x���S�Mn�/������h�M˲���}|�B)�=    8��   �Ϋu��Z��y6���D�&��#�4��lz;    @V�    �E��群��u]��w����9{�    @V�    ��և��,˛��w�    ��     ����TJ���k�M˲�     /�    �7��K)SΖ�8�'P    ���     H)M�~����    `V�  �.�R�j���Z�夫    ���    �A9穔���֦eY��҉W     ��    �~��K)SΖ�    `/V�    �I)�i�gq;     ���;     �@k��K ��|   #�      �7(   �c�          A�   ;2��X~�       c�          ��   vf�8   ����  �8w           B�      t�D���]  ���           � p  �70�       �'p   ��0  p5�   �L�   o"8   ����=   O�          @w       ���v   8��   ��f8       <N�          @w       ��'�  �y�   �f6�      �1w           B�      ���$6   8��   `s       �'p      ��u   �@�          @w   8�)p       �5�;           !�      �<O^  ��   p ��       �ww       .́t   �C�          @w   8��p       �9�;       �� :   �"p  ��<      ���          ��      �K�5   �G�   '��       �      p9�  @Lw           B�  ��L�      �	�          A�      ��x�   �%p  ���T      ��      ��   6�;   `s       �           !p      �<A   ��          ��   �0E      ���      0<�  �w   �f;       W&p      `h�  @?�           � p  �`L�      ��           � p      `X��   }�  @@6�      �"�;       Cr�   �#p           �;   e�       W#p      `8�  @��           � p  ��L�      �J�       Łq   ��          ��   ��s       \��      �a8(   }�  @l�      pw           B�      0O@  ��	�  �6�      ��      ��9   c�          ��   :b       #�      �5�  `w           B�  @gL�      `Tw       �� 8   �E�          @w   �Pk̈́:       ��/    ��;   W���   0&�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�  �v���/       ��       ��ɠ   �'p  �6G      ���       
   A�  �al�   �d�  �(�   �f)       �7w       �0	   �D�  ��l�   �`�  �h�           � p  ���   ���   	�          A�  �iL	   8�u   ��  p*��       �F�       b�    �	�  8�MU   �cX�   :�;           !�  ��0   ����  @�   �a�       �M�       �3X   �^�  �f+       \��  �pD�    ���  @O�       0(q;   ��  ��W       ��;       �    z$p   ,��       p-w       ��   �J�  @h6c   �c=  ��	�  Ϧ,       \��       aP    ��  ���    _�~  ��           � p  ���   |κ	   ��          ��  ���F   �'�%   �D�  @wl�      ���       �)�    ��  �.ټ   ���   #�          ��  �n�R   \�u   F%p  �k6s      `w       ��   �L�  @�l�      ��   A�   \�5   F'p      ���  ��;   ð�       }�      @p�  pw   �b�       �%p      ���  �J�   Ǧ/   0
�   \��  �!��      ���        �  �"�;   ò	   �ʺ   W%p           �;   C3�   ��   �L�          @w   �g�   ��   \��ξ    8��a       ��w       �}   �  p!�5�   @H�,   �w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�          ��          ��           � p           �;           !�          A�          @w           B�  �W���/       ��;           !�  ��)�    <�z   ��       ��  �*�;   ߲1	       A����w?-��Y�Ͻ7"��l�����O��ͬ\.ܸ\���r>�nu'�Bt7�Ѕ��a`GQ�g�q����?��q��E�M����32"�=�<�$�m��ǹ  "r   �m�  �w           R�       [q�  �]�  �`�       �>	�  ؈�   ���  �Kw           R�  �1W�    ��N  ��	�      ����  ��;   �b�	       ��  �G�   �&�B   ��          ��   lŵ.   ���=  �}�          ���  ����       ��          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�  >Sk���    �Q�	  ��   ���   �}���  � �  ^�*r�m    vB�  �p��   dT_m����Z�    &a;  ��\p  x3�'    �Q��   �#p  x�Z�E    �o�   �'p  x )    �!�%  lG�  �@S    ���$  �n�  6`A    �λ!  ���  6dY    L�  ��  �|n    �F  �{w  �-X`   ��q   `�   [��   ���=  `��   ;��c    IDAT`�    ��;   ��	�  v�g�   �xy�  xw  ���   ���  ���  쁅    >�|   OO�  �'�_    p���  �!p  �#�/   ���M  ��;  ��   ���   hO�  �D,�     /�w   9�  ��%    ��j;  @.w  �'fa    9x�  �G�  Ј�    ��}   '�;  @C�h    ����  �%p       N��   7�;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )� ���Z�~c�9     b�Z}�z  ��f�   ا������~����Ϟ=����Z�    �R�����.��[�  В�  8z�8�~��?�����;�����[�    Qk���������GDm=  @kw  �d���O>���Ϟ=�����_���L    �i������.//�k�u�y   ��  'g�\~�\.�����x~~��]�-Z�    ���j��˗/8���,   �� �SU���>��������?���    �[)��ŋ߻��y�z  ����   �Tk/..���?�nD�0    �������H�  �v.�  DD)e5��뺾����Z�    �Zk�RZ�  p0�   ��Z�8��]��^��     ����   �p}�   2����q��|    61]l/���  �w  ��(�D�uw?     o"j  ؞�  �+L��    _f��  ���   t?t����8    @cӛ���   �#p  �P�5�q�   ���  �  �����    NG)%J)�  ��w  �-�R""���躮�4    �>�Z��  ��;  ���R���{�   �c!l  xZw  ����8�Bw    8p�v  �6�   {0���֣     *���  q�  `�J)�u��    �W)��
  ���   {Vk�Z��    �����  ���  ������o=    ������v  �<�   O���8
�   �a;  @^J
  �F|�    �(���  ��  4�R    <oq   �	�  ��X   ����  pf�   ��MK���O    �A�  pX\p  ��DĪ���d    ����}��    -��  ��D��"�[�͈8���V��   `�GD���z  ���  �)�iD|;"�."� "~��8��rBw    x��_F�_G��Fĺ�,   �	� �S����͈����Z�q6#t   �/:�}���g  HC�  ���}�������������mH�    �9����������    �� �Su�ߊ��j:�#�   8U��w]�iD�QD�{�Y   ��[   ��O#�����O[�X���   �M�Z�=�����  ��   qvv�~��q�=    �*޿   Nì�    �δ�뺮�$    ��v  ��"p  8BBw    ��  �4	�  ���   �C#l  8mw  � t    ;a;   }�   x:��    dSk�n  ��;  ���0    �T   �n�z    ژ��]�5�   �S#l  �M\p  8q��    <_  ��  �X   `�?  ���   �Ǵd캮�$    a;   ��  ���    l��   �շ            "�           $!p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�  D�8��^\\�`�^����z    �x�Rb�\�r��q�Y   ���    ����uD|xuu��0gϞ=��gϞ}}��m=    pxj��^�c�Z���mDD��x�x,  ���   �����������ggg_[,qvv]׵    Hl��ooo���6j��H  �M	�  ��ާ�c>��b���l&v    ��xw����z  ��&p  x���R��1��b>��|>o=    �@)%V�U�V+Q;  �	�  6tq�u]����b����[�    �Q�5���ݵ�M�zK��a���������j����
  p��   [���r���r�0�b���b]׵    ؁)j���Xk}��v]�0�0Ӂ�_y�s������  �"p  ؑq���:��e�f�X,1����    p��q���^J��w��}�=M  p��   ;Vk�������bw     �RJ�V�X�VG��[`���^   lA]  �G�b}��b���b1}�    h������Z�&���a|�  `��   O����2��e���"���Z�    'g�ڧ/1�Z��S�>�C   { p  h`Ǹ����j��nt]��    <�q��˗QJ�������l}�{�  �#�;  @C�ֻ�i)��    ���w�q��}�0�l&�   x*�  Hb��8�w�]�   �ǹ�o���!�ap�  ��;  @B�obw    x�m����c6���  �  $'v   ��{l�~?j��  ���  ��LK:�;    ��Q{D�|>��L2  ����   ���    ��m��qcǨ���  �  ���   p��O�SJ�q�4   �&p  8"bw    ��6a�t�  ��#p  8R��}��   H�Q{)�.l��w  �E�  pJ)�;    �ls���r�  �q�  ����B�;    �l�O��E�   �I�  p��e����   طm��)j��w  8,w  �7-����   �3�D��Q�  pB�   |��i�颻�   �M=6j���K��;   �E�  ������   �U���^k����Z;  �i�[   �ċ������X5�%��s�ӏ%#    ��oG���Zc�^���m���zw   "\p  �����W?��]��nD|��P�L��߾�]u   8A�\k/��]k  ��	�  ��2"�3��~�z��J)1��   ��ZcǍo�ڧ�$   x�;   ;1]��   ��\[/�܅�   �Pw   vJ�   p<6ۧ凜GE�    p  `/,0   �c�u�q�q�	  �5�;       ��RJ�Rb�֣   pD�       ���Rb�^��  ��;       �F��X�ױ^����z   ���       ��Zk����:J)��  ���      �;7771�c�1   8Q}�       �<��y�   8aw       �N��qvv�z   N��       ��ab�X�  �$p       �`6��|>o=   'F�       |��|�٬�   ��;       �F��<�^^   ���(       �F]���ٙ�  �'�O       ୦Ƚ�֣   p��       �W�"w   �'�;       � }��|>o=   GL�       <X��1��Z�  ���       �!�ah=   GH�       ll6���  �9�;       �(�0D�K   �e       ��u]�f�躮�(   	�;       �h]��|>�  �w       `+�%w   ؖ�       �Z��"w   �&p��ػ� I�������<�=?�eYw�]�vY@�B���P1�4���%��;�R1��\�n��RIʨ�YI!�ԅ���Quw�ǲ��5��V���P�C`vw�{�y��w�fv��y��׫�k~�|f�Z��ϻ?      ����  �-�       ��iHӴ�1   �)�;       0PY��$�$   �yN�       ��5�;   ��$	       E�e!�X�   Ԉ�       �ch4"w   6L�       M�1dYV�   Ԅ�       �$IB��({   j@�       ]�$6�  ��       �H�i�4-{   *L�       �L�e!I�
   �Ή       �F�!r  `UN�       ��eYb�e�  @��      ���1�F�!r  �4w       �"w   V�       ��1�,��  ���       �J�D�  @A�       T@��!MӲ�   �dw       ��,I"e   �dN�       @e4�;  �s"       *%˲c,{   J p       *%��,+{   J p       *'I��l6mr  �0w       ��b�!MӲ�   `��       @e�i*r  � w       �Ҳ,�  L�;       PyY��$�9   �;'?       ����  `�9�       ��eY�1�=   C"p  ���7    �D1ƐeY�c   0$w  �
�   �%I�ͦ��   Ɛ�  �f��y��=    �*��4-{   L�  P3EQ�=    TB��"w  �1#p  ���   �tY���  ƈ�  �&ln   ��eY�D  0��   j �s�;    ���h�c�c   �Ew  ���   ��4�M�;  @�	�  *��v    ؜F�Q�   l��       1��h4lr  �)�;       0V�$	i��=   g@�       ��4MC�ee�  �&9�  �(����sυ4M�oY�y�d    �4MC��!��G  `��   %�]`�t:���=���    6.����vO��yZ�VHOr  Pw  �
�   ��֊�W�n�C���  Ԁ�  �&֋޳,[�E�    ���}c��}iii͘}5EQ�v�Z����   *N�  PckE�����   �:)�ⴭ웍���s{���_  P]w  �1��yh�ۧ�O�   @+f_M�1�CQ�  �0�;  �X��.�����K    ��(BQaiii�6̘=I��n   ԃ�  ��z��{�B{:��S2�������w�    8Sy�/oe�mh���5H���?j��  ���   �۶ޓ��r��۪��Y�����[�   ���  0(w  �Z��F��.�G�i�n�{   Pbv   �I�  0&F��y�<?-z߶m[h4��߅F   ��ѻO�w��s�=7��Ӌ���   �M�  0�֊��<_~}P��W�Y+cw$   ��?f����[�2dO�d .   �'p  �01Ɛ��i�������j����w   ��x��}P��   l��  �U/*�Gｍ�[%z   (O�b�Q��=�    �G�  ��������2�w@   6o1{o�ʠ   �B�  �����{J{0u�T�   �q���C��<�C��r   C#p  ���?�t��"��   `pF���W����p�   4�;   �24�   ����>ʊ�  `��   �z���/�����  �*�f�����:   T��  �R�oZ�7��d��r   �U����   ԑ�  �JYmۺ@   `}bv   ƅ�  ���   |_�ދ�  `\�  �������.�   �?f��~   ƙ�  ���r�{�Q�   Ԋ�   �   ���ѻ�   @U��m�]   @!){    �  �*�2��    �;   B�   TY�$!I\�   �c   ƞ�   ��,�B���1   �Tw   ƞ�   ��cHӴ�1   �Tw   �Z��e�    �ai���  �D�      @�dYV�   P�;   c��v   ���$	I�r>   �ɉ  ��TE�#    ��4M�   J!p      ��I�D�  �D�  0v����   ��,��   FN�  �X�   �D�  ���      @E�ib�e�   ##p  `���   ��F�Q�   02w   �F��e�    0p1Ɛ�i�c   �H�  6�   �,˲c,{   :�;   cA�   �;[�  �w   j/��G    �4MC���  �xs�  ��ln   &I�ee�    C%p  ���   �$�1��  �Xs�  ����   �$��  �q&p      ��1��  [w   j�(
�  ����i�1�=   ��  �Z�   ���h�=   ��:    IDAT��  ���   �ci��=   ��  ���   |��  �q#p  �V�</{   �ʈ1�,��   F�       5�$I�1�=   ��  �ڰ�   ��lq  `��  �q;   �ڒ$	I"   ���n  ���(�   ��lq  `�      `�E�   Ԟ�  �J+��w   �J�4��   Θ�       ƈ-�   ԙ�  �ʲ�   `�$	I"   ���h  �,q;   ��ɲ,��   6M�  @%��   �\��w   j�i  �J�   l�-�   ԑ�  �����    �B��e�    �"p  �Rln   �4MC�H   ��X   *E�   0XY��=   l��  ���   ^�1�iZ�   �!w   *�(
�;   ��dYb�e�   /J�        ˲�G   �%p  �t��   _�$!Id   T��+   ��   ��-�   T��  �R��   F'��4-{   X��  �R	�   F+M�c,{   X��  �҈�   F�w   �L�  @i�    �H�4$�d   ��qZ  �y��=   �D��  �*�  0r6�   �/I�;   �#p  `��    � p  �j�   ���   �:b�!˲��   �ew   F�(
�;   @Ťib�e�   !�;       L<[�  �
�;   #a{;   @u%I�DB   @��N  	q;   @�5��G    �;   �'n   ��4M�  �	'p  `��    ���i�1�=   L�  �P��   �#��,+{   &��  ���   �K�$!MӲ�   `B	�  �<��   �3��i�1�=   H�  �P��   P_1F[�  (��       x[�  (��  ��+��w   �1�eY�#   0a�   ��   `|$I�DZ   ��x�5   [��tB��!����=I�姲�1zZk   �
�ݧ�[^��v�~   �;   [������B����n�kz�{Q!Ƹj��v����>.�   &��g�������#���z�e�kb�
��F�2�   ���	  ��lf��06�m6����    [�b1z�۫�}���ۈ�������K   :�;   ��v7|AtX�������?��j�4M_��   @}��kXZZ
�Ng��+��0��N'4�ͲG  `�	�  �Ao���lI������>.�  �սXH����C�h��aaaa ��U���n��  �A�  �e�n��j�L.�   �ă��7oiiI�  �P	�  ز4MO���qx��Wې���   �9��c\�/�����[�}�}-   ��  ��[��V���΋�  ���Jh�b_;�Y  `��   ��0��6�o��   ��Ӌ�mC  ���  0�Χi�$	!��.T�X(��}{��r=   �qyv�����SSS�O�   k�  �l4�_����ne�.�  `��y�����  `��  �&lw  ��K�D�   c(){    `�\�  ��4-{   `��       �R���   ��i   j��v   ��$IB���1   ��  @��  ��lq  ���      @m	�  `�8�  @���   �K�$��   �;       ���i�#    "p  ���   ^(I\�  �q�   5��y�#   @%�C���1   ��      P{i��=   0 w   ���(�   *-I\�  �q��      @��E�   0��  �lp  ���i�#    [$p  ���  ����   ��t      ���  @�9�  @���   ��i�#    [ p  �
�  ���C���1   �3$p  �
�  ���C��   u�T   %n  �3��i�#    gH�      �X�1�c�c    g@�   e�;   ��$q9   �ȉ      ��#p  �zr�  �
��   �&I�c,{   `��       ��4M�   �$�;   TLQ6�  � $�K�   P7N�       ��c�1�=   �	w   ���  `p�4-{   `�   P!�v   �4Mmq  ��      0��   Pw   ��  `��4-{   `��   P�v   �  �>�   Pw   �cH��  ���      {i��=   �w   � ��  `�lp  �zp�  �
�  ����   �'p  ����  `4�   P}w       &B�1��   X��      ���$.�  @�9�  @Ɋ�({   �i��=   ��;   �(��G   ��c��   *̩      ��"p  ��rj  ��EQ�   0��   P]N�       L���   *ʉ   Jb�;   �G�   ���   %�  @��4-{   `w       &��   �G�   %��   ʗ$.�  @�8�  ����  ��$	1Ʋ�    ��  `��   P��  @�8�  ���  �Z�   P-N�       L�$IB���1   ���  ���   Փ�i�#    �#p      `�%�K�   PN�   0"��  @5�C���1   � p      ���i�#    A�   #Q��   PaI��9   T�:   ���   �-�(r  �
p:      �B��e�    O�   Cf{;   ԃ�   P>�s       ��;   ���   ��w   ��4M�   &ZV�    0�������{��-  0��<?���i/W���$Ib�Ν   P�;   ���+�"E��n!�n���y��<����t�2w[   l�z��<��χ�r��$���4MC�Q�B�$�gV   `�\)   �?T_�z/d�  �No��z�v�$!���I�,���i*p  ���  `H�-����EQ�������  &E/��\M/pϲ�|��q���s  `��   0$u���{��z��W��   L��9����9�����#|_I���   %�  �T)n��WF��u��{[�z�D���  ��w�����{���7���Ra��7��-�i���Ǘ��i*p  ��  ��z��j�֋�X�	��+C��ޮ��  0(�3�jz窞,˖��;G�������п�?�v������  �I#p  �
���ھ^����������e��M}   U�b��g�
!�F���^�w+[�ܻ����w�e�"���g*M�uL    ��   �`��
���1^_m�z�N  `m���ރ�����ίe����t��������޿�?�_��   FO�   ��y�v��/Wnaa���jVF�+7�WA��>  ���X��9��oZ��C������P}�~�   -�;   ȩS�B�o����-�EQ�.T%^  `u��7������\k#|�#�,�B��(e.   �Dw   �ކ�2�����   �_��w}0�z�{�v�Q�v�w   !�;   Ш��?�S�   �֌�p�g�ރ�������8�E��nH�t�6   �Bw *�رc�c�=v���7�ͳ��8��� �<?��>�`�cP3[��޿e�(
�����   �^�$��\�wV,�b����f���3L��������� `|��m��Ϯ|��}��~�ر� V�0P��rKs���/!:�s����l�Z�[��K����7��m�fs��j5�F�$Il4I�$1˲�$�iwL� (�׿�� pg3֊�W{*���   6�yrm���"�V��Wn���v��=�k��᷽�m�= ���`��n�)�y�<KKKE��E��ɋ�(�:�N��n�\\\�_XXxnqq�v����<���?���_j�����#���x`��	��!p`���ַ�?==}���ܫ�:�˷o�~�m�榧�ggff��V+i6�1�2q: c�V.�D��:   ��̹u9��o��a�1�,�o P	�{�ޣ!���٫}rQ���n��v���8q�}�������x���y������������g��'F�s PsNH ���n�|ǎ�۽{���s�eg�}���۷����6��fȲ̝�  kXo+ñ٧�  ���%  k�=H+˲�j�b!ݵk�t�nn�����N'����|����<���=����x�g���o�����?p�=�|���J�L��o������/���^�9�|ǎ��>��V�Պ6D     @��=� �ʋ1�f���f8묳{��}I�%!��!�[;�N���[���|�駟��SO=������?���|�c�����_z&��`��r�-ͽ{�^�o߾[v��y�K^��ܹsfjj*�8     �%p `4��h4z�����µ�N�W�򖷄g�}v�'�x��'���G}��=��C���?�){n �G�0f��7���/}����u�w�޳cǎF��I��=     0@1ƲG  ����[���0�pa����[o�5<��3�'�|�o|����G���{�}��y�;@��~��ssssw�߿�'w��uѮ]�ffff��  L[
 �I'p `Ҥifgg���ls߾}���ʃKKK��z�œO>9�������������#�ȳe��������>�o߾;����{��9�k׮�V��l     �@�  @Y���۷��۷�u���k���k���7�i�[������׿��?�����{+{V 6F�Pa��v��={��������ݻ��s�9'k4e�     T��  V�j�={�={�\|�W�����/�|���o|�_}�G����#��N�=' ��Tȱcǒ'�|�փ�����_�gϞ����� �J*���   J%p �����
�~���Ͽ��k������_��W�x��G?�կ~������e���	�Jv�m��ܿ�{8�������YgEwH     c� `  ؤ���p��^p�7��U���'~�'��{�_���������o��}��&����z׻�8p��_xᅯ9��f����	     �!�;  lM��a�Νq�Ν�>|�WN�<�+ox�����ǿ|�G~��{��j�3L�;���y��_|�ſ}�Eݽ{w3��     l�g� �����	��~�С���~�MozS��Gy�������*{>�I���;��'/����8x���ݻw�i��=  ��	  �K�  ÓeYػwos�޽׿�������׾���?~�W���.{>�q%p�w��ݯ<p��\t�EG�=�ܦ�     �;  �F���w^���{�ѣG?��?�㝿������?�o��O��+e�0N� ��w��.�胗]v�k���ZY�W     `��  0z����ػw��^{��?�c?v������K_��/����.{>��S`��n�!{�k_��/{���ܿ�ٍF��  `bEQ�   � p �r5��p������7��o|��:~������رcy��ԑ�`��뮛/��߻��/;묳�k<$�nw��� ���   P%1F��C�E�����1��#�4�$�mff&\~��/�����~ꩧ~����_����'�'�.{6�:�l�����/��?r�e��ynn��$I�#UVQ���<�C��]~�w�v��(���W��ｷ�
���o�=�
�/  �N��v�ԩ�裏�= ,�z-L�q��$IB�1�i��v����L��R�1�ڵ+y�k^s�ѣG?u�M7��җ�t��?��_���?�){>����u�u�]?z����C����-{����N���nXZZZ���     �謵�  6���p+�c�4M�_6���'u�d�����袋~��o��+_�ʗz衷�ٟ��˞��� +�r�-�Ç��+����{�NM�S1��N���������  �fB     ���R�Ng��佭�F�[/�w1ưcǎx��^q��W�G~�G�������{��~��� �F��=o}�[�����?����_�cǎ�_u�����������  �L�  p:� ��^�n�_�$I���f���2��3ql6���K/=�K.��o��?�����_~�_������e�P���?�&�u�]?z���/�䒗�Z����v�:�Nh�ۡ�n���E!;     �	�;  u��yX\\�����?I��l6C��
�fs�6.b�ann.�馛~��k�}굯}�?|�_���{��\ٳ�I�L�cǎ��W\�����73NOs��t��_\\�vۆK  Ɗ�o  N'p `\�y������z�ާ�����F�Q�[c۶m�x�+>|���^{�?�ӟ�W��{�_�=@��D9v�X�h4>t�ȑ_���k���ޣW���<��     ��_�  ��Xm�{����j�V�������V���⊹�.������?���|�7>����� FI�L�;�cۅ^xߕW^y�Ν;k��=���n�éS���v�+ �$~�  X]�љ	 ����v�ɓ'�ɓ'��׋�{�$IJ�p�,��9x����u����}�s�����B��?0���X��;�]|���9r��۷o���2�������ɓ�ԩS��n�=     PAw  8]o����>B�n�>==���k��=I�p�������ޣG������S���/<��Ke�0,w`,}/l�/G�yS���ކ�ޖvwF     /�.q  ����;�	I�����0==���B��,{��$IسgO��7��G���믿��O~�Bw`,	܁�����}ǕW^�?>|C]���-������=  T��  �N�  ��y8y�d8y�d!�F����}zz�ҿ_�Þ={��o���|�+��믿����x�������!p��7ܐ�|���������:��KKK�ԩS�ĉ�� �&���  ��*8  Pu�N't:���sυ$I���t���	���!MӲ�[U�1���e7�|󻮾��w^p�|����+e�0w�֎;�LMM}�������;w�U��vii)�<y2�8q",..�r     ����5  ��<�É''B�1�Z�0;;fffB�U/��1���;/{�[����]w�/��_�կ�����`�slE���ؠ������W����{����[��t��m��e�  �灢   ��1z�+  ��(���BXXXO?�th�Zaff&���V.vO�$�߿���?������3��������/{.�3Q�a6��}�[�=��}���VqI�����a~~^�  $�      ʲ2v���
���avv6�iZ�x��4�\r�����#G�<��O~���w�Ce��w�6�����ȑ#����Kϯ�/�!|7j?y�d�������     `�lp ��Y�o۶-��̄$I�-�B�e᪫�:�e/{��~�~�o?�����O|≲��?{�%WY������[wWW�;�+� 	I�FBB�	���u�qft�Pg�<,=gd����AA�`~Q��Q���0��8#���0DZ��-hȥ�����뮽�*;���]]��k��4!��'��v��ٟ����Լ}�C�7n�񩧞zj8�vw�<�S6�U"�P2�d�        TU-�|   4:��N��N�e�Z[[���D��5IRKK��nݺaÆ�[�l������{�ǩv� �h��i����z�Yg}(��̌�mۚ����̌��|��   $�/�    IDAT4�   ��p   ���<%�I%�I�AE�QE�QՏj�b1�mo{��7n|ײe������o�v� ��T��	 Gp�7�sӦM��t�Җj�E���g"�P&��vw         ^��;   P;l����&''��ҢX,���֪��0-[�,x�UW}yÆ�x���/��;��j� ���)��GWnܸ��O>y�eY���Q<W"���3   PM�aP�    ���;   P�����������ŪZ�ݲ,�_�����ϮY��?�zꩋ��t�: �A�@�����M�6���+=�S:�V"�P:�&@   ���   ���   �-��kzzZ�x\�����b�D"U�O[[�.��-�ׯ�/[��l߾���u f!��ꮻ�K�9�{�/_�R�~x��D"�x<.۶��        ����   P�<�S2�T2�T0T,S{{{��.^�8p�UW}y����������wU� ��T͇>���3�8㱍7�Q�-w�����fff�8N��   ���    ��p   �m���Ԕ�Ѩ:::dYւ�ò,mذaѪU�^9���馛�+���� ��*>��Oݰy��:;;�j�!��hzzZ�t��^             U�8�������F��
������e�]v��'���|��o~����� ���XP���{�<��_�|��k���P��٬����J��r|    sǢT    (�a��   �y�<O�DB�DB������T8^�>����?>��~��u���䡇zˣ�>�_�N hj�,�[n��g�}���X�*3�333���V.����   �&��+۶���e�Z[[��%   4�L&#�ueY���`����   �#�J)�J)����S---z�H$�7����Y�&�v��˿����xA; �ipPq���m۶m�I'��l�'U=�S2���Ԕl�^�c   @-p]W��C���"   T��8rGҡ
���{ �i�U�]}"�   4�L&���a�B!uvv���m��m�V�^Y�t�֮]��]w�u��� A, E�@E}�ӟ��֭[o�F�:��y^�b;�v    ���<���b��   j�����C!�`0X��.�   иr��<X��{8ֹ�{Ί+�<�ȥ����;8��C�@E�����<������`�BN���SSS���v\    ���a�|>/��Jz��j�   �B;����y��r��r�T��nY����}   ��{WW�Z[[丆ah�ʕ�?��?~tٲe�p�(��� 0��������s�9玮�.k���y�R��&''��   4�R����u]���b��ܠ:�-   �i�����w(2C�@��;~�0��  �&���422�`0��������ҢK.�䭫W��?��#[��o<� �4��ͻ���Л���_�z�r"9�Jibb�`;   ���y^1�n۶/A�4}�   P�³�rlz�W�?�d22M�vM�K�   h.�m�����D"���R$��1��	'�x�������[�g�
�ip��?��??�.x|``��wG�G&���Ą���B    D!��8N�J�|�!�0d���(   �˲�y�<�+�NTN��B1�0����=p�h�/   �C2�������ڪ��n������ݸ�+�Ǌ+�}�}�m��~0Y�hx����>����s�9��B����8���T2�\��   ��f	a�����y��av鍫��   �6{1fA!��8NY�ƞ�)��)��IR��{!T���F��   8�T*�t:���6uwwwЪ˲t�g.;��FW�Z���o���= ��G�@ٮ����駟��)���b!&J]���Ԕ��x�\    4.�u��狡�����������<�/   Xp���>Բ�b(�����yF�8Nqg$�0�7��   x�����R)������sN�����g]}�������'?���+z0 ��;����_���۶m�Nwww�g}=�S<����   �-��v۶}Y�;�B{9B/   ��@zA!�^�BQ����LF�i��@�⁏���>   ��u5==���uww�����c�p8�K/���+V�}衇N�ַ�5R��hX���m��v��͛��P(T�c�R)���+��W�X    �7�qd۶���/�����|�<�
�   �;�i�4M��=��
�sUx�mے�w��b��cv�   P�8�FGG����ݭH$R�c���SN9�w���޻}���+v0 ��;�����w�yϝr�)k*=�k۶��ǕN�+z    �����������y��f�T�*���  �1��c��E�����8e��z��\.�\.'I����   ��e�Y)����[�eU�X===����ouuu]��O~��@�!��$����9������̭�y������4!    5��b�ݶm_�1���
��FEG   TK%�C-�*������r8�#�q$��

�r�^.��   ��̌R��:;;��*�{U8֥�^zՒ%Kλ���O���ש�@C!���>���޲e˖���4��L&511�|>_��    @�
�v�qd�v1�2�+NVz�,   �V,T��4M���@  ���y^1�^N�����t:-�0jꞾ��   �6�����	��̨��G�ʇ���SO=uqoo�HWW׶;��9��A��Q}�+_y��3ϼ��H���&&&�L&+v    ��������y�ivu�Z��X�1   �f/.��Ϯ�^ν��y��r��r�T�oYV���   �*��ihhH�hT==={~�lٲ�������������~���@C ���>��w�z�/�񽕜 ��㚜�,{[P    ������P�|�+��� M�0��;   ���CÐeY�P�k����G�q�;=��@ pX�}!p   0W333J�����V4��1�Ѩ��w����q���_��@�#��u>�O�{�������b׈l6����bE    ���v۶}	�̮�^롒Z   ��H/�]ݽ�������LF�i��@��`k},   �69����Q%�I���6N�K Л����������u?���P��8�-���۶m�L$�H���ijjJSSSi    ��hw�X�}�fWh��	w   T��y5�l��L�T ��y���>W��ٶ-��8"�~����   �m�TJ�LF]]]��b��o��N=�ԁ�����˗�~�w���  �w E;v����g�}U����d2+N�   �����f����n�f�T񪋕D�   (��E�����8e�1<�S.�+�v[��nYVE�    0W��j||\333���S0��˗/����}����On�����  �w ����e˖nܸ��JL�z����IMO��   ��Ắ��|1�^Nu��
a��Z�  P�P��X,�*��_[ݽ��l�q�;L��@ pX��ap�   `޲٬��߯��.utt��~gg�q�UW����q��7�|�� Pw�M���x�)���+WvV��l6���Q��   �(������>_�+��{��h�   ���H/(��]p�y�lۖm��d22M�v%/�%�   �/��ibbB�TJ}}}�����D�����c���o�����8��C�hb���6\xᅃ===�_<���Ԕ����n   @�8Vcv�=���;�1�B{��m���   ��*��i�2MS�@@�置��\^W((d���`1��F�e#��    �#��h߾}���Q{{��m]|���vuu��;�RUhR܁&��O~�/�������}����rU.��i    M�u]��yٶ�[�}v��fE�   ��ًi
aw�q��x��\.W|S��nY�a�w��   T��yS*�Roo�,��m�4�iӦձXl쮻�:����q u��;Є>����m۶}1������&''�    `^Ð�y�@�m۾Uhm���1~   �eY�P�����՞�8����@ P�   @��R)�߿_���jmm���u���>������Z�����/��8��ǌ�d>���o?��s?�����8U:���]    �)�N��+��
�T.<2�   ����H�ݟ����;��<�+.6C�H��.   @��8Q4Uoo���+V���O���X,v�W��՟��0��G�h"�7��M�.�{�8�Nktt��"    �Z�/fWh'0S�r3   �|y��=��v�)��Aw�q�@���   Pi333��r���S(�ݾ�>�=�y���p��v���O�5��p��W���?�3��=�999���i*�   �U�c�������7   T����!˲dY����못�2v"�   `��r98p@��݊�b�����n��]��ǖ�����z�g}k@�"�4���x��O>��6���FFF����l    ��P�pv��Âe   ,4v*�a
~��wvu�7z_��   ��<�����2�����|[p��Ң�/���H$���o�Q 5��;�����i׺u�N��T*���Q&�   T�� ��
�T�a   T���0MS�i*���Ux���   P�dR�\N���
�B��
�������P(�w���ȗF�$J��;������~w��p���<H�   @E��AY�%˲�Tc<   ,$וQ��**���E�P��   ���m[P"���`0��.��_����[� jw�}�;߱����q�7�W���hhhHSSSL<   �8�   @��9��),   �j�<Occc�m<hY��=��+w���/�9܁s�7FZZZ&�.]��W��LF���W&��I        Ф�   @�I$R>���=˲�y��K�o���/�)܁�����3�_�xq̯6�񸆇��8�_M    j�a�        @�e�Y8p@�tڗ�L�Ԗ-[�۾}�/|i@� �4��|�#��;１���V?�+l3>>N�    ����   ���    м���𰦧�}i�4Mmݺuӎ;��A 5��;� �����m{����~��8�����H$�h             ����	����R|�0�s�9�o�N�h܁:w���]x�{zzz�~�W�&����    ���Q�.   �ɰs,    @�������8μ�2C[�n]��/|��>t@�p�؍7����K_�����^*���А����    ����   ��,    �LF���W.��w[�ah۶m>����܇��"�@��������O?}xѢE?ڋ��:x� US    �	1  �Bb�%    `6�q444�T*5�L��y���[o��g>t@�p���>���s�=wxɒ%-�m��<���j||�@    4!�g       �js]W###����w[�i�.�v�M7=�C� Tw�Μ����[�-^��u�m�����a�����5              �611����y�cY�.�䒷�p���C� ,0�@����?�wٲe��mǶm8p@�LƏn    ����   ��    �&�kddD��ͫ�@ ��.���_��>u�!�ԑ��|eժU�m'��ihhH�m��-    @���1   0,�    K*���АǙW;�`P�]vه��/��&��`p��w���֭[5�v��/?�    ��
�   XH�    J��f})�
�t�e�}����ϯ��k *��;P����7�9�	ߙ����P             P�l���Аr�ܼډD"��+������O]PA܁�cǎ��v�iη�x<���1��    ��+�u]vP ��9�Üz�P�    0��hhhH�Lf^����+���k���S� Tw��}�_��͛7`�����g"    ��8�R������l��  ʔN��ǕJ�X�3�W     ��u]+�Nϫ�X,f\y�O����^�S� T@�� pd���g�y��g�4�ebbB���>�
    Ј�öm�r9ٶ]��B�W�� P_\�-�#�r9�r9�A�B!��*�����˽    �,��iddD����F�e��h�"�=�y�K�����z�/Tpj�M7�t�֭[�	�B�jgtt�p;     �y�l�V<W2�<,�^����3  0G��n۶�ɤ��r��    ���466�D"1�vV�\�򶷽���jL��\����l�򋖖��˗x���jf��e     T��y�d2J$J&�r]��.w  �ϑ���(�J)�H(��t/�    �Q�Ϸ���������/�ڧn�Q�� �{7�x�y�駿���a��F!ܞJ���Ps�Q&��$e����d2)I�,K�HD��D�����V��   ���<�Y%r�8)�=�m[---�  ������;�LF�lV�`P�HD�Im�cq��]    �N:���r]��	��rŬDkk�ÐeYŹ�P(�`0X�>abbB�穳���66o�|��7�|�7�p��]0O܁r�	'��dɒ�r_O����<MMMiddD�x\�D��{"����L�����	�F�jooW{{{��X,V����vuuu���_�hԇ-   �ze��a���4M�B!9�#۶�.�7  ��8r]W�e��c��=�S.�S.�S0$D   ���i���jll�uy�#�*u>�XZ[[�C��K��XL}}}���e�]�Xp���r]W���e��0]x�����������>����L܁�կ~�{k׮]U��=���Ȉ�鴟�|�H$4<<���Q<xP,~=::�ۀl.������455U��oiiQ������קE����O���P8�p�  ��1�
�G�y�l�V&�)���th7�P(�@  �0��x�q� P'lۖaşݖeC良ֶmY��p8�`0(�0*�e    5"��kxx��\���DU��J��J�4<<|̿kY�zzz�H�^�h��������LOOKR�!�`0��.��T*���o��!?��<܁�cǎO�~���W���<O����d2~v�3�qt���۷O{���+���}��idd��]��t:�={�hϞ=G��]]]Z�z��/_�e˖i���Z�t)   ���n�
k���`0�`0�@���B�#۶��
 @�p�u�t˲dY�\ו�ǼwrG�T���K8&��p�	  �F199��{�j߾}ڽ{w1+Q�"~r��?���V�X�B˖-���˵z�j�\�R�Hd�{
nzzZ�a�����U�]v�ccck������; sE���[o��7m�tC�!�B�v��Xh�mk���z�����V����8 �q�ݵ����������|�r�\�R�V�Һu�|�rd  �&y�������(��ʶ풂W�a(*
���V˲d�f�?� �Yx��|>��?�MӔi�Ő��ù��L&�l6�`0�H$��E1�  ��^��/��W_}U{��Q2��v��"�J������?_�3�0��߯�+W��Ӊ'��O<Q---U�)���Ԕ�PgggY����5�����^z饮��A&��*"�T�_��_�mڴ��ʭ��y�<�t:�sπכ���K/��W^yE/���~���8�l6��_~Y/��r��"��V�\�u��i�ڵ:餓���V�^   j�`�m���r%�q
�X��`I�eY�m[��6}� �Z�8�<�;�����7MS������y�b
�uwV  ��9��={������ݻ�k�.���U�[5�P�sddD���/$/-Y�D�W��I'���k�j���U�)����$�r_�zu�5�\�����:?�`n�Ut��g��Ŭr^[��R)��H:���駟����^�����:�    IDATP���2��a+�-��ʕ+�v�Z�_�^�ׯW8�r/  Ќ�-h�y�l�V&�9f�Ղ@ �`0�@ 0��*ȶmٶ��>  5.�����a2C�i��ǪP^�/�,K�p��Es    *#������3�<S��r�jw��}��i߾}z��$I���Z�n�N:�$�v�iZ�hQ�{�F5ߐ�Yg���S��Է>�O\�g� ���;P%�����ҥKc弖p;*�u]��w��3�<���A���5�Ul p�ǘi���CkE,˒a�UMr�X)<d���h���ڽ{�x�Y��N8Ag�q�6lؠU�V�p   ���+�u�b��R���`�l/Ga����	� P��p���3�u]��{��+�q�J���Ä�a�  �255�_���ԯ�����&�8���s�ҡy��׵������	=��z�'$I�-����a��z�jii�r�H&''e��b��G���E]t���ď�o�~g���U�cǎ�9餓֗�Z��4::Z�7֨���ڵk��|�I*�LV�?�@@�HD�pX�H�"�&)�Z�kt�m+����m[�\N�lV�LF�L�8�[(��+��u�]���Ԇt�gj�ƍjmm]��   �9�62�q��fK��d����B��LӜױM�,Vu  ��P4�)W�g��yŰ�Ѹ��L&�l6�`0�H$2���Z�l;  �68���^zI���z�g������s��a(���������_�e)
)�{|0;1;+���d۶��2�LU�֏��hddD?�����N:�b�}����4���q�����9�6
��.�cbb����7���p܁v�m�]��7���-w�v||��!dԷ��	���?�Ν;�R�ݲ,������M����D"�P{����0���X�)>\J��J�Ӛ��Q2�,���|LMM���c�=�`0�6h���ڴi+�  �ض�l6[��U˲��?�W�@@�\Η�  ��BuC��
�M�,)��y^q��`0X�    (��z������LO>�dU�I������Mmmm�|D$Q(Z�>�cf<�+�f�J�RJ&�J&��m����m[�<�y��u�]Z�l�6oެ-[�h�ҥ?>��ؘL�T[[ۜ_���a\v�e�ܳgOǣ�>��U2�&G�X@7�xc��N�����Ą��ϽB3H$�կ~��;wꩧ�Z�`�$��aE�Q���)���T�ǲ��`�2�Lq0�J��Ǖ�f+�۶588���A��   �]#Up/��2�L���Q�
�B�mp �F����TN/�-�*ݏu�R��hYV��c=ͫ   �⺮^|�E�ܹS�?������ײ,E��bF���U�h�����PKK���m+�LjffF�TJ�D����ۧ{�G��sO1�u�V-Y����Ec�ajmm��kW�\�z�W>��+�5 o�~~���{�]�bEo9������Ą�]BK$ڹs��x�	�ڵkA�*---���P,S,k��u.���̌�񸦧��H$*�އ�a�q�:�st��S�	 |t��]w�uU�C�� T�i�
�Bu�v]�X��ԅ��ꨕ�w{��D"�`0XV���������5{?+#ׂF:��vn�Q��W�u�ȏ�ca.o!>ץ�
�j�p��?��t��k x��7��k��v7 �ny��g�}VO<�~��_.H��P(����b>���������q����x\��T���W�.Vv������8�����"�Ȝ_�8����>��O�]p��S����������O��r^�H$466�w�Ѐ<��/�����gz�ǔ��*z���6uuu���K����@�O��*�HhrrR�����������ڴy�f��-o�ʕ++z, h�4�z�;��l6[��4M��%�I���X,6���b �k�@t9-D�H���M9j��J��t��<z����i��,x�W���0�AE"���� � �G� �399����g����V�X�`P������TGG���pE�W�<���̌���599����4C�ׯ׶m۴y�f�B����4M-Y���⑩TJw�u�y_����@� �Fs�V��n{���{g9��TJ###���Ԕ}�Q=����~�,K���VOO��2ض]�MLLTt��իu��k�֭e�> p�\�P8����m��f����%�}˲���d2��r�F��
P�b �k�@t9-D�H���M9j��J��t��<ڶ�d2Y���)9�.��`��vt$� �G� JW�����뗿�eE+�G��bѿ��hF������W&��ر
� ��ַjŊ;C ��ŋ˚ڿ�}�w�|��߯�V@��.Pa7�|��m۶�kii��lm6����PEW3�~-Ԡ-���W���M��V%V/���ittT�l�"�iiiі-[t��k���9 4*� �I��=�S.�S&�)y����m[�tZ�Hd^�Pk1���5R ���n���h��x}%�^��~S����|M|��K��1MS�pX�P�.>�����������������Cill�"�0MS]]]���SWWW͍�]*���Ą<�d2Y����{�T��
�BZ�xqY��'�|r��o���
t�,�?�Թ�}�{�˗/���l����PEW��>��i=��#z��4::Z�c��b�����.�4�T*���1���Tl��	'������zӛ��C$ (w �&��D��H\�U6�U.�+9�
�k���y�������h���b �k�@t9-D�H���M9j��J��t��<��qI��ϴ�yŰ{)L�T(R(���� �z���=��s�����SOU�@�a���Poo����jn\ب2��&&&466����#���/�[��VuuuU��o�HDs�s]W�����n��V�k D�����ۿ����:�s}��8�mە����Ԕ~�����J�@ ���~���Q�����b�=����~__�.��]r�%jmm��} h�4�Z���ye�ْ�Ȧi*(��&�L�u�ymi\�L�����h�u#��F;7���+�����躮���@M~�t7C�`P�H��<�S6���� ���; ��<��{��K/�T�c*������X�٤R)�������)t�9��+�Њ+|o�-����w���T*������Y���d��4=f��
��g?{����os�Pw]W����f�����~�;�w�}������T��bZ�x�����⡂�yrG��ߏI:l�����4��˲dF�>�z-��466������Znii�\��/�\===�� ���;�f⺮Z[[k"��y^1�^�O˲
�j�^?��(��)�����(]#���h!�F:��vn�Q��W��1��)�J)��+���V�,,�������rM���"� ���i���?�}�ݧ��1���Z�h�����{���8N1#�y�a���bX����0^����gM������hE*��[�NW\q��8��%(���,����={�_��c�>����+��fj�q�7��u�Y�-g2}||�p;$IO=����������@ P��J���Be�B����q�������P�Ѳ,��P(�`0�p8�P(T�Նa���O}}}J����Ȉr��/��i=���я~��[����/����}i   �+�ue۶2�L�/��`����"*���d� �fe�v݄=
�R���U�4���qT"�  ��7>>���_�<�����wuui�����P��y�\D.�S.��m���w�u�_��P����#�=g��ѡ���Y�F��АR��o�?���z���r�J���oז-[�fn�355%˲�����+V�\q���裏��B]�Z�b�����o׬Y�r������H�fԗ�^��ַ�k�.�ێF�Z�lYY[����<�r9��ie2e2�b��ρ��
� C��"��"��ZZZ���>���i���J$��m��>�l]u�UZ�d��m@=��;�fR�
���z*ܣ��5��<%	Y������� _���w9�Jx#��F;7���+�K7������aU�I�bc��ALӬ�}T��	 �pTpЬ����>=���y+В%K�}m�T�|���H���9P۶�ҟR��`���hmmU$�ڼA<׾}�4>>�{�}}}���+u�2�nr�ah``@�HdN�����{>|�m�}�B]�Vs�V�cǎO�s�97���nffF��������?�o������ݭe˖������߈�yJ��J�R�߳٬�ث�0�bؽ𫭭mAu����W_}�/^�k� PO�h&�㨭�mA�]�|����a+�u�����iٶ��������D�)]�FQ7��l�sS�Z��p/]��G�u����3�8N��a+�=Vح p8� �M"�����}=����f����D�d�,�=��iff�fO�����0����2�htA��tZ��Ȉ�㊥K���x��m�V�cC��4M-Y�D�`pN����t���/<����� q5|t�m�-?������9}�2�����ٚ�I��⋺��{588�k��i���WK�.U4���#q]W�dR�TJ333J&�f/U!���ڪ��6�����Ʒ�tZCCC��}�,K[�l���iѢE�� ���;�f�Pw����R��!�4��C�4�Vu��lV�lVmmme�j1���5R ���n���h��x}%�^�r?��lV�tzA��J��{����������m7�1 w �"�N롇����=�R)_�^��=�S&�9,#�w�z���֦��6E�����������}�W�X�w��]:�쳛~��Y�A-^�x�sO?���|�+*�-�)q|t����X��{.����ڿ?�M�W^ѷ��m��W��]�4�x�b-_���$<�S"�P</�BƑ��aE�Q���+�U���m�ڿ��ו`0��.�H�|�;����[� P��h&�몥��b�>����R�V�P�k$�{�=��+�J)�������Z �k�@t9-D�H���M9j��J��t�~��dC}�g�<�v/E�+
U�z�wuN h�4�t:������|�wtt�㎫����tZ�DB���J���|�@0T[[�b��b�XE�ٞ����ڻwoɻ������UW]��7��.�CKK����uu������n��
uh:�=[��+_��76m�t�\^㺮����vg�J$������?�u�c��-Z��˗W,������le(Tx/����*r�J���.��r���h��V �F�h&�
����l6�\.7�`��Bf�p�<O3332C�Xlί�� &Jר!�R5Z����g���r�����{���<����n1���<y�'�qJ���i*
)
���p�##��Qy��������7����q_ێF�:����=�:�%+����V<�=@�,��p1�F+2��y�����ꫯ���ڰa�����i�

s7���Nuuu��5�dһ���O��{^�P����ܳՀO>��ϝ�u�֧B�М^w��A%��
�
��q=��C��N�}k�0-Z�H+V��H�#�JijjJSSS,ƨ�`0���uvv������\.��޽{544Tr��===���u�y���& �"� ��뺊D"�-d����f�%?�1C�a�L����th��������(]#���h!�F:��vn�Q��W�+����533�@ �4������b����"��o߇����hD/�����N��⋾�[�`{>���Ԕ&''�J�|}ƎCϼb��:;;��|�9��h߾}���kY�.���������}k����΅+_xᅉ����=��Tc����|�#/vtt�����Ԕ��x�����O��[o��?��Mt__�N>�d-Z��ׇo�TJ���ڻwoq!F��}07��*�JibbB��r�,Ks]0�F,�Rww�������}[T�N���_�R�v��ʕ+����K� Pk��~��W��i6M�@�Y�5����y���J�R�f�%�&d�f�b{��)�0j.�8W�������c�\׭�����5����s2�v>�ܔ����اZU��1��5�B�R�J��;��l6�|>_�bģ�m��5 p$zӛ�T�n �/&&&�o|Cw�y��U�#��N8��Y�F---�����511QFS��r<�S&���Ԕ��Ɣ�d�;H�1N0MSZ�d��C����y�^y�=��#
�BZ�z5c�&�J���mOOO�q���'?������g����}�k�'�i�!�Nkll�R]Bٿ����/��������ѨN:�$-]�ԷPG.�����o�>B�U2;�>>>.۶
�|9ǁ@@������.���0::��~X���Z�n�"��/�@� ��٘�Y����y�f�J����r%U6�j��u������cil�V*�*~�ՊFD����m�|6ҹ)G�]_]���̌�C�К��K9��l6�p��R�Q�K:���뺲m���g�ߓ��< �p�4�l6���__���{�n�ڵ,K�w�֭[7�J�o��<MNNj���ڿ���8;�/�B�}rrRccc�f��4MS���Z�h�r��R��=>��y�駵s�N-Z�H�/��]Զt:�h4:�=g�r�~��g'*�=��1���-�ܲ������\n�l�ցJ�b����d��o}K?��}=��`P�w�|y�y����5>>���U����E��������a����v�����mmm��?�]t�E<��08�뮻��}�KEc ���
��� �u]e�ْC�|	���pxN�դBh1���u�|�!���y���dq5˲jj��f��Z��5Ԙ���g���r���5�N�nL�T[[[�|�U�\?���)��nv��<�]��
������i�o 8��7��k��v7 �l�����׿�k�vI���תU�|�=����P[��zzz�����=�k�����X��}�ٺ�k��	D"�9/hصk���ٟ�W�K@S`&���~��/wvv�\���<s����~�i�r�-���]r��XL�Բe�t��'+���ac6���Ȉ^}�UMLL�����y��q���)��)*Ϋ���V-^�X�a(�H��j۶���j�ڵs� @-��;�fR��Y�C�|>�t:�t:]��O�aȲ,_M�R��q9�3�-xk��p-�m�u;�y�������R�l�to�h糑�M9j��꺮��t�=ϛw��F7��c>�W.������������{�nɯ��; �ԫ��i}��_�]w�u�f�:::t��'kɒ%�^�뺮��ǵw�^)�LR���9��D"���Qe2Y�5�b'�pX
��J$���}���'?��B���?�x�:�0��DJ�	����m����?��OX����;P��}�k_?��ϙ�k���|��GmI&����;��o~ӷ퍤C�����@}}}����ڻw�8�T*Š��x��t:���qMOO˲,E"���/�Pgg�����J���d|���ؘy�9���k��̃a (w ��h��B�)�L*�͖4�(TD�;8�(��{Z��Z
`�
�u��#-�u]׷J_��h��r4ҽM���F:7娥�k&�9b��|>/۶kj�N����Ѷ�څ�O����a�0�c�pG�l����h�)w 82� ��Ν;u�-�襗^��@ �5k�h͚5����r֞={4==M1�:��d499���I�����y�#�Ѩ���}��n۶�~�i=��sZ�vmM�$	e�Y�B��R�����M�e}����JT�{@Cb�(×���e��v�?Z�U�]��̌���*�-T�Ν;u��7�7���omZ��U�V��㏟����<MNNjϞ=�Z{���󚞞��Ą<�Skkk��`0�E����USSS�,|p]W�v����j͚5���w� P�4�0^79�y��٬��r�\I��B핺�5J��0��m.�Z
`�۶�J������5m�@t9�ަ��g#��r�����Р��s��f    IDAT����X(�P�V�ޅ����뺲m��ߟ�m��pPOFGG�}�v����������r�)���W;�tZCCCڻw��ɤ/�����)�z������R�be�4��ӣ��.%	ٶ�K��������B�.�N+��|~��������߶W�k@C"���k�����+���r9���T�K����Q�رC������f}k���K��r�����~@�8���ƴg�MNN��A�����_rmmmZ�h�l�V2��������O�t:�u��5D	@s!���̮$�8�2������|���B���׮F
�۶-����n�0��XUۥC
�w��j��{����H�6�v>�ܔ�V���J�ҡ��ot�������y�<O�L��V	
!������sf��Tp�##���������۴�~���B:��r��y����ꫯjhhH�tڷ��v����)��̩��k��a-^�Xҡ�?8��]�v�W����?�xuuu��.jG� P4-yl�������;�������w`����/d���T���<O���G�"���s�N}�3�ѫ���[��@@'�x�V�ZUvX�q��6[�xܗjܨ}�r�m�������eY���U4�����yz�����\k׮e��p�l
כB������ʞ�k���th�8���`��_�0�)��)�L����eYjmmU(���_sy�+����h�{�F;��tn�Q�W�u���=F������Q����yq���pHE�a˖û�u�N��Ev��. X��7�&�^�����H�EZ���%S�)9r(��dK�dْh�A������p8�g����q��I����ê����/Mu��TwMש���$�c��w�O��b���^3�GUU)�Ϸ��	+qW�{�<��1V���(t���ϗ�i�> �� �t+++t��z�L��o��"�Ȗ�ؼ��Yi��|�,���*I�D�@`K�w�Q4�X,fj�{<��^z�t]�������h�F��S0lh�㨿�������D!@P�Є3g�x^���?�0fB��$�x�z��L�9���C�QWWË�4����iff���4���`�$
�C�Ж��Aڶmɲ\sI�f�R):s�n� �UP� �FQ�BR=<���-)�k�w��"�����8� �U���Z���|>
�����w'���[A�V��w�v;��tn��	��\.W�fm�k��Ks�������qs�5�VZ�n0��Ԛ����i���;�=
 P
��Ɍ𿅅���x<�o�>ڱcǖ��R)���)�v�)�����
e��-��|>ڶmm�Ro��?�>��C:x� ��aS�g��r���^A 
�^�����Z|h m� M��������G�?�NS<���f�1�z�t��y���8����h�޽[���+�'�I�C�$I�Y�[)t�y�������S<7�e��]�p�:���V �VA�; t�Fۍ¤V]�ک���y����q\ÅםZ��Lj���&��*1�H������n�[�N�m��|�ӹيV__cE���mކ4�r�|%I½V���o~�X͇�~������ ���I�D?����?����===t�С-����KKK(l���]��-�i��h����M[�`uu�Μ9C����s�NS�g�e��Z����Q����{��Z|h m� ���?��O|�7�GIQZZZB�q��4�N�>M���w)�N��n(��R___Ӄ��1ZYY���iJ$x�AUF�;c�B�P��p8L}}}�J�
I�������K���O�����	 `�@�a�U��0
�<�#�K�T��q��J�����o�w��L�5�����IŪ���L��>o4Y�
�V��������g;���h���Zz{)��W���1F�,;�;��+p߼� ��n��'
� *C�; 8�ŋ��[o�?�д69����qڳgOل�Fd�Y���Fa;�$�2������[
E����UU���z��������-_a��+N6r�+�b���ԩSߴ�� �
����|�]]]b#�2��ڵk�B�&����ȑ#���/�ZD><<L7�x㖾�&�I��������c�N�i}}�<������m۶���L&M9&EQ��7ߤk׮��Ç[Z` P
��Ӕ�o.TrR�\;�mTj�F����{�.��S���^����KA���n�[�N�m��|�ӹيV^_륷�j4͝1�1ō~�	 ��]�J����o|�)�~Y�o6 @�B�; 8��i��SOѽ��K�Tʴv����ަ����t��e�r助I��޲�,�������ټڽ��������k����8�����&�����q�bC%��F�����3g����Ch(ph������}����F�___�L&c�!�M�y����[��ի��)MLL���H���\����hqq(`K4M�D"A�d�DQlj��q���C�p����L������7�x�8@��ݦ�	 `�@�1
�x�'��k�ǶR��3�HUU����N(po4�=4��؜�ND-�d�n�[����V���l�s����������K�Ks�4�c���<�r���[j�f�K��Q��q��1.  ��w p�d2IG��_|��𿾾>:x� �����c����iffƴ$m�,�1J�R�����6\�l����(��V���f��_&��C�����Q�e���`Cc��Q�g%I�����y��P�PǙ3g<������|��K݀��N�N��|����@�<H===M�������|��(EQhmm���|��r�A���x<n��#�N��/�LCCC422bJ�  f@�; t"� ��מv+p�y������F&��{Q^��v��K�@��u��IӴ����[A�V8��Ҭv;��tn��U�W�X!0����R����{qq���l6{]E۝ƌߕ�Ez; @u(p�V�t��r�-433cZ�����8���7�=0����4��qS��3i�F�x�2��B��Ɩ}>P6�%I�L9���������馛�j��SɲL�p��k�(�� ��s�=���P�P����W�o߾��}u]���E�u����R):z�(�9s��vc�<x����d����L]�� I���� �w^���m�F�\δ+TU��_����馛n�CF p�@��8�לv+p7��5M#��_��k�����d�N�6�zEqK�����H[j����
���יF���l�s����n5��T���7�y�u�r���   �@�; ��/�@w�y'��i���z�t�����o�ߩ�J���t�ڵ�� [���iuu�c#m�o� ��M;�˗/ӛo�I����.����N����nw�����~��Ň�j(p�ᮻ�:t�M7�������
ɲl�Q������[n���)S��={�4����*����իWq��b�Q2��T*E�p���㨯���^��7qSSSt��y�ԧ>��  ��� ��ڭ��hc \�4�x<u�۱��Hm�`��_�y�y�TU%�X�
��n�[�N�m��|�ӹيV\_�7��T'��7�yT�Ei��VB�; �=P� ��(
;v�N�>mj�c$�ÇS(j�߭������i)� �d2���ZQ����E]]]���f�g&�Jѯ�k�;v��&�F.�#QZyT
�B��O~�#6�k����/}�K��F��F��f����n�!��^~�e:z�(%�I���n��Fj�anܠE���5�8���`���H$B�H�0�������k���������& �V�� ��ڱ���8R�x��; �N�ͤ�����	)��V�,UU]�ZD#��|�rn���W�������Kջ�h�4�F>��,����(p �
��n���t�m�ѻ�kj�t�����[dY���)S�7ԣi�����iM�����������2V����t�����q;Y�)�4t{zz����ɗ_~���P�P�<��۷�/���i]�v_�]J�4z衇�ĉ�&��|>:x� E�ц�M>����iZYY��	Z�1F�T���dSi�@�b�X���$�+��B}}}466fJ�  �B�; �3�k�{>�'""��_s�v)p�e��٬��6���N>��ֿ��\X�(
e�YR��߻U��|�M��|[<7���L&C�1S��Km.L�4�F�Q����  �w �ӹs��[n���ES��ݻw7|o����%���-L���h*�b�qY��륁�J&�U�;��455E7�|sC)��<�J���`�quww��'n��� \	� U|��_~'
5�maee��/,`Y�鮻�W_}��v�� :t��%���8MMM����*����q7���|>���d2Y(̹^���[o�E�L�>��O��A+ �
� ��]�u]'UU���׼����]�uJ��U\���^�}�A�QTj���]
�����)�����1����|f2��g�H�6���쾾*�RC13��T#i���7��z�GM�(��Y��nG(p �
��.�������H�e���8�&&&h����EQhjj����L;���4����IQ���j螑�y�\.G�Lƴc�z�*�����O����i�}��<�����>#���s�Α�^z�)�u�;R	`����w�ٳ����d(�[|D`���u���[�������M�"����������-.."�'�NS:������d	�@�����fI�$ӎ��ŋt�����]�� ��  �Ԏ�DR4M#��S�{���Im���_A
�v���KAt3r�\�=��i�/�%j��)�r�DuUU���4���k6��,��T�4w��7����<����{�w  {�� ���S�N�#�<Ru\f+A�P___����T�$Q"�hx�{�㨷��x�7�v,�H�ٳg������cZ�`Y�)7t?=00��l6{�����I�h#�(�����s>���_M��ڵk(Jv���9��7�AW�\1����Aڿ�I��4]�t��ٜ f��󴶶F~��DQ��?�����O��P:�6�8._�L�Ν��|�3/ p�P� �L�Z�N�Q\�q\�t7�k�F�L�jj;��e�����q1�
��<����j���fȲ\5NUU['X���SQ���E!��;���뫢(�b;��9ͽ��1�˹�3�
(p �
��J������O�>���튢H��H$��������,����TU���5�����n�����H �2��ꫴs�N6�]��1�
������9A��s�=�C�U�5:	`��;w>522rC#����`F�}��t�m�Q"�0����aڻwoC�c���H���i���`]�)�����Dz��b1b�Q2�4�8VWW��7ߤ�n��� ��w  gj�w��
鹵&����]�e�$�nj�݅�� R�5M������+%I�;v��"w7�O]�	���n��[���W;��K��d�Jܘ�^��(I��� �3  {�� ���d�;�~��v� >|��@�ǁ�?p��!��PwwwC�D�p�B�����v���ٳg)�О={Lk��������1�����<����{ϼ�  � 
�6��w�>x��q��Sw�>�ɘ���㥗^��|�;e�._��۷��ݻ�W�4���6u�&�]��,%�I���j��k45}9�t:M���*�۷����  ��  �ԮŖǑ��iZ͂_��;-����w"�-������f�e�/�`����)���ŵ�<�q"7��L&Sx��<O�`�t]/+xVU���-���캾��ڒ��RF�r�"w�����<��Z���UsP� `��������]�t��vC�:t��U�WWWiff��:�|����)74v)���ʊi�0����ߧL&C���'qO�2�,7"��xH���駟�ϦCp�H�������m۶�z��NKKKU����N�:E�<��K]���Ү]��W�$������3���J�������&��C���C>���g����8m۶ʹv J�� ��ڵ��hぅ��5�	�^���\.����R<ϗ��[��э`�U�������A �狒�5MsMm)��OY��& �x<��z�1V��UU�c����(����l�t]oIz{�vJs��y��󅿯�� �� `���9���Z^^6��p8L�"��Ww_������Ғ�� `']�imm�<�����F���]�x���o�=��0ƈ1��{��������7�x���
������G{���l#��������c�����t��I��޵k�ܹ��}�����ŋ�������t��%�z�jC�o߾�&&&L}����;�7�xô6    Z�(���z�t��Q:�&Y�+>��y�� GI�<_(��uݵ�w�`�Q6�-7�D"���U�9
�(�E��`=EQH���Ϣ(&qW��f�\�(}�FQ��g�I�y��Y����)�L��:�i��~�     V������릮�M�q�С�&?��y���M?�V`����<���5T����E4=��W^��G���޼S�R����j|>�t�M?�� \Q ����������믷_.����U;	L���~��y���޳gm߾��c������E���Z-�ɐ$I���]�8%�(����fZ���ӛo�I���466fZ�  $� 8S;'��<O��c�j���Im��|�����
i⺮[������z��������n
��e���~�e�����*�|>W}�q���u���la�����M60�����5M#M������<5ʎ��wBz{)���W�<2�H�$$�o~o  �@�; �err�n��VJ�Ӧ��F�СC��$	���B��I�(�LV)�������u�z�*}��G���~�m���Q>��H$Rw,����������g�^��� #R Dt�}�M�ڵk#����XG�u������g�5����q����i499�I���]�x��Y��{�nS��u��������sS�    hAH�u�4�Շ�UU)4�Rۍ�n�Cm>���!it]�T*UV��F)
U�7<�S4-ڦiZCiF�u���y�/+n7pG�@����C�TU-\c�x=4�[�������    ��ϟ�[n�����H$Bh�;���
MOO�f\�Y�$�G}D�L�H�<h��s�����N�$��.X�K����Ч>���� \�Y�  -��/~����ޞz�%	�o�����w�M����m������H����<]�t	_(�#��J�x�"�H�%�}���M=�>��� MLL��. t6$� 8S;'�m\��J� T��tJ����^���Hmw���)�����W��^��[��Q�^���bj�[A���B�>�Ƙ� �K���M�S����FVT0��K�I8��n��u�*N�;��4�j�GEQ
W�yHp ���z���{t�w�c�!7����+W���⢩�8��������W0��~�����eS�VVV�7��}����|EJ0G.��p8\�;�C�й7�|�w6�caD
:�w��}ccc�����Ř`EQ讻��_���w��A;w_6���?��c�QE��/R"������0��U����=��#�����v    �f=��a;����J���^���FmNX��t]�t:]�p��8����p�`�O6ۜ2�P���*�b�֢(V|Pj\p��y�7�C���(���    4��ٳt�ȑ�I�ft�������1������S�p2]�iff��]�Vw߮�.:p����SSS�����gs	]�iuu��~� ��>��c6��!�:�_��_���b��[YY1�f ̧(
9r��}�]���ݻw��/�c�-�X�1J$��x(�ܷ��������f\�p�8����. t&$� 8S�'�sWH����eZ���N���|>���nl����kQU�2�LQq3�����Wwe�R~��dY.jKU�TP    IDATU��|�����z�gv�FΥoc���]q�a��u����sK�{��#c�$IB
�u�� �Hp��:{�,�}�ݦO>E�>�O�QU�&'')�ɘ�?�[��iR����j���H�p�� �d���}���>�$wP�DQ�;~�F]]]�y���/�th ��)�hw�y����X݊eI��e�t]�{ｗ>�����={���oyy�fff�\�1F��󴰰Pwߝ;w�����p��I���~fz�     v�c��<�Hj{0tMj{)��W(�U��	���(JYq� ����tq;��{'�m�4+�dsa5��M���+�c�N�u�r]��7
�1ͽ~�     �|��t�}��^��������u��eY��>��$I2� �Y]]��������X�&&&L�~~�n��J�Ӧ��[]]��^�y�>��<d�!8F����ܹ�F�YZ�1F��{/���릷�Fi�޽u�[ZZ�+W���?�[---���l�/�w料�>����L���/Lo    �F����c$�2���L}>�B!ץ��D"��Fque���%�{<�-�|>uwwm��r�*�u#Y���#�;���V\�M�u�d2��f9��bAp�º�**���c��dj��a'�=�ƉW     ������#G��~�,�x�u��%I���Iܷ��D"A���u'���ؘ�������ߎ	'.�(
%�ɺ�������o��Ol8$ �B�;t���{���hݪ�D"�/���|�^}�U�������@J��4����OLL���1F?��襗^2�]     ;��ND���.��S�Ky��B:���-��;M>��L&St�������ה��P�,]|s�84GQ��Ϯ(���'��C�`��3o�c,�����I;�����4wEQ���    @D���[R��q�߿���p��2�MNNb�3@�L&C/^�;�822B۶m3���/���N�\����\�x��5��y��?���6�#aT:�������5M�x<n��V=����_���v}>8p�+W���Ғ����x<N���5�܍$��.�^c������ٳgMm    �jǑ ��jKpMm��Om/��!.R�/��Q6�-����(���H�F��SF����D���Į͓7���x(�3�(�Ͷ���I6_Gܞ�^��i���m1    �033C��~�%c�w咽������i�t�B �0V7�W��gϞ�����p�=zc3��:�����o׮]}����6�#��:���ǣ;w�<Po���5$D9܉'詧�2��F�mc477G��˦��n��$]�t����F'�4K�u��{���3�]     ��<O�1�Ӱ:-���(��B`EQ06D�����H�X��dd��)�m�4���9���y�'��.r�d2���M��m�5���S�܍��v�[    �inn�n���d2��=22BCCC5�I&�455���:�"�Z��Ɗ	�P������w��LDq�L&S7m_����� �}GTj��|�x�ޚ���yJ��6l�O�Sz�',i��n�H$R�u����64� 6��i����Y�i����?x�4���N���~gj�     V2&�� �1F�$udj{���:��Z����A ����
v}>uwwm��rH�j�,�Ec���bLx��L��f;~I�\.Wi���RNLs7�(p   �vp��5���GJ�R��=00@ccc5�I$4==��v�ɲ\7�]:p������z�-z���*�í����gbbb�+_��6���:�;���\��P��lgϞ������1��b5�����x<nI� �,�����T͛�h4J��������ȑ#���`z�     V0���(�UU���d�bTA(
�mj{)Q�~����R�r0�h4j���x�m&IRǞ�F)�R4!a�{�*<�W-r�4A�S0�
)���^��4�T*e��6EQ:�w    �+�N���nI�B8�������R)���A�,@�r�]�x�f����o�ђ��_��Wt��)����r���rx<:|��Ol:$ G��t���ϟ���5�H�T��28ǅ����橷��v��Qs�����f�@e������}��i���(�H��6    ��8�#AH�4� 2�(��R:��ڇ��Z�ڮ8��p8LD��NK�f�Q:�.���-��h4ZT���:e2<P�B���1M��kIX%�U�NȲܑc����^�^���Y����:1�:bR    �7UU��;�$�����-�M��4==�{q�-��rt�ҥ��tF"KB ��N�>M��կ,i̱��V�{�7���/~q�M��(p����v���������u��5:z��%	?�@����W����ի���bz� �&�H���l�/�{��)��iii����ou\�
    ��QY+�g�����"��}�B!���Y 
���|�c��J�s�H����l=��)�m�4�c���f���{����f�{�޲�I�j'�'�tr�x�4wEQ,Ks7��Ŀ_    �>ct���ӹs�,i����������fizz��\'I��ҥK5?K��ôm���ˌ1z����?4�m0�1N_�(����|q��q:wd:��?|{ ���L&mY��J���n��G}+A�����LSZ\\�k׮��7@����t��媯�<O7�p�%K�ONNZ�    ���BQ3�u]Gj{8��P(DD�����L&S66���M�H�%��������h[.���]	Y����(�����8E�⽼�(������Z�殪*q�w    p��{�^~�eK�+�T��Q�[+u ��f�ҥK-	�4����o��ܜ�m�9�D���7��?|�ӟ.O� hc(p��2<<�׵^g�Q<��p�	���w�AW�^����{�ZW���B����������j.�hbb��o��=�裦�    `&� Ьb^UU)�JUMm�x<��^js����v��:�R����h�昉B�PY�$IH��w����W+0��q*&�+�B�l��?K�5����Kٝ�i��   ���9s��x�	K���������r9�X �����t�q��h������H�D��ַP�P���|�D"ܟ���g�!8FW�c<���K,��'�L���n}��G��?<<L���U_O$4??oI� @���D+++U_�7�r=�z�)���nI�     f�8��^/�~]ż�1��o�qn'1ƪNp;����=��
����F�����\(�]�I������|>_�h�Q�^�XE�y-r�|>_�,�zZ̮4wM�H�u�   �k�ۿ�;v̒�EQ�}��U}]�4���2u5A ��d2Y�IE��,�{yy����ov�J�n�H$�^{<��m: G@�;t�m۶=Xk@[�u�Rs�S�N�+��bI��`�v��U�uI�hvv֒������)�HT}}�Ν���eI�?�0�;wΒ�    �`�gluR��(�L&�g{�^
������|��,
�1�1�]���bc�㨿��,5��x�/[:]Ӵ���N��f��<�S h�E��EӴ��*�n�D�Wgu���    n���HG����|߾}U�Wct��%�Xluu���������C��Ö�=55E�����n��0�j�����կ�W�	��0���ɓ��u��'��{���}�]:}��%m�<O�����CQ������&�����f��>11a�R\���]w�E��˦�    `�{p��~Fj{�$\��HE
(����B����m�⮪*��颱�穯���^o��2��G���E�r�ܖ�`�N�墂Q�X���+N���r���r��	P��i9�     PO.���G�R&����z�b3335���yh}}������
�,���ٳ��3�X�6\�z�9���o���6@Ka�:��i'k=P�4��ɤ�G�X^^��~����ܵk��ኯ�NSSS���t]���骟�@ @�����J���ѣmU�    �C�8��{T#��Vj{("��g�a��H$R(��e�-�E�L&ST\��x���ב��P(TV,-IR[I7BQ���zQ-�n��W1]�1F�tz�+T8	�۷��4w����w    p�|����,i;����H���&�����(�NW|�㸚�����G�?�В�a�c��k�366���/��M��R(p����GGG?Sk��;O>���G�R*����X,Vu9�MMM�$I�� ��[9app����-�{zz��?nI�     ��H�e���؜�^i_��o�q��$Ƙ�'�+�B�l��P���P,stq�!�sI��0����[y�^WLV�z��܍�9�ލ��|ẋ��昙�i1�p    �u�y����mI���n�ᆪߓWVVhiiɒ��:����T)	�B466fIߺ��=��C�����[�N�k�?�@������2x�m�G����W}�#�ݙ�;F��Ӗ���zi�޽U__XX�:C �'I���V}}�޽���-���^�_|ђ�    ���\k`���ڼ$��'�����"Q��G����N ߌ�y�F�E�4M�\.ע#�W6�-R�<_�h�d�u��Q����#��B�>��(��"3�܍���    n��Gѣ�>jY�{��z��d�ʕ+�� ���Z3p�����,�;�Hз��m׎Ǵ�z)�7}��w�`.�u���m۶��Z�'��Iwr+g&mܼU{����N��˖� �I$USA�9I�z=��C499iY�     [a�WJ8f�Q:�Fj��A�`0HD�Mq��r��f���|>��b���[�|>���.�&˲+�K3dY.��S����6V�p�9T�0ƌ�����4wUU]��    �ζ��Nw�y'i�fI����UW�VU�fffP3�b�,�����,�brr+�;P��H$�����	�%0�
m���t___���How����[:39�Q___��dY�˗/[�7 4gaa�R�T��zzzh``��~E�;Ｓj�     � �<_���H��T�N������n�p���LnKq�e��EQ�X,�ڂ�P(T�@'IR��+�S��N�q��61���x(���c��d��D�THo7�V��c�i�k�i    �yTU�o�۴��nI������S�5�MOO�r�1@;J$U9�^/���Y��/�K:s�e����Kq߿�_�t( -�Q>hk�p��k���vg�d2t��Z63Y��7o�����t�> p���٪�������Z����
�s�=�    �"�N�����<�S pe���y<
D�1������$Fm$�����4�%X���v?��z������+� T]Y"��R.�k�Q5OQ��u��'�i6���	    �'N���?�ز�w��U���ʕ+��d,� ����@�t��kCCCe�������9�ڇ��Kq߱cG�o��o�G	�vm��u������o��:�۝�رc���bY��v�"��_񵙙�<4�$�����tŇ�^�����-���>��޲�    �e$5������PȲ	��ns�{iѸU*��F�b����F��i��v�<�l����4�ޭA�`0X1����'2& ��:���!	�h     np��yz��-k�����m�V񵵵5Kk3 `kc433S��y�޽���*�Bw�}�k=:E�w�������l< �a������^����d2�4y����ٳ��_��mii	� L�$�r�J��(�Y���~�#�R    �0
@7�o��v{x��B���i�}�c������ۦ�������dYv�i�,�EZ��3��|�"wY�������1��+�O�6��UUm��    �/cu{�jVA������ɲL���� �OUU����x}422bY�sss��c�Y�>4/�NW�!"ڽ{�����=Uw p9��B��/�^�u�r��5z�G,k��y�����pC�$�z��e}�9VVV(�HT|m���Un^/�R    '�j%R��
�
�]Z@��1�f�e?"�uuu�訬
��R�%I�8�ME)J1EѲ{�V�8�j�{.��L&ӂ���87Ho�����x��=�y     7�zu��������c4;;��{e�v��dhii��k###Ec�f{����?��}h^�Z"�p8�����7l< [�����������E���J����!4M�����$��۷׼yC�?�;\�|���TQittԲ~����ĉ��    Ќ��O������+S+�R3E�n�1�d2eu���)�:\���(y<�,�u��٬k�~t]/3�z����ZxD�2��+M�Q�2���Υ�(�i!��nǑ 'D�o!    8�ի�ھ}{���J ����"e�ٲ��ў={,�1F��w�R)����R��T%{������`+��B[E�x��l�����ɓt��E����|U�癟�/J� gSU�fgg+�6<<\q"�Y�y�z���-k    �Q��w}>R�[hs�x.�k�����J��
�Ѩ��NN��<E�Ѣm��:��4+��B:x�/K�oGǑ(�U�ܝ4a�x_!��ux�'��[4� �    �ɬ^ݞhc��J�(�T����-� �SkŅ��.��﷬���uz��,k���9�`dd���꯬K�h!��A[�l���鴣R�:م�?���}���UL�I$���ji� `�j/<�Ӯ]�,�1F��?f)   @�y<�y�B�������z������8ɹU���҇^�X���`���~>�������ɲ\�h�t�,�av�*F�{��zEQ(�N���}��(�n=#��    �L�4��{,MP��b���S�ﹹ9�� k�r9�����ڮ]�,�~뭷��_��}hN"��8فh���C���� l��>h;?���s8.�h���D"a�!A�\���ު|��Dh``�l���t��e�� k-,,T\}����,��L��������    �q�B�����~�S�[�J���eE��QG�~�2&�l&I���PfR���$�b�}�k�k�Vq2�����<<�w��    ���'���?�ز�9�������κn�7 lX[[�x<^����ӎ;,�����a��T311�l< ۠��N4�z��$Iv�x��hii��>v��U���˗���b�R\������-}�|��Yz��-k    �(�t��������VUUJ��E}�<O}}}��zm?��F���x
?�N�l������^����z+yw
Q+%lVm�;����v     h���=����1<<L�@�l���%�IK� k���W�s�8nbY��رc��ͩU��ż_��W�����F_���<yR�Y�u��;���$=�쳖�100P�5Q<�� �H�Tq�p(�m۶Y���>H�l��>     �=Z��(
e2��"_��C���]�N�Qx\�ʗ����m��f���)BG&�����1J�Ӥi��ǃ�v     hc���~K��^/����m�4�,� 졪*]�r�l;��466fi�|����+���Q�j�
�q���o�|H �C�;��l6�5��[�B�Ҿ���ѱc�,MW�y�v�,���z�/| �N������˶���Z�$���:�8q²�    �]DQ,$�ۙ�n<�؜H���b>�������ɲ��eY.J�E�����UL"�u�2��m�5j�Vx� �     ����Ӆ,�ctt�h3V�h���=([�����&����Ν;��x( ��,��X,�ߪ��?��������-�cpp�b�����c`@�t]������>�����,�ێ�(     p��
�c�$���y�d2E��>��z{{-���F����_�$�&"4�4�CE��^��f���~�9Bz;     4b}}�{�1K������&�I���� �����8�U)�L�T�~��Y�4F����]]]�7�񍿴�� ,�whgΜ*��i��i�	J\�pd��    IDATz�N�>mi<�ӎ;ʶ��iZ[[��o �_:����ղ�;v쨘R`;�     ��{�|>oi�t.�+[����Q,CAt��⺮��߷���$IR�g��K>���G�\^��B�PYq9c��٬��麮#�     ����R&������Ѳ{$]�i~~��~�~���իW˶�b��U����/ӻ�kiИT*Uq;�q4>>�5��R���q��廪=�K�R�y`թct��1ˋA�m�V����˗/[�/ ����B��z^���o�ny�O>���}     �;pG�P��6�!���%�Ȳ\TM�Q���Pp[�qe�E��ڒ�߈l6[�!Bŕ	��A�@ P��g�Q&����g|���     �x����߶�Qipp�l��e�F �Z���e�D�]���C�@��N�IӴ���ܹs��0pmO=�m����Y�ת�\����t��9K���޾���� `>M�haa�l���)�DDO>�$]�r��>     ���`!%<�˙� IR��@ @===(no@��qY�[�2�,�E��EQD�t<O�"w��	f�"�     ���d�����S)�]�$ZYY��o h�˗/��=���Pww���.//��?niPc���t�ׂ� w뭷��6�e0m�̙3b___��k�L�,��%I=��c��344D~��h���t��5����Z[[+����x*Nz1��������>     �JS��,��T�)���	>���^o�6I�
��vS�h҂(�Tm�J('����&�\�-���    ��N�:E�D��>� �m�����_ h=I�hmm�l�Ν;-���瞣˗/[�ԖL&�������͇`�C[�����Zr��[��ɓ�߼�<O###eۯ\�Ҳ�� `�JI�CCC�������{�Y�     ���b�|>�)�FO���p��[TZD��:e�Y����u�$I*���z����z��y
�B'Ȳ\�;�*#���yL@     ����矷��J���x�2���}@�-..��Cuww[��i=�裖����Zu�kddd����
ܡ-�b������$��]7o���e	\�l����-� �!�ɔ}�=m۶��?��e�    ���b[�����Iqg�Q6�-[�0�PWW�ug'�8�DQ,ڦ�������f����� �4��8
���s��uwȲL����#     *9~�xٽ��|>���mc������s(�B���eۭ^垈��ޣ����~��j���`���׿�_m> K��\�w��������Dr�ӗ��E�����p�v,��y�^�Zv���\����     �
�
	j[Mq7��K�T���)��r���RA�,˶M\�e���AE��_'�Ƚ4 �h�o&���gqsz��+�    ��ٵ�������#����V������\���(Z��#�<B��Y�TW)�hc�l����O	�t(p����~��Vz�`<����ok��[�/gkkk��f-� �%�����R�6��O}}}��}��IJ$��     �V�����e]�)�J�= ���)�����CK�T����JW��ǡyF:��bEQ(��6]���
�현      �h�F�<����@CCCE�E�k׮Y�7 8K���Hq�r�
B �Zm����n��(p������J۳�,f����i��������ۋ~f�����]�v���o��$It��I��     �D"�bXY�.�5��K��c�ӏ�Ӊ�XT\��������:I�T����VL���8��@�$�t:���e�Q>�Gz;     4��矧��9��*�(���h��m p�D"A�L�h��� �|>��>y�$�R)����R�Tű���n�k_���ւC0
���c�����J�!���~�_�r��D����h���j�< �9t]/��
������_x������     p6��
��1�HQ���FӴ��[�㨿��DQ��X;���������+e��B�� 8�1��+=��4��$�J��     ��d2t��i���8�,�=����ښ�}�s]�z���J�
+d2z���-��SU�h���������|8 �C�;�ډ'�������UU�l6ۊC�H1>u�-}!� *YYY!UU��ّ��:=�裖�     ���]�!�AUU�d2EE�<�Soo/�-V��\��{��Uڦ(�(���(����˶W[)a3��r9��    @CN�>mK�q�I������D �N�˂`�����/}��
��^�B�����|( �C�;�����#�����_�Ֆ�7��K}}}E�VWWJE��V)�=�R ���>��Ο?oy?     �l� R�u]�:^�(JYq�����^[�"��W6�`s���R�h�C ([N����+�3�(�N��i���    �Q�����_�Җ�J�s������7 8[i���㡁����4�N�<iy?P]�ز�����w�w;[pH �A�;�Z__�'*mG�{�d�Yz�gl�kpp����`������m۶�ҷ]�X     ���KqW���lQҚ��X,��v���XTt��)+D�N�$~�z�8�6���e	�D�&�ɔ��3�(��#�     ��OP.����`0H]]]Eۮ^���v  ��"��0���A[�~��hvv֖��c�2�L�v��idd�-8$ Ӡ�\�駟�D"e1V�,#����zꩊ4�P�Elyy� 
*Mz���e�s��ѹs�,�     ����
k5M+*���r��d�D�|>���EQmpWV��jŉ	�؜/B�Bk���竸��Q�yL1�ˑ�������     5���Ћ/�hK_�A^�,S<��o p���������
+LZ�1F�O�����tr�add�?�|( �B�;�V"�������N*��g�}֖���hї0�---��7 ����j�Cj��O�X̖��q[�     g�D"��6��eY.J�&�(���bE)�`�J�,�%|7��ߊ�����z��2�(�͒�(�q\!�I�     P�O~�[B�8�+ \\\��_ pI��
��Z���7ߤ��[��r�\��ߣ���"$�
�������c�jKn�=~�ӟ�=��J�����-?l��������mv��]�p�~����     8���-M�३�(R,�e�)����6oNao��(E�9`�x<
�e�qeI���     Y^^�_��W�����_��[>��D"aK� �.����2��C`�U��E�n���҂�0���+1Ƹ��������_2��_������x����h[i+ �aee��oCOO��~[�>q�1�l�     �+��4I'POO��DŢbt]�)��6��u]/
��z�Hw��C�@��gNUU��    @C�q�B�����~^^^�3H �(�N�Ky<��볥�w�y�.^�hK_P.�NWܾcǎ/�|( ��Sp�S�N}���M/�v����'?)K����@��D"a[� �>�����j�6�R�/]�D���-}    �s�|�B��f�`���(���㸲�e��7bs� �=�V�"w��    @=��+��җ(����U��ҳO �͖���~��>����ɓ���E�|>_�}pp�@�(pW�u�k��@���iz��m�tfa�3 �R�)v�P&ژ      �9������U�0]���|�����s�P� P0,J�Gz;     4��'�,ZA�J���E?��^ P*��"���m�x�|@������*��������/���p �
���b��gJ�mNF{=��s���l�����N�$�2��-}�{��y��ㅟ�� �A[�����.��     8���#��GDD�H�h|����=��5�(JQ�{ (*���y�����  ���w�O�]�}��O��LO�E#���m��d��8H`"	a��$0&%��<IA���E��T���[�R�ۂ�mb�I0�d�e�B����s�{?/�iuό4������rU����-M������ �|^��x��ko{�������^��@3UU�������^��2{��_�zmc�ӹ:t����w���ā˦�N�<��ˇ��+9�1�N����^�xG��������:s��s����  �k���q���X__O����o~�^�elnn���;�v��`�$����z�o�>g  ���׿��d佴��kkk[ߟ<y����f{��Ww�Pg?�;��Ύ�=���f�<��رc�� \6w���>���R��/��Ϸ����"ﵣG�n}]E�c�6w���s������K/�6  �����/��_�׋���6��v����d�~�+++�e�������  ���x���7j����No.TQ��k�m}�����%����k����p������Q�)��8�~�g����fTU�"N�UU��?����[^^����<����^��\�W_}u�����s�^���  ���UX�F[��F���f[����Ei  ���?��8u�Tm�m/��F�s����~DD�� ���Qlll�6o:}��Yv�С������ �.Qp�q>|Ǚ�!>��~����H|�UW�x9x����<yr�Ƙ+�������O�$~�_�6   �gii)���?�g�澺��~��x   챲,��_�zm��۷/��۷���ہ�u�-�u�#��a�7^��l��dǟ-,,�����%��L��F��7��x�����VU��1���?��Z�;r����g]p>g^õ}^�k��$���o��  ��ZYY�Q^/�r���*�  ��/��rm�m�YUU�<y������~x�bii������pǭ���\��_{�O&��E��F����ę' ��(�2Q������������6���b���o}ow2p��/����w�5�{����z�NY   �����������r͉   �K� ^q�[_�<y2���u|�μ�~�ܲ�^{�����]�x��\�+���Q�(��(eY~��?���L�����/��w�����z���X���z�������Ç�6�/~���w�S�x   �~�Β�����gW   ������������6ޙ n?��bE���C��:~��2�0�Nc:����Ç/���o�'��D��F9p���ۿ��J�=�������w���kN�.�k����u����o|���  ��ZZZ��`�����j�y�$   �Q���� ���s��p��o��>���瞋��ǵ�Ǜ������~�t�M��(\w�СC�?�L\Ô���ٟ�x<�m�^��c���������v�>�<x0�{$�ۿ��������  `����D��?��  @������?��Z��~ �~p�666b6�E��7D����j�7���૮���	��%Sp�1���o���`��g���i��౶�KKK1���N.�d2ٚK�����o  �l�^/VVVbyy9u   ���O?}�)�{m��
��n�>��}������z�*o�FQ��?;r�ȭ���%Qp�1^z饳��Pp����?/��B�c��x�����vJ���ַ����1  �]�~��+�  ��7��Z�ۿ��Ma�Ѩ�r=�N������u�#677�g��uL"��:�w�W\Q���p��i����m�~6��d2I���^�ED<xp��'O�>>�N�7�Խ�;u�T��_�e�c      �����g��u�C�m}��v`�lnnn·���������o�ه��������ݛ(\4w�СCǷ�������x��k���Ł""b:����F���5�N�~��۷�      ؒ� @w`7m�S���=���?�a��?�c�c���o�D�K��N#|��\ܿ���?�F��t��O?]��Wkkk���#���}�[!z�^�߿�ֱ������ӟ���1     ��N��g�g��;/��C�`W���u�h�������1��(��L&;��+���Dq�)���/,��q��hM�7�������@����>>�n���/���~B���o}�[��	      ��3�<�O��u��������͘N�Q?""�O��O�(����3;��>�(
\4w�ԩS����x<��,S��W_}5~���>��^�elll�>>�n��d��;�S��       ����~��1�N���[�s���z�z�Z�~�������U똜]p?p��J�(p��i�����m�����{�駣���ǝNO�:�d|��N�:ip/��r�����	      ���p����kwޏ(�"677kh�y?baa!���j?�桮�F;:w���������&�L��FX[[�a��
����w�S����˱��v'{g~�_�ߏ}���>�������      ��/��/b:��>�����n�5�.�<�L�f�����b4m}����ꫯ�F���N����8p`u��1�SFꜟ��g�����>�������� �mcc#ʲ��7?4�ӷ��m7T      @&RP�����oTc܁�������lll������>n�m/�GD>|��'�E����ɟ�ɭ�~�7���k3�{�ʗ�pF�QL&��������M4)NpO��      �icc#~���>�� @`o�7�l�w�������:t�DQ�(�������Sۿ?sG{/Ճ��A���k�y�      ��g���lV��������I��c^p_]]�^�w����{�gb:��>n�M&���8p M9.��;�[ZZzp��
��z���^H2��;P�ӧOGDڂ��I       ��|�;IƝ������+��0���^�����p����k�˪��ѹܷo������$�D��쭮��:������)�t��O?�d�~������e��4��(�X\\ܚ{��ꫯƳ�>[��      �N�:�7�d�y�T�����FDD�߿?��n��������B�|��K.��;�[__�b��x<v�m;���&wmm-z�^�F#�o�H}�{��      �����EQ${����@��'�GD����?�,�$cw�p8���W\�d�(p�����O������4�~�U�ӧO�s�=�d���m�@��R�P�����d\       ����������~?�� �Z� LՏ���H�I�3^__�'a� 
�d�رc7/,��c���������d��VWW#B���|7����/�ɓ'��      ]VUU��?H2�����J��6���d���t�������L&[�<x�ڄq��(����^zi�UNp�W�ӄ܁��p+++IƯ�*����'      ���矏�_=������ԧ,������^/I���o������_K.��;Y�����_O��d��wQUUI$���b6�9��MUU�����R
p      P�����p)�u��؈^�������j���kkk��d�)Y[^^�u���s�^x�d����$�ݵ��KKK��������}�f.      ��_��_'{ee%ʲԋj5�T������?�A���j��~���?��{Ɓ�Rp'k���z���z�\����X\\ܱk���0z�^,--%cc#�{�$c     @�>}:�;��������i��Z]]M��-����fQ���W\qœ	��y)���}���ͿVp�W�oY�u��;����H��      �&�-�+++�@���qTU����7�UU%���w0����O�K��l��_��`ee��ƕ$��$u����܌g�}6���b�܁��p)��     ���|?������
�@���h��q�ԩx����E�����9a8/w�U�?��z1�L�֪�������n���[Q u*�2&�I���?��[K      �&?����=/���0��#""��o�6��]�������_�0
���;������_;��^?�я�������Ȧ ��pKKK��/�"��ޯ�j    IDAT�d�     @W�����ӟ�4������R�FI�
�u���ܷo�j�(p^
�d���_���^����R�F����4C�y      � �����1�L�(��9�n��3�Ͷ~��۷��8�-w�5�5��N��E�=�\�����9�L���     @�.V��FI3 �5�cqq1z�^�'O��W^y%��]4?lx0���,'�oI��l���_;��>?��O�/��;�R��1�f�я~UU%�       m���)� ��dUU%?��?�a��f�{����ѣGߛ8�%w����r8��_��#���'�iM��䋷���x���f      �6�N���/$�0܁���i� R��<�.	�=w�����/�_��'�C�׋��E�@2��,z�^�+�"���      �f�=�\�n� ��r��>�Y�d�����;F����N����#�N՚�.T�z�XXXH���-�S�-�      `��GD8�Ho2�$/���⋱���4C�l�孬����Q�m)������k�~���:�<y2^}���1b6��� t�d2�����I�>�l��     �͞{��baaA�Hj2�D��O����x���f蒪��:����Gǁ���N�&���۾N�S~�����^Ϧ ��t����ӟ��u�      �Gr�HTUEQ��tX FD��?�C��2�d.--�O�R��	���?��?�x�A�i����A��d ��$z�^�UUŋ/��4      ��x<����g�c�� ɍ����������'�#t�� ڕ����Q�-)���S�N���DZUU�8��C����Y���f�,p9��      �6?��O��8�H�(
���@;���[Rp'KUU�+�͝B�#��p
�@r��,�+�r��     �mr)R�e�:�q��#^|�E�~j4�e.//��ˇ����,-..�pS�����^z)uw �,�r�`      �$���܁�r)�O����O�:Fg��y�<�=��p�[p�~���:���KY����z�<8�U�eWp���      �I.M)�9��*u��Б�SY�QE,,,������y�\��������7��`����w ��,����S���ɓ�c      @���⋩#DD>''ݖ�\�K�+�����_I�I��,-..�F(��)���UUe��tWQv(     @���q�ԩ�1"" d!��V.����w3WVVޙ8
���;YZ\\\Qt��K/��:�8 ���i~     ������~��\梜��.�������i���)����`0�N�ٜ��/��r�[ʲL ���~���      �5rz��� � _y�}��Op_ZZ:�8
���;Y�\~qv�+���:BD��x�� ��(��      �@�`�\���,^{��1:c^p_\\<�8
���;Y����	��w�ԩ��cDD>L ��G9}�      M����\�Iݖ�f� �g~ �`0�"q8'w�SUU������^�7�����f��      M�Sy2�w�@��4�H�g6�ED����Z�(pN
�d����jě({���l�l��q�ԩ�1      �r*O��N趜梜��.(�"�S�sQp';EQ(��,�w 9-�rڈ      M5�L���_OcKQ�# d��ʩ����4�R�sQp';�^o_���:�T���	讲,���,�      ����+Yt��;I��r����c낢(���)��%w�SU��k�Sq���AUUY}���<      M��{7	 9�E/��r��2��bqqq1u8w�SU�zY�Y���?�y�;���)�y      ���W_Ma� 9�E���ZVyڮ(����
�dI���>}����=�_���#��!H-����N�J      O?�l9�EEQ���f��Q�e,..��%?�dg2��)�����ө#��C@�     �����M?H-�y(��Hm6�͢����%?��h9��s�l8�l6Kc���n�m��6      h��J�����'�yHG�>eY�1y�IvF��Jn��6�m����-�m��x     ���{��r��t$�SEDD/u8wr��[���r| �����.��H      �4��w��$�=9��r쳵UQ����ɒ�;9Z��� j����8 ��p��8��i�      �h��&��ґ ��qʱ��V��=����;yr�{�r۝�_����s��      �&�Ҥ��R�s�~D�FL��ɑ�{�,� v�u��     �KWElnn��q���#ǎD�����;�Rp'G=�f}r,���H)��[D��5      4���F�]�\�Oݐ㼨Q��l�:���;Y��g[M&����� �J���t:M      +��m����!�M6���mU�_DdI��,�����r݁�g H%���      .]���r}?	�_��O��u[�f3w���N���H�3r} ��
h�\�\�k      h �����|�V�{�+w�SUU������*�(��r�d��|      M��ReY���B��,��z�e�YRp';��t�:C���@�k�h������(��      � ��m��L�v�u��uCR[��+w�3�NG�3tI��\��v�y     �K�k?""���@{�Zl�y�n#'��+w�3�L��^��,����<��<_     @�r>P*ג)�n�v$r���(ןPp';���	�5����/O�n9p��|      ���@)��n9�;9��m���ݦ�NvF���{�r~ ȹh
�S��9��      ���߷���h��{Y �WQU�p.
�dg8NRg�^��:�[��A
h��?8�y�      .]UUY���'�9G?�^9�,�m
�dgjV�SGxK~yu*�"�*�M�9��      ���`�:��r P������ɹ+C�)����(��k�sa������v�}���     �K�s?""���@{����}���Nvf���{�r ��a
h�����k      �Y�J���h��̻���|�6��<�]
�dg<{b�Q�p@]r�o�     ������,˨�*u��#8�_>dI���T��r�ڡ	�!	      r�{?"BG�G�sM�k`�)����t��^����ʾt
4_���k      �Y�j�{K��r�k�0_�IY�k�'w���^�&<�f�����}�ь�      rՄ����h��(�?l�	�5��ܡ��@���&�3M��      WMx�ք�)�lM�H� @ B�:oyy9u��j�\M��hii)u      h�&�#"�q8�\M�c�#�w������p^UU)�{�)�ˁRG      ��Z[[�����RMy	4OS:X���# ����SMy h��A���2�4e�     ��z�X[[K㼚��h�&��#�#�7(�C�5偠)X@�4ewr��kč      ��&t$��h��l�i�\�=w踦<EUU���LS>ڷo_����1      ��8�:�i�{L�Y܁&Qp��k��-�9Y@s4e^qz;      \���w�N��# -Ӥ�E܁w�&=X������ܛ�	      rՔ�neYFY��c -Ҕ~DD��l��Qp��[ZZ�����1.H�v�kҜb�      ��)'�G4��
�I�6e3��܁F'-���Ҥ�[�>h     �\5�Ѥ��@ޚt `���w�Q��,���PUUE�:�k�<      �j�{��,�,��1�hR�j0���J�@܁���+SG�`M�Q�is�UW]�:      4^���*����f�#\�+��2z�^�@܁8z�h���\M�G�6O     @���ޭI�T OM; �i�4�w܁�=4��
䥪��}�w      �|W]uU,,4�.U�eE�:�`M�Y5����<�{�i�I8�r4m�a      ������ÇSǸ(M|�	䡪���!����;����=|�h���������c      @+4�#1�N����1�jZ?"�y�{G�h��-"b6�Y��(�(�2u��b�      ���	���Ă{�h`o(�������O�TUe\4�7      �&05�LRG �� F�H oRp"��M,��4ucL�g      �U߿�eEQ��4H{UKKKq����1�L(���\Qp��N�QUU����3      ��ꫯN�4��
��� ������z�c �Pp""�nH�X����ES�g      �QS߿5�@/�~M�/�:?{C�����n�)u�K2�N�,��1��5y���     �ݳ���N�L&���h�\q�7�� dD���f? 4�Tf�>M�'�9���c      @�4��&��ԧ��DS�f`o(�q�5����J����f��+�"��H�X�     ��k�!�UU�l6K�XSOo�Б vRp""������_�:�%�����3{�ɋ��~�      9kr����?��5�͢,��1.���j\y啩c Qp�X�mS�e�O0h�      �j�ASM
�&��n�����z�c Qp�4y�w�\��q�����2      ��뮋~��:�%k�{P`�EEQ��q� �I����8`���\���ǎK      Zg04�]\�߅���) gRp�4�����}�����x���bqq1u      h%� m����#܁�)�[����k�I�L&���*u ��(b�-�ܒ:      �V��Ǖe��4u M�������xG�@f܁���w��pY����Zq�C��c      �٭�ޚ:�ek�{Q���f�Ɵ���w�3���S� 2���ІB�Sܡ��pz{D;�c      �����cuu5u���w�]ڰ��}
��mx`���o��i��[���G���      ����7�|s��m<;:���G8 87w`�cǎŁRǸl��$ʲL���      p��r�Sܡ��p `D�-�ܒ:�!w`�^�ך���<��-���     `ﵡ���{R� B�����k��6:�:�!w�,mY���$g�´e���      u���[ca����d�:P���Z�o�-=5`���	�Umzp�F�# 5h��myy9�?�:      ����j�p��c��t�@��xUU���+ �w�,7�|s��1vEY�1�NS� �X�o��rK����1      �n���v�x<N�cEQ�����w�,�� n����1vM�����ڶx���SG      �θ뮻RG�5m{w
��MY�9�]w]�@�܁s��{RG�5UU����i4�����     �>w�qGkn��p ��d2��(R��5��w_�@�܁sjS�="b:��l6K�e��8ʲLc�9r$n���1      �3�����nKc�TUպC��,c2����� �w���;W_}u���.eh��.�z�^�      �)m+Y�f3� B˴������W�WS� 2������+u�]��2,tYOh�g      �m��>���m*�B�M���mZ���buu5u c
��[j�n2�DQ�c �������~�q��c      @�\��q�UW��������x�:p���o����(�o�;��`�:Ʈk���%m���[n�����1      ���X�l���5m������K�xK���q�m�����ʲl��F�
�7      `���}][߯B�u�ʑ#G�nHȜ�;�N�8�:�L&�| ����QE�{���K      :��;�����1v]UUn��j����w_�z��1��)�o�=�yO,,�s��K��(��L&�c�o�1n����1      �����[{(�l6��t�:p��kz�{ߛ:� �l���СCq�m����'�R��h�����?u      �6���FQ�e��h�����w��]�c ����<�:��f�=ڤ�����2      h���/VWWS��3��0u�<�|�}�=���U����y��=�~��:ƞi�Gh��d��,u�=s�����R�      ��q�}����gʲl����tUU�~#J�Zv��;p^�_��_IcO�è�*u�EQ�x<NcOY�     @>���n:��t:M8�����9��rK�@C(�����OaOua$4MW�]�}~     �&���c߾}�c��h�{�L�]������R� B�� ��,..�����pR44I�w&GD���k��&u      ���A����Nc�u�},4EWnVx�{ߛ:� 
��Y[[�;�3u�=7�Lb6����ׅ����      ��%̮ܨ�+˲r=z4���w��4��;p�z��j1��,��1����3���������1      �3�}��q�W�����ti�7�t�6��~8z�^�@�(��ĉq����1�\UU���ى�G�MQ1�RǨŉ'�СC�c       gXXX�|0u�ZL&��L&�c@'��N�٥9�=
����i�J�P��,;u�>���      ����#���B7�U��8f�Y��)��0��H���{o9r$u�a���~����.�,�Μ$�u�ڭ��#G�ĝwޙ:      ���No4u�l�umS� �K��\����:n����1j3�͔�a��oL�µ[s]:�      ��K����d]zo)L&��L&�c�����q�=���4�fp�y��j5�N;�`	u�F������Ń>�:      p'N��Ç��Q��ݼu��f1�SǨ��?�~?u��܁�����?�����1j5���a��N]�q�=�ĕW^�:      p�~?������Q��,��aE��0u�Z�z�x衇R� J��h���s��7J���4uh��hԹr{D�n�      �&��>�^/u�Z͋�J�;�Xn����;�ꫯNh(w��<�裱�н)���\�m]�0r��Ѹ��R�       .е�^��sO��+�"F�Q��x]���Kh��S�]q���8q�D�I�C%w���8&�I�I<����      M��㏧���l6��Ӱ[ʲ����N�ۏ;���A��Ѱ.�G?����Qr�K3�L:[n߿<����c       �W�W��oN#��l�$w�].�GD<�����R� L��d7�|s�z뭩c$��g2��x<N#�}�C����:      p	{����N�Nr����r�������S� N��,]��kn8�t:M�7�;]n�}(u      ����q�W����l6Sr�PE����>�h��1��Sp.˯�گ�5�\�:FR��H���h4��d�:FR������éc       ����ǣ�>�:FR�٬��]x;EQ�p8���������?�:�
��e��z���kN����7�ɏ|�#�c       ��G�}������/�� ox��c}}=u�܁���Cy0���x���TUU��Η�#"�瞸���S�       .���j<��#�c$W�"/l3��b8������R�]��\���e���x<��h�:$5/��f��Q���<u      `�<��㱼��:FreY���F�e�:
$5�L���}�{_\}�թc -���G}4<�:F�ө��tVY����EQ����{�7n���1      �]r�С�Ї>�:F�����M���Y��(��q�YXXXp  ��܁]���O<�D�٘_�e�2]��~�^����'R�       v�G?��X]]M#����i�(P?�g{���رc�c -�����q�W��H(�m    IDAT�'Y�%n.8ۉ'��oN      �e�����8u��8ɚ�����\�~���v`�)��f0ēO>�:FV��qٱI�����F�cd���      �nO<�D��������d����h�VQ�����3|���G������;��>��Ƒ#GR���h4R �u�8&�I�(ٹ�������c       {dmm-{��1�3��bss3ʲLv����m0�o��o�����;��<��5��IQ���iW�9,,,Ŀ��"u      `�}�#���������,css3f�Y�(�+l���
�w`�=��î�y�*��5�?����}q�uץ�      ����x��'S��RUU1c<����,���؈�t�:J�����c�X�@K)��nqq1>��O������bss3&�I�(pQ���+�<���⩧�J      ��c�=W]uU�ٚL&n���f�������h:t(u��܁=q�����ߞ:F���E�QElnnڕ|��G}x      2x���g�Y�(pA��q�C���q�ȑx���S� ZL��3����ca�4�v,�h���z���ޑ#G�'�H      ��<���*��a�F#�a�5��L&��Q����~6���S� ZL��3Ǐ��z(u��Yđ��,css3��q�(���|��      :�!�f:����fE�:
���w뭷���ߟ:�r���=��O~2��ۗ:F#Xđ?��[n�x u       ��Ǐǃ>�:F#�[sJ69p�����z������RGZN��S����c4����i�R��.R�׋���o      �q��;����0�ccc��k$3?�����{衇��oN� w`�=��q�צ��(��4666b6���B��n~�.΃>h�      ����~�R�h���S���]����xꩧR� :B��s�����}.u�Ʃ�*��a�C��)�K������'S�       2�裏Ʊc�R�h��t�@6j��K��O|">�:�
�@-��x��R�h��l1�NSG�e���p�L����-�      �-�� ���/F��K�qʲ�:�,��qh�y�f2����HǏ�G}4u�C܁�����b}}=u�F��*F�Qlllح̮�N�n����o�|��c       ������GI���Ed���l��|�~?���/E��O�w�6������~6u�F�?tonnz��E1�|p�A|�_p�      pN���g�ȑ#�c4�d2q�=�l�����<�?�x���H�w�V>�`�u�]�c4޼�l�2�����O|"����1      �L��������1o~����fE�:1��V��w���������1�Rpj��/~1VVVR�h����;o�,��Fv$n�)�x��1      ���{����'u�V(�"677�y[��T�f�z������˩� �����O|��c�FUU;v�z@'b�U[�k�=�^/���/D��O      h��/�e���������l6�����Fn��E?�p�y睩c ��$�|$n����1Ze{��K�5�98}����=��c��-�ܒ:      ����~���c�μ�>�;l~b����w�����g>�:�a
�@�կ~5VVVRGi��gW.uGY���{��믏O~�c       ���ǉ'R�h������Љ�2/�;�}o�z�����_�}HJ�H�k���oUU��$N�>큾Ŋ���p���=6�_�j,--��      4З���8|�p��5��bss3677c:����Ѓ�χ?����{S� :N�H�7~�7�R���+��Xn��t��8��f��ާ?��8~�x�      @C���Ǘ�����z���ZQ1���s�}�e��(N�>��������S��T� 
�@zv)�g�c�B��ʲ��x���f�z�u�]��8u      �����x��GS���������j{�ũ��p�=�w 9��뷽(�T��٘�΁��~���O      ���ԧ>���UU�uC�w���gI�3��L�t�M�c D��;�	���9�<]�e�H�צY���	      `79!9�3oM��f�#olB�L&6!$v��w�o��o���E��Ƨ>�)� �~=��{eY�d2������ܴhK�7~�7���~w�      @�\����O:u�N�N�1�����?�;���K������/���@V܁l������ƾ}�RG��e�y�Z�}o�Oj�o,���[g������}.u      ��~�73x���1:�̢�h4R��#��֛��6ddaa!�����SG�A��ʵ�^_��W��ș����◦����f1�����6dh����}͕�      ����z�/})n���Q��3���_��(b2��(��@��O}�Sq�]w��pw ;�~���c�X��CY�;v.�C��0�$0_��ØN�6	d����W���8z�h�(      @˭���׾�57�g���s���@��wf�dss3��R{�N�8�?�x� ��d驧��{�'u�c6�m-�/L����/r�;�O�:���ۂ-��;�w�}w�      @G��ʲ��d�U���؈�h��Ӈ����hk#�h4�to�)�;f����di~���W_�:
h{�{�N����(��-^����l�c�frs�8q"�|���1      ��q�}��O*���1�Lb6����^EL�ӭ���������f~{���j�( oi1u ����������������x<N�KP��gnaa����в,���(�2ʲ��(���v���k��_�r�?�      @{=��S�?{�[u}�q�}zzhK)�(�\,:'�8��:aUG�^�/���˦Y�e���0˲���[\�9�˜��\�]�2oh�:e����Ѡc
J�|�>��I�����<���?�x<��C����8 ��7��z�P(t5�b�-?�jG��yG!^�=
�B�{�q������@�ƌg�yf|�+_I=���.|v��w<�걷l߾��;_��x�w�����/�8���z
      �G
�X�ti,_�<^x��s��o߾˃#����6bo6��#v�$v4����Ν����g �+�;����:*�y晸�[RO����~w\������{�3}[YYY,[��7�     ��jjj�K.��.�,6mڔz�h���ݼ=t�Fb�B���&O����'R� �-���`',�����3��ۿE����q̮,^�8�L��z      @DDp�q��G�TJ=�L��G�N#����G��رc���Ϗ�2�(�3x�z�B�K�,�C9$������9s椞      �|p�{u7s�w3dȐX�reTTT�����@�Q^^\pA����� =\kkk,X� �      �]:��#���x�@׿�X�bE��֦��G�@�RSS�^z�]�{����w��      ��͟??���S� z�b�]tQ�5*��=&pz����X�b��� {��      �S
�X�dIL�0!������tw�Gjjj�O��QV�m�=����       �(�b1.��B'0{�SNq�GS�=ִi���sύB��z
�������Kc���O=      `�TWWǪU�bĈ�� =�q����K=�}�=Z{{{�q��g �����.�,<���S       ޓ��ڸ���c�С�� �3gN,Z�(���M��x�g���إ~�����ˣ��)�      �����>V�Zuuu�� joo��O?=���B��
�w\�x≩g )//�/�0>����      �W444��ի���6� #�Їbɒ%Q(RO�+�@�q��'�G?���3�����ҥKcҤI��       �UÇ��.�,���SO2p衇�g>�(��� �5w�W9��Sc֬Y�g 	����y�ӧOO=      �[�3&V�\UUU�� 	M�0!�/_�R)���J��*�B!�:�8���SO(�q�y�E[[[�)       �j���q�WDMMM�)@�vX�X�B��Jw��)
��O~2.\�z
��J������      @�1v�ظ��+���.�`�2eJ|����~�����-�@����)r�>���"V�X�~x�)       ��ȑ#c���Q__�z
�y�q�E9����@����g�uV
��S�nҿ���ˢ��%�      �$�k׮�����S�nt��ƲeˢX,��Э�@�w��Ƨ?�i������/�<���SO      HjȐ!�v��5jT�)@7�;wn�y����;�'����ҥK���<�`/�����k�FSSS�)       Y����U�VŘ1cRO��SN9%N=�Tq;�g܁>�#��K/�4���SOާQ�F��W_#G�L=       +����v�ژ4iR�)��T,��ώ��㩧 �Sw�O9�C⪫��!C����G---�v��<xp�)       Y�����˗��ٳSOޣ���X�|y̚5+��}N��9p@\}����Ԕz
��>���%�\���O=       keeeq�g��ŋ�P(���A�Ś5k��K= 	�;�'��~�z��:uj�)�n(
q�I'Ź��b1�      ����#.����ׯ_�)�n=zt\}��1f̘�S ��}VEEE\t�E��ёz
�J�R,]�4�ϟ�z
      @�4mڴ��+b����� �`�ĉ�v�ڨ��O= )�;Ч�����ŋ���Ow*4d���6V�Z3f�H=      �G7n\\u�U1bĈ�S�]8��b�ʕQUU�z
@rw����G>�W������S������\sM477��      �+���q��Fkkk�)��+�Jq�y�ŢE���L�	!p�����]w]�?>���9����>C�I=      �W������??/^�n��ذa���k����:*����vRWWW^yetvv��}R�T�O}�Sq�9�Dyyy�9       �R�P����X�jU��֦�}ҤI���k��Q�F����;����X�pa,[�,***Rρ>���>֬Y3g�L=      �O8����뮋�:(��3
�BtvvƊ+���:��,	���3f�ڵkc�С��@�7q�����MMM��       �)���q�W��G�z
�z��+W��P(���-�;�;8����믏����S�W*�q�I'�%�\555��       �I�R)�,Y^xa0 ��ƍ�]w]v�a�� d�<� ��UUU�ҥKcʔ)q�7ƦM�RO�^aĈ�lٲhllL=      ���6mZ455ŗ�������z�
�b1�͛'�xb��9�`w�vSkkkt�A.�`/hkk���>;***RO      `'��իWǏ����7�o��f�I�c:4�-[�ǏO=�G�����W\��v[|��ߍ�[���=JMMM,Y�$�N��z
       �C�P����?~||�K_�g�}6�$�q���⬳Ί����S z�� �Ceee���k֬�����s��8��C�n�      �cǎ����q��G��=FMMM\t�E�t�Rq;�{�w��hܸqq�7�~�����b۶m�'A����'�|r|�#�B��z       {���2�,YӦM������/��ٚ<yr�}��1hР�S z4�;��PQQ.�#�8"��կ�c�=�zde���q�YgE}}}�)       ��vX|�_t �B]]]�~��1mڴ�S z�;�^0f̘������o��o�9�lْz$��~��g���      ��q`kkk|�k_��<�$H�P(�̙3��N�����s z�;�^R,�����"��GM=	��B�3f̈ŋǀR�      �466�5�\� @��aÆ�9��rH�) ���`/khh�U�V�]w���ַbӦM�'�>1bĈ8�����N=      �n�� ��S�ƍ7���_RO�}�T*�ܹsc޼yQ*�R��� ݠP(ĬY�b���q��7�O~�غuk�Y�-������3�?��(/��      �/1bD�Y�&x���馛���O=	���ɓc�����Аz
@��B�F��ձx��={v|�߈?���'�^S(bƌq�i�Emmm�9       $4eʔhii�;�3~���믿�z�5#F��E��ĉSO�� �����c�ʕ����M7�O?�t�I�r�!�hѢ=zt�)       d�_�~������q��7����ؾ}{�Y�0 N:餘3gN������g�����������'?�I|�{ߋ�^{-�$�#Æ�Dkkk�)       d���.�9�8�c⦛n�u�֥�{�X,��ٳc���Q]]�z@�#p�Ǌ�btttđG��rK���?�͛7���hРA1o޼�9sf����       ��;vl�]�6~����7���d���,f̘'�tR444���g)� 8p`�v�i�����~{�y���o��oQSS��G���#���z       =L�P���֘6mZ��7���|�;��Ϧ�oQ(bڴiq��'ǈ#R���� �80.\s�̉�n�-~���Ŗ-[RϢ�����9s��	'�UUU��       �ý=t�����=�\�Y---qꩧƁ�z
 �O������X�xq�p�	���0��غuk�Y�1UUU1{�����>���O=      �^fG�~��ǯ~������6lH=�>���%,XcǎM=���df���q�9�Dggg�q�q�=���͛SϢ�4hPtttĬY���       t�b����1}����/w�qG<��өg����hmm�N8!S���d���!�8���'>���/��[o��^z)�,z�ѣGǜ9s���=J�R�9       �1�R)fΜG}t<��#q�wƃ>�z�Leee}��q���ǐ!CR��]�2׿����c�=6�ﾸ��[c����g��577�ܹsc���Q(R�      ��+
���---��O�����w_lݺ5�4z����8��c���#�z �I��C���G{{{����C=w�qG<�裱}�����!J�RL�>=N8�=zt�9       �Kcƌ��K��)��w�yg�s�=�iӦԳ�A<��8���#���r�$@O���)
1iҤ�4iR<��s��_�2���x��SO#S#F����:*fΜ555��       �n2dH|򓟌�<w�uW<��#d����b�ԩ���---�� �>�z�aÆ������O�G}4�����~��\D�T�)S��1��      ��T*Ekkk���Ƴ�>w�}w�s�=��+���Fc֬Yq�GFeee�9 �w�^���,ZZZ���%^~����{�?�i�������566F{{{���ŀR�      ��j�������'�������{z(�mۖz�P���c���1{��3fL�9 �ew�^���.:;;c�ܹ�nݺ�����׿�u���L=�n2t�И>}z�����z       t����S�_|����o���[�.�oߞzݠ_�~1ahmm�iӦEEEE�I t�;@/U(���9���cѢE]��}���]���!Cb�ԩ�����ͩ�       @2��������#~��߉�{�R�---�v�>F�����v�i��#��}��<�@��_�J=�������������s        ;��ݟ{������<������***b�ĉ1}���<y�����1�b1&N�'N�m۶�O<?�p<�������R���b	���"j      �=0lذ�7o^̛7/^y����>�`<��ñiӦ���ICCˈ�    IDATCL�0!&O��zh�J�ԓ HH�Ї���Eccc466Fggglܸ1}�Ѯ���_N=���q����'N����ԓ       �ǫ������hoo�:���|0�q�c1~���<yrL�:5��z �Х��&Z[[���5�o�����O�S����u���ƍSO�ub���]'�744��       ���Ο??^~��x�G������������8蠃���9>��Dsss����5�! إB�MMM���s�΍��6�_��׮�3�<�n������ã��9�������d       H���.��ڢ��-""^���������[�.6oޜxe�RWW���]�DSS�����7 ����!���=""^}��X�n]<���~��x�'bÆ���(//��#GƨQ�bԨQ1v��hjj������       �wPUU---���[�n�������c�œO>O>�d�_�>���'^����w�cƌ��������S����80�N�S�N�zm��ͱ~��x��'㩧����z*�|��ظqc¥ݧP(�ׅ�ȑ#c���Q,S�       ާb��ƍ�q��u��}��x��������b۶m	�v����9rd�=���=ztTWW��@/#p`��������hjjz��[�l��^z)6l��?�|lذ����s��k���h񻫮��:����.���~>|xTVV��       �C�B��8��û^ߺuk������/�����J��������Q__1t����$��B!�L � �; �D�T꺰ە�7�+�����j��_���7ƫ��7n��7v��y��x���#�?��oٲ%""6mڴ��X,v蕕�Q^��_}���QYY��FMMM80555]�A�EEE����        z�b���766�ן�8 pG���x���^��_=�m�۶m�:8��7��j%ޮ��*��ʢX,FUUUD���������&bG/��QWW�}�1 �� da�����e˖x�7�.�        r�n��۷�k���������Ы�J�(�J�g        t�B���թg @�p�-           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;           Y�          ��;        �;wl���a�Ҷ�`;�J7i2@jO`��(#p�c���OPa�y��<|�_�� ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @���������          ����s���          ��	��yxx�         �
	��y~~�         �
	������fo           NO�N��          �I�N������          ��	��clgo          8gc�����;9�����          ����#p         8:�I��3����          p��w���1|p         ���3Ƹ��         ����N������          ���S�c�1{         �����$�;5���         �U�r}}}5{          0�����~�a�         �s7���� ���r8�          �RwR...���           �!p'e��v�          `�;)w          X/�;5w         ���� ����;          �����;          �����         `���lf           ��          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          ��n� �o����,���;~����ǻ���3          ��n���,���;~�����o�Gp\�c���l����Wl�����f�         �5�{Y�/�G���p|of           �e�          !p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w       ��{�    IDAT    �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�         ����@A�?eI��>��gQ��0 � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p       ���  ��;       �����  ��;       ��;  �N�  p�    �7�;  �N�  pp]��    ���   ;�;  ��}��    ���  ��   ��LO     >N�  ��          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;         ���;�n[I(���-��$�|U��O%��� ��@�w�  U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;           U�          P�;  �o\���+        ,��  �7��}�        E�  ��ݮ�
        �"p  x�f�I�0�^       `Q�   o���G�        G�  ��8�i�Z�^       `q�   �<==�qK�       �8w  �W~��Qz       �E�  ��m۴��K�    ,Dι�
   U�  ��Ǐ>(    a�q,�  @U�   ��sN?�,�    � �0�^  �*w  �����m��k     2M�wI  �_�  �����
    ������s�5   �!p  H>"    �x�  �/�;  @J�i�t��J�    ,��pH�˥�   U�  ��~��Yz    `����J�   P�;  �x9�Z�J�    ,��  �_�  ������}�5    �;���t:�^  �8�;  �x.#    5�V	   p  nǴZ�J�    ����Rι�   E	� �E[�Vi��k     ��m��x,�  @W��    IDATQw  `ў��K�     �?�,�  @Qw  `��qL����     ��(  �tw  `�����4M��     �������)�  @1w  `����J�     �?�]  K&p  �����nK�    �?���Sι�   E� �E�    �U��i�ٔ^  ��;  �H��ϥW     ������+   !p  ����4M�5     ~����_( �E�  ��^�}    ���}��v��   'p  ǯ}   �9�	  ,��  X�q�f�)�    �_�V+�  G�  ,�f�I�8�^    �ڶM���   ��  ����/    0'�4 ���  ��sN�ժ�     ��M  X�;  �MӤaJ�    �n��)].��k   ��  ����\z    �{yy)�  @�;  �9�^�K�    �aw  `I�  �"��u]�5     >��&  �$w  `���K�     �)9�Z�J�  B�  ,��?    ������^   ��  xx��)].��k     |Z�4����k   ܝ�  xx.    s�sN����   w'p  �j�*�    ��9�  ,��  xh��-���k     |�f�I�4�^  ��  �C[�V)�\z    �/�1�v��k   ܕ�  xh�ͦ�
     �f�^�^  ��  ���9�   ��"p  ��  xXMӤaJ�    �m��sj۶�   w#p  ���    �#r�  xdw  �a�V��+     |;�;  ���  �Cj�6����k     |��v��q,�  �]� ���    �iJMӔ^  �.�  �C�    ��(  ��  ��q�    xt�ժ�
   w!p  �v�M�8�^    �n��K���   �N�  <��    ��[(  ���  ���Q    Xo�  �#�  �|>��mK�    pwMӤ��K�  ��  �CY�V�W     �sNMӔ^  �[	� ����nK�     f�ٔ^  �[	� ��1MS��v��     #p  ��  x��.��Xz    �0mۦ�mK�  �m�  ���n��W     �m  x$w  �a��    ,��Q  ��� ��0C:��     ��lJ�   �m�  �Ch�&�K�    ���t<K�  �-�  �Cp�    X��v[z  �o!p  ��7    ��y#  ��  �������s�5     �i�&M�Tz  �/�  ��2    �t�8��~_z  �/�  ���lJ�     P�c   �#�  ��4M�     ��  �@�  ���|N]ו^    ���~��q,�  ��� �Ys�    �_r��L ���  ���lJ�     P�;  0ww  `֚�)�    @5�  ��	� ��:�i��k     T�|>���K�  �iw  `�v�]�     ��s�v
  ̚�  �-i     ���S  `��  �l5MSz    ��x;  �L�  �R۶�z��^    �:��!��Xz  �O�  ��    ��r��p8�^  �S�  �,�v��+     Tˑ  `��  �,�8    �{�P ���  �s����r)�    @���}�9�^  ���  ���v��+     Tm�t<K�  �aw  `v�Z    �Ｅ  s$p  f�G    ���7L  `��  ����N�S�5     ��4M�9�^  �C�  ���     �>}ߧ��Rz  ��  ��K���6    ���)�  ��� �Y��W�U�,    �{�|S  �w  `6r�i�߇�[��a�     �!�M  �;� ��8�i���y.�    s׶m����   �&p  f�p8���.�ǰy     ��s}[  �*�;  0������g�,    �{�|[  �*�;  0�a����f    ܓ�  ��;  0�0���6O�    <��~�rΥ�   x�;  0��!l�0i�ل�    ����S�u��   x�;  0���]��i���y     ���
  �w  `"/������    � p  �B�  �B�Ǘ�j6     B�  ���  ��.]�װy.�    ��p8�i�J�  �Ww  �z�����K��1l    @�i���t*�  �_	� ������Y��    ����yL  ��  @�"?��   �H]ׅ͊<&  �Yw  �z.�    ��z����  s p  �v:��8�a���u�,    ���6�r������  |��  ���p����C    p�^�0!�r��x<��  �,�;  P�ȏ-///a�     ��g�ȣ"   �!p  ���V��Y     ��<�q:��f  |��  �V��r]p    J�|��|s  ��;  P����0!��iJ��&d    ��"�����i
�  �Qw  �Z��!l�f�I�8��    ���tJmۆ��9���2  �3�  @�"?��V��Y     �E�Q�ǰY   %p  ���e�݆�    xm�ل��  5�  �:a���u�,    ��"�ȿg  |��  �R���z����9��iBf    �%2p?)�6  �#�  @�"����S��a�     ^;a��8���Bf  |��  �Rd�y	    �-9��n����Y   !p  �$p    �&��t:��  ��;  P%�;    �4�o��o�   !p  �3MS:��a��    @"�*�C�,  ���  �9�N)�2�m�t�\Bf    ��v�{�^�����Y   !p  �s:��f���Y     2C���a��c�,  ���  Չ����_    ���<�!p  j$p  �s>��f	�   ��l�۰Y��%l  �{	� ��N��Yw    �&��#�b  �K�  Te�t��BfÐ��}�,    ���<�!p  j$p  �r<S�9d�f�	�    �mۦ��2k���#   �%p  ���&����	�    �^��6l��|�  �w  �*����    5��va�"�d  �C�  T%�Z��    �Q�ۥ�  @m�  @U"?�D^A    x�ȷK�;  P�;  P�i�R۶!�����]    �J.�  K&p  ��z;    @J]ץ��Bf]��4C�,  ���  Ո�#/     |�+�  �R	� �j�N��Y.�    5�  K%p  ��E�    �,�3��  ��� �jD�׏     >*2pw�  ���  �B�9�m2k��t<Cf    |F��;  P�;  P��咦i
�����f    |��|N��-dV۶iǐY   #p  �y!(�׾     ���y�\�f  ���  �B۶a�"�    �Y��{�-  ��� �*D^r�    ���c.�  ��  Up�    ���|�t�  ���  �B�u��s���!�     �"�o�.�  ��  ��S�u!���s�1d    �W�N�4MS�,� �Z� ��ڶM9�Y��!d    �WMӔN�SȬ�m�bz  �?�  �E��V�    �I�fԟ6  �D�  ��[�;    0'�o���H   ~G�  �;    ��"�4#��   ���  (�w    ����  ,��  (N�    �6� ���  E��>�t]�n�[�,    ��p<�f��  �@�  u���8�!�\o    ����#!.�  5�  EE^�    s��9MS�.d  ��� ��"/	�   �9�|�t�  (M�  �;    ��E�mF��  �E�  ��[�;    0G.�  K"p  ��    �Y��f�-  �[�  @QQ׀�a�k]    `�"���6  �-w  ����2��v    `�ڶM}߇�r�  (M�  s�^�4M!�N�S�    �{�z��.�Cf  �E�  y	H�    �Y��4Ma��  �"p  ��^�a���s�,    �����v  ��  (&��    ��ȿTF��  �&p  ���H��    �E��  %	� �b"s�;    0gw  `)�  @1�I�    ��E��2�8	  �kw  ����$]ץaBf    �Cd��;  P��  (&*p���    p�0�  (E�  q�^�4M!���s�    �{�z�^�)�2  �5�;  PDԥ���    �c��[�4M����Y   �	� �"ڶ���    ��"�yt]6  �Ww  ��    >F�  ,��  ("���    x���<R  �+�;  P��v���    �^"�y� �R�  @}߇�r�    x��<"��   �J�  u���4�c�,    �{�<�y�  �Ww  ����?mۆ�    ��a��s� �R�  @����    ���<���	  ��  7C�9���    ��뺐9Q��  ^�  �"m+p    Iԛ�0i���Y   ��  �"��kF     "�z\�װY   ��  �"���6    ��"�ȷ\  �� �p.�    |Nd���}�,  �� �p��{��    �{�<��;  P��  'p    ���7O�;  P�� ���{����|�W���{��$#~#0�pg��ď8 ;�hG�t{D�6����A EY8�D�����ǀ�G� ����%aǱa+�*�%����5�uomb�5�]��VW�]U�j�����H'�    p2�3�/~�i�   ^'�  ��
�ƽ{�Rj    d����  mp  �e�]o    ��k��MӤ��|�  �u�  @:w    ��i�&^{�Z�  @� �Tu]�h4J�%�    ̣�٧�;  �w   ս{�Ҟ�p    �Q��{���  x#w   ���aZ��%    @���u]G]�)�   ^'�  �p    �L��3s�  !�  $�|���ݻi�     �d�>3g�   �  @��k?�    �<p  晀;  �*3���/~1�    @����h4J�  !�  $s�    `2.�  �L�  H��p    �Q��3�h	  @��;  �,s��L/    @��٧�;  �M�  H��q�    �G����W9  "� �dYː��è�:�    @&� �y&�  ��Z�d.x     2e^pp  �	�  ���!�    �Lu]��Z�^�  x��;  �J�    `rY�X�F��:   �p  Re]��Z�     �!�ȇ�  @6w   M]�Q�uJ-�   �y�u�#�UN  ��	�  i2!�    �<s�  �W�  @��h�V+�z    @��u]G�4)�   "� �D�wW�    �y���e�l  @�  HS�uZ���ôZ     �2g���]   w   M�w    `�e�@]p  2	�  i�    ��w  `^	�  i�    �#s��;  �I�  H�y�G�    �g�3Pw   ��;  �&3�n�    �3w  `^	�  i2� .�    �,s�y�  @�  H#�    0��Vw   ��;  �&s	"�    �3� �y%�  ��\�d^/    Ȗp7o  2	�  i2� .�    �L�  �W�  @w    ��p  敀;  �&k	R�u�u�R    ��w�V   ��;  �&k	�z;    0�2����  dp  �d�-[    �y�y���  �$�  ��Z���    ̻�hMӤ��:^  !�  �!ׄ    �� k��  �p  e-A,[    ���,  �G�  @w    ��1s  摀;  �&k	R�uJ    �6e�B� �L�  @ׄ     ���  �G�  @�    ��1  摀;  �&kْ�,/    @��\ �y$�  �q�    `z���f�  @&w  `�X�     �Y(  0�� �4.�    L��+  0�� �4�-     ӓ5��:�  @��;  �Ȳ    `z�B �y$�  �q�    `z�\ �y$�  ��l    �3W  `	�  i,[     ����:f�  @&w   M�$k�    �&GE  �y$�  ��    �<p  摀;        o�(��[   �w   M��,��    �?�s  `I}   i��-�:    �y�  0��  �p    ���๙+  �I�  �;�-    �y`
  �#w   ��     �c�
  �#w   M�$�Y^    �6e�B�\ �L�  �kB    �y`
  �#w   ��r    ���  �G�  @��%��r   �� k*�  d��   Ҹ&    0=f�  �<p  ��    L��+  0�� �4�-     �S�9�3W   ��;  �F�    `z�\ �y$�  ��Z�d]-    h��;  0��>  ��c�    ��  �<p  �X�     L��+  0�� �4e��'H��M�    Ц�Y��;  �I�  H�p�t:)u     ڒy���  �$�  ��Z���    ̻��y��  �w   ��;    �t��  �+w   M֕��(\    暀;  0�$>  �4�KW�   �y�9uP  ��/   M�D�    �g�E\p  2	�  i\p    �� �y�/   ��;    �t�  ��_   @��%��;    0�2g���K   � �4�w    `�	�  �J�  H��q�    �g�3���%   �  ��    LG��w   ��;  �&�ʏ�;    0�2g��  @&w   ��B     �!�  �+w   ��     ӑ:Ϝ�  �  H��p��zi�     �e�@� �L�  �d���~Z-    �lY3Т(Rg�   �  @w    ��)u�� �l�  @��'s��;     m�:�9�  �p  �e-C\p    �Y�����  x��;  �*�9[w    `�e�b)�  dp  R��    09� �y%�  ��Z�d]/    ���v�^��:Z  �:w   ��;    �d2_�t�  �&�  �ʺ�S�e�#    �L�  �<p  Re.C\q    �Q��S�  �&�  ��\�d^1    Ȓ9��z�  �u�  @*w    ��d�>]p  �	�  �2�!���    dɜ}
�  �� �T��ٺ�    ̣��g�L   B�  H�y�G�    �G��O� �l�  @��eH�3�     Y� �y&�  ��|�V�    �G)u��p  �	�  �2�!���i�     �d�>;�NE�R  �u�  @�^���p    �Q��3�EN  ��	�  鲖"�    �<ʚ}����:   o$�  �)u�   �yS�eڌU�  h��;  �.k)"�    ̛̹gV�  ��� �tY��KF     2�^/�  ��� �t���N��i�f��     |���!N����9�  x��;  �.��O�    �e^pp  � �  �;+�#\q    N�qg��  ��p  �	�    p  �R�  @�T$    IDAT��`�V+s�    p�� �y'�  �s�    ��qg���ɗ*�"z�^J-  �7p  ҝ��;    �,ɚy�z�(�"�  �	�  �ʲ�n��R�w    `�d�3�   ���;  Њ��m���    � �  �;w  �Yˑ������;    0+��~t:��Z   mp  Z�����]�p    f���rZ-w  �-�  @+2�#�K    �Ӳ���VK�  h��;  Њ�`�Vkҥ�+�    �,�<�9�  x#w  �i�\p    �A���.  �	�  �ȼ�3i��w    `��  ��  @+2��Lz�H�    8-Ǚ?f�]p  �"�  �"s9���    W]������<���v����  �r�  @+2$.�    �踳Ǭc��  mp  Z��$�t�#�    �����A�z�S��>w  �M�  @kS�������)�     �U��؟ͺ�!�  �K�  hMf�|���    �i8��qee�;�R�  @�� ��d.I&�n$�    L۬^pi�   ���;  К��ŴZ�^7p    ��8s�̀��  @�� ��d^�\�     ��8�I�x��;  �&w  �5�K�I�.�    �V��؟��g'  �r�  @k2�$�.�   �i;��qii�;����E��I�  ���  ��v���vSj	�    ��i�c��.�g��	  ���  ��Z����EQ)�     �8�����c!�  @�� �V��:eY�����;    0Mu]��ٵ��S��Ke�l  ތ�;  Ъ��ŴZ�.���   �i�Հ��  @�� �V���;    ���F�lsii)�  �W#�  ��,�]p    �eV/�g�l  �w  �U�׀�   �Y1��� ��	�  �r�    8�f�{�׋^��R  ���  ��v����Sj	�    �b܀{�ߏ�`p��q�  ��  @떖�R����XXX8���   �iw޸��~ʝܗ5�  �Z� ��e^r�    h۸��#&�i��  �,p  Z'�    �'�pw�  ��  @�2�&��     ��fV�.�  �@�  h��    �yr������)v�\p  f��;  к�t�]�    ��,^p/�2��~J-  ��E�  h]�ߏN��RK�    h۸s�N���˧�͑���(�"�  ��"�  ̄��Ŕ:KKK���N�}w    `R�^p_[[K�g�h  D�  �	KKKi����D�r    &1n�}�Y�qd�h  �w  `&d^p    �2n�="bcc�;�R.�  �B�  �	�ׁ2�B     ot����  �y$�  ̄���    @[f����;  0+� ������Vkҥ��;    pR�܋�����S��HY�����R  �A� ��0����Z]]�N�s���    '5n�}uu5mf���EQ��  xw  `f�����)�r��G�    �I�p����}�/l  <��;  03����jM�w	    �F��766N���� �Y"�  ̌���/�\q    ��i��g���3g�   "�  ̌�+A�.��   ���Fc�w  �p  fF��w     []�c6�{Q����R  `�  ��X\\�N��Rk}}=��8���   ��7ྼ��~���9���e)>  ��   3eii)�N�Ӊ��Չ~C�    8�q�Y��#r_�  ��;  0S2�)}_�    8�q��.�C�  �5�  �LYYYI�%�    dr�  ��� ������Vk�%��;    0���Ǟ)��  �g�  �Lɼྵ�5���   �q�{�="bss�;�R�  ��p  f���R�eΟ*�p    �5n�}uu5��)wsdqq1:�NJ-  �q	�  3�(�X\\L�U���O�
�    ��Fc}nҗ'���v  `	�  3gee%�֤�"w    `�^p��g�b  �%�  ̜̫A�    @�  �#�  ̜��մZ�    �ik�f�Ybf�=s  0.w  `�d.U.\�0���   ���z�������hY�.�  3I�  �9��vSjM�0:��%    �|�Fc}.�z���r���  0{��  ̜�(R��O�4p    ��q/�g�3g�   �!�  �$w    `^�������Z   �!�  �$w    `^�b��w  `V	�  3I�    �Mӌ5C,�2666::"�  �*w  `&-//GY��ɲ�������p    �̸�ۇ�at:�S�����b�z��Z   �%�  ̤�,cyy9�ޤW�뺞R'    �<wvx�S�侕���Z   �%�  ̬�'r'���    |5�^p���<�N�˜�  ��;  0�2�	�    �a܀��3��p  f��;  0�2�,�>�+�    |5u]����/�r'�	�  �L�  �Y���QEJ�������'���;    ���kv8'�OG�Ӊ����Z   '!�  ̬^���h)�b�+��^b    ·qg��.]:�N�[[[K;,  p�  �L[YYI�5��w    ��F��X��������  8	w  `�e.[.^�8���   �77�>�l�82��   ���;  0�����jMz%i��   ��a��{�Ӊ����n�d�\  NB�  �i���i����ciii��p�    �8��s�Q�9�N��;  0�� �����cqq1�ޤW��   ���GD\�x�;�omm-��H�  p�  ���|2W�    ��q��$�#��L  ��p  f�Y
����0    0�f1��9k  8)w  `�e^�x��DO���    D�p��s� ��@�  �ykkk�Ώ����p8��7��   �|k�f��3�����XXXH�  pR�  ���t:����V��ŋ}��    0�Ɲf�]o  �
w  �L�\�L�Tr�    η�h4���  �R��8=��6:���u��t:m�  Y[[K�%�    L���p��M���qd�X �4MSTU��˲|�ڵk���~8�s���ۏ�u�?�M�|��  `R�˗����v�c/��\�4�4ME1��    ��`��kkk�����MDQ�  ̅�=8�o��骪~�(��k׮}�(
��戀��x����޽�]EQ�x]���v?  0m+++��t�~�weYƅ�3��̉C�    Χ�i���~����	�YZZ�^��V  �#��i����_�n������g�y�ϵ��p?�����1"�q��ݧ"b�o�e
  ̝�/�Իz���w    ���HǕ+WN�������j @��(���z�UU�N]��~����''�~ݹs�pp�=��4��"�YH  ΅̀��˥�����L�    �7�~���S�侵���Z  Т��x�,�ǫ�z!"���'�|���8�3��۾w���������  �����'>�R����Qŉ/���    ��8�����	�q� �s�ш����/����_���?^�~���n���ϸ7n����om�f����{����  �V敡~�[[[���~�ĿQ�u�e9Ů    �Y7N�}�$��,�XYYI�  3f="v˲ܭ�ꅦinE�{{{��n�7',=�>��^*��_E��4�׵�  ̂������q��ݔzW�\�(��;    �/M�D]��\f�}mm�!  8�hQ��������ht����/��_I�}�ܾ}�Ѻ�w#����v?  0k��a���K)��\���'�����t:S�    �e���c}��ի���}���i�  ����4ͻ˲|WUU�������x�'�)�g�͛7����E��u][��  �,���H�O�dr�    Η���y�^�[[[	����H�  gL�E�cQUճu]����9�ޔ�{�nݺ��EQ�E�;"b��~  �,�i�c}}=��/��ĿQ׵�   ��'�~��崙aQ.� �xv"�˲����~�(��k׮}�(
��Z ����͛��`���G��  8�����v�c?�;�+W�Lpw�    Ώq�W�\I�����R����z  0��x�4�����֭[�w���O=���m7v��'y��g���맚������v?  pVE��0>��ϦԻz�j|�#9��뺎N�3Ŏ    �Y4��:x�p���H�  s蛊�x�h4�QUկ�u��ׯ_����:�Oѝ;w:����?����G��?����  `d�']6��    ��8�N�e�.]J���p8L�  sl!"�^��۫�z!"�#����>�r_sK��TUu�i�'���\;  LS�Rfmm-�����W_=�o�ueYN�+    `֌F�~��ŋ���E5\p ��{4"��xoUU�V�����?i��y#�>%7n�(�����4�nD|oQ�� �)Y__��,���zW�\��}�c'��+�    0��	�O�b�q,,,���BZ=  8g�#b�i�kUU}(�������޽���B�z���w��}""~�i�om�  8ʲ����x�WR�Mp��::��;    fI]�c�z�jB7G\o �ED<��������/6M󁽽���r_g���	ݾ}�Ѻ�w�޽����v?  p��ô���K'�   `��s�="���˧��}��0�  W��ywD����7Mssoo�E!4pL����sϭ~D\������  γ���x���j-,,�k��v�ߨ�:ʲ�bW    ��8<<|�g���b0$ts�w  hM�E�����Goݺ�lQ����}����
�1TU��EQ�����nD�  f�p8��(R��E������Ŀ�;    ̯q.����$tr������rZ=  �M}}Q���귋������ݶ��u�o�Ν;����݈x[�4E�=  �u��XYY����N����3Q�����t:S�    �M��\�}8��  �2��Ǜ�y���?-���w��sO?��ߴ��,p�2UU���(��#".��  ���aj�}M�D�4Q��,    ̓q��eY�իW�9���qz  �a��4��v�����_m��?��?�?�nj��Gč7����6M���ig ����O~2����Z���N�p   ��sxx���\�|9�ݼ���;  �	��[�nUU/D������K?��?���k۹�������t~�(��MӼ��~  �����L�����gv���ueYN�#    �m��'}!�8:�N�����  ��ш�����]UU�8����w���m7Ֆsp���DďE�?��^��   '���cii)>��ϧ���ޞ(��4��    ��4M�F�~.3�>�$	  g�0"~���<SUՇ#b�ӟ���q�ƃ�e�97����#�EĿ����r;  ��lnn��']B5MM�X.   ��'������ŋ	��~�  8eD<�]�z�S����t�޽�?��ӟl��sp�}���u]�F�D�r��   ӵ�����Rkqq1677��_>�o�u�Ng�]    m9<|�ŝ��(�2��#�  0w���yw���W�n��oeY��ڵk*�bn���ˀ���?�p���������  pz666R�=��Cܛfn��   �sg�����	���z����V  H�)��;��������}�֭��}�g>�vc�6W����o��wܽ{�ZD�'�  p�z�X[[�����J�����Gt���u=�n    �6�p���I�����fE�V  h�7E�^�w����)�bww�w�njZ�|��Ν;����ݦi��R �sfss35�^��DA���S�$    ������/6.--��B���   �3�x�4�WU�BD�/..�ʓO>�jۍM���?���E��D�Cm�  �gss3^|�ŔZ�n7.]����gN�Zz    �������y��8��;  �k�FD��/|��WU��#�?����϶�:�3p�q�F����֦iv#�{��  ������������D������L�#     �8����N�,,,���RZ=  `f�E�nD�VU�B�47���ս��{m76�3�}����h��EQ�5M�um�  ̖�,c8��/��Rogg'^x��w    8ۚ���h������$tsdkk+�  pf<Z�/D�{���~4ݺ~���m7� 3p�}���u]��u���(��  �]���i�K�.E�׋{�N���뺎�,��    �e�p�p8����n�lnn��  Μ�MӼ�,�wUU��������'�x��ܴ`��7o�\�O�u�mm�  ��˛�,cgg'^|�����;    �]������?��ɑ�(� �q��XD<vpp�UU=[���_��Rۍ���ܫ��{��<"VZn  8c��֢�펵X���~x�;    p6�Z�}yy9��~Z=  `.�D�O�e�SUU�VQ�׮]�PQMۍ�p�y��`0|wD��ѿ   8��/��R�?*~�[���{�7�o��    gO�41���g��n\�z5�������Z  ���G��M�<�����[�n=��vo?��S/��P+�[�n}CY�?�4͏Dą6z   �Of�}ii)����s��܉�iZ�G�    �1�s�����N���͑��ʹZ  �\���(�3�nTU��u]������ ������;w:/���?*���"�mM�Y� ��!{����Op��:u�    Ln����?��ɑ�(bcc#�  p.,D��˲|{UU/D�~D������3��z�����M�<ypp�΢(9�z  �������k���{�G���O���i�i�(
��    ΊY����;�  ��G#����VU�kEQ�������,x*�7n����om�f7"��(��K�  �������ԧRj]�|y�@�+�    pv�uu]��lnn���JRG�/[  ��zD�6M������MӼ/"~soo�޴M5x�����޽�DD�D�4�2��  ���VZ��(���ى�}�c'���i��    p�ƹ���#���_�p!�  @�4���������,?��SO}bZ�?����۷��z��ݻ?K��M  ���p�BE��G&
�?��    0;f-����bmm-�  ����4ͻG�ѻ���pD�oll��O<1��GOp��V�?"��u��4  0-�n7����W^I����O���:ʲ�bW    �ixP�}0ĥK�����  �eeD<�|�֭[�����{�;���N�c��WU��EQ�����nDl��(  �i�p�BZ�}aa!.^�/��҉C�    f����]<��C���.��  ��E�{���LUU�]��������
�߼ys0�;"v#�I.  ��.�G?�Ѵz�<��Dwc   ��{������E[[[i�   �i�7M�xUUZEu�޽�~��y��φoܸQ��w��t<��g�Nz#ɲ�1�Ι��<fL���YU+�h#h��Z� �hHi�5��k�4����$w7ӂU_dFҝ�A���ٹ�k<g��^� p�MNN���X�z7z�(
!w    ���gY�4�>33�z=Y=  �8.�����j�߿�˿���|m�}yy����n�5  ��,Kz5���|�����o�y~K�     ��(���z�,,,D�umN�֤<  �%G�����u����׿E��~k-  $��jޛNfp   �����\�'���w  �aʲ���_��O������?�s-"�="��{1  �-y��yT*�^Zuk666n�|QQ�-u    ܦn�{힛����l�1    IDAT���d�z   ���eٿ��O����oڣ�n�/�;i  ��U�՘��KVomm-j�ڍ��)�    p?]p�������D�\Noϲ,Y=  �[�]����~�W��򗿼β����   ����ϓժ�뱺�z��!�    �O�۽��ŭ��4�����|�z   w���_��_\���_���z�e�oD4�-  �;�rbR��_bEq�2     �릷GDloo'��R�R�gϞ%�  pG�,�������|�	����%  �;6>>�����mnnF�r�EYC3�    �N�3p}ll,��v�n"fgg�V�%�  p�V������_%/��׿����9YK   w,�U���"K�    �<ϯ=���ظ���Q���  ���������_~�a���k3"�#"ꩻ  �+ϟ?OZokk�F�EEQ�N3    ��t��k�loo'���g�   w�(�����^����po6��GD|UJW   w�ٳgQ�V�ջ��Y�    p?t:����z=VWWu�j�bbb"Y=  �D+��������?���?D��PZK   w�R�$�h411q�+����    �{EQ\;�}}}=j�Z��"����  H������_GDT��?�c�R��{D�i  ��M���ں���    P����7?���R�z   )E�o�ӟڕ����{e7  pW"˲d�vvvn�7��   �\��+�Jlll$�&�^����l�z   %x^���Z�����N   �R�^����d�fffn��I�    ���t����F��H�M���b�A   %�/+��  ��-..&�wӫ��   �<�n7���g{{;Q7���  (K��   RH=��6^n	�   @9�����,�bcc#Q7�j5�?��  @�� �'��l���T�z199y��!�    ��t:ח��b||<Q7�獕��  �4��  <KKKI�mmm��yw    H���]{6w78�baa!i=  �2	�  O���b�z7�G�   @j�Mo�����aU*w  �Ip  ����񘘘HVoyy�������n    �at�݁닋�155����gϞE�ZMV  �l�  ���r�{�e���s���繐;    $��y�z��{���us)�͔   ep  ���/�vwwo�7�<��N    ��t:���Y����v�n.-,,$�  P6w  �I����V������bLOO��o��    i\p_^^����D�D���E��HV  �>p  ����vvvn�|QB�    p��<�^�7p�m��8
�� ��H�  xr�ֻ��^y��B'    @?�Mo�T*�������K}�	  p�  O���l�k}�?sss7�&�   �ݺ.ྺ��V+Q7SSSI�  ��  ���eY�}wvvn�|QB�    pG���^�7p�m��8
�� ��J�  x�R����_y��B'    �箛�^�Vckk+M3�����  �}!�  <Iϟ?�F������l��Ϗ��/����    w㺀���z�����阘�HV  �>p  ��,˒Oq�����_Nm/�B�    nYQ��v����K��%�� ��L�  x���v�z_���P�/�    ��]7��V����F�n.�s�>�  �O� �'kvv6��ƒ՛�����K���   ��.ྵ��Z-Q7333I�-  �w  ��ʲ,��������C�B�    p;�<�n�;pϗ��݄��  �S'�  <i�_���D�e#=SEE��    ��]7���h���Z�n.��  p��  O���L���'�7>>���#?�˩�y��   �-�.ླ��j5Q7Ϟ=�f���  �}$�  <yKKKI����/�W}    F��y�z��{��,�&R�8	  p	�  O^�F[[[�h4Fz�(�_Mm7�    n���b����tҳ�,�bqq1Y=  ��J�  x�&''crr2Y�Z�;;;#?�˩��   ��t:��멧����G�^OZ  �>p  ��Sܿ���/�W}    �����=_���O�ͥ�����   �+w  ���gY������H�|>�]�    ��u��WVVbjj*Q7�J%��  ���  "��j%}a�e�Lq   ���.��%70����|T�դ5  �+w  ��k��I�}�K����    \���Q��b{{;aG��&  �3w  ��K�ijj*���Gz�(�_���<r   �\7�}gg'��z�n.���  �w�   �l6�ٳgIk~��^���σ�M    �Eqm��K��nbqq1*�  ��	  �F��~S_2��@�	�    0�n�;�<mrr2����J�z   ���;  �/,--E�ZMV�^��������2�^�)�    0�������eY�n"Z�V���%�  ��  �B�Z�����5���cS�   `4y�G���goo/Q7�RO�  x�  >S�ē��#=�y�=�s!w    ���\o��1;;����,�bee%Y=  ��B�  �3sss�j���˲,���G~�������w    ����_r��M���&=�  x(�  >�eY���5�����v�   �j�^�7#~�V����N��v  �>�  ����Y�%�7333���(~j/��w    ����������h4����T*�����  �C"�  p���񘙙IZ���h�g>�:e�;    �V���~||���KKKKQ�ד�  x(�  �X^^NZogg'Z��H�|>�=�s!w    ��N�3���ٳg�������6G  ��D�  �����V���U*�������B�    ������멧�7�͘��KZ  �!p  �Z����BҚ'''#?�y��w    ���yt�ݾ�Z-���vt9�=˲�5  w  �����֛���z�   @D�������f3Q7�R�9  <4�   ������XҚ_r%r����gS�    ���b����Q�N.������DҚ   ��;  �5��v�z����j�Fz���y��   �u�݁7>{�,���v#��  �	�  \#�K�J����#=S�o�^�   �cw���/�I�&*�J�@=  �C$�  p�������MZ���d�gz�ޯ>�   �TE�n��z�V�����E,..F�^OZ  �!p  ���j�z���#O��*�.�   �S��t~s��/���D��L�Q���Z�z   ��;  ���v�j��5������    <E׿���&��Ǔ�	  �P	�  �R����rҚ����j�Fz�����sQB�    <)�^�7�d�4;;KKK	;��ޞeYҚ   ��;  ����ד֫T*qpp0�3EQ����AW1   �cs~~>p���$Q'���  �	�  ibb"�5�GGG#?��t�<υ�   x���n��w�V��<T���h$�	  �	�  �`uu5i�����'��y>�w    ��\\\�����<l�����  �C'�  0�v��Z-i�/^����vw    �������_}�U�N.���'�  �p  A�R����5���G~	���~�;    �Y��x���Ϟ=K�����,˒�  x��  F���������H�����U��    <f�Mo���o��a   ���;  ��&&&�_+|xx�Fc�g>��^��;    �RQ��t��ONN���f"G>�  @�  �����&�W�����`�g�
�>�    �a��gY���K��  w  �/�n��V�%���W_����)�y��   ��
��j�8<<L�MD�Պ����5  w  �/P�Tbyy9i͙��X[[陫��_�    <T�Ng�����A4�̈́E���%�  �X�  |�����5��꫑�E���    <&���GD���$��R�R�����5  w  �/411���Iknll�\����    <4�^/��n�����x��Y"��h$�	  ��  �@S�G�8u���ϧ�   �Ct���QoD�e�  <&�   7���cccIk�<���EQ\|   ���(��t:}�'''css3aGSSS�o}  xl�  n ˲X]]MZ�^�����H�|p��z�;    <o*|��EdY���������   #w  �Z[[�J%�ϫ/y9�y��w    �����k�Z-v�h4��n'�	  �	�  �P�ш����5gffF�o�;    �E��x�����f3aG��   x���  �e\=�����E�+���    ����kY��˗/vsYsԁ   \M�  �LOO���lҚ���1???�3��   ���z��v�}�777���---���XҚ   ���;  �-Y__O^�իW#����7ۯ�    �����|xʸ�  �p  �%eLi��ى��ɑ��jb�)�    <EQ����XZZJ����333Ik  <f�   �$˲X]]MZ�R��˗/Gz�����;S�   x�����z��m0�  �v	�  ܢ����T���:>>yr�)�    <D���������f�n"�F��   ���;  �-*�V�V���㑞�7�    �����~�:�,K�Q9/   ;��   nYW�x�"��������2�~U�    �A��[�V���'�&"˲X[[KZ  �)p  �e���1;;��旼��*�n�;    �Q��8�a��aii)��fҚ   O��;  �X__O^s�+��<��JgS�   �o������j�8>>N�ͥ2�   �w  �;���cccIk�������H�\f�*�    e��z��v��%?�+�G  ��B�  �dYV��W�^����)�EQ��   ��1hz{�e��ŋ��\���N^  �p  �#kkkQ�ד�l�۱��4�3y���;S�   ��<�N��w}ww7���v�j�baa!iM  ��D�  ���j�XYYI^����#�jZ{QW�    �A��#F���6lnnF�e��  <�   whss3*��?�677cvvv�g�
��   P��(No_]]�����E���R�Z   <%�   w��lF��NZ3˲x���HϘ�   �}s~~EQ�]���vsicc#��j�   O��;  ����J^soo/���Fz�0��;    e(�"...��/--%��^�Vcmm-iM  ��H�  ��MLL$�*�R���   ����tNo��]�n.���D��H^  �p  H��)�1999��~avw    R;??�6??�|�z�e�����&  �S%�  ����\���$�Y�T�իW#=c�;    e���x��7�$�����B���'�  �	�  $RƄ����^�Eq����    �rqq�w���祜�mnn&�	  �T	�  $����|�S�Z5�   ����\y>�o߾M�ͥ������M^  �p  H$˲R�K���D��z�禸   P����k����������+�&  �S&�  ����J����5k�Z�|�r�gLq    �n�{���,�v111���Ik  <u�   	U��X__O^���$�����Mq    �����k��ӱ�����K��  �'�  ����zT*i�5�x���HϘ�   @*�LoO}��l6��n'�	  ��;  @r�F#VWW��}��e4�����   @*���}�&''coo/a7�������  p  (E/��F�����L�)i   �(z�^t�ݾ�eLo����   @�  �ccc������W��^���w    ����Yߵ���888H�ͥ��ͨV���   �  P����䓧���ne����   `X�Mo��M�3�Z�kkkIk  ���;  @I��Ƣ�n'�����h4C�7�   ��r�����Ä�\����D   n��;  @�vvv"˲�5����ŋ#=c�;    �����޽�j�����j�Ik  �k�   %j�Z������W���l��ߴvS�   �R���������~�n.mllD�VK^  �O�  J�����f�шׯ_��)�    ܖ릷��7Q���4��  p?�  �lbb��)�/^��V�5��~A�<ϣ(��j   �'`���gϞ�2b}}=�F�   ���;  �=���Y�%�Y���͛7#=3(�    �fz{곲J�bz;  �=!�  pLMM���|�'''1999�~S�   ��A�����ckk+]3����f3y]   ~K�  �����I>��Z���_=�3��   �������߿O�ͥJ������  p5w  �{bzz:�?�����aLOO�P�]�   �AMoo�۱�����K+++166��.   Wp  �Gvvv�׬T*��ݻ��1�   �Qu�ݾ�J�~�m�n.eY[[[��  П�;  �=233sss�����ųgφ�����(��|_��;    W4�}mm-���vsiyy9Z�V�   �'�  p����&��eY�}�v�gLq   `X�Ng���o��&a7��,�����u  L�  �������ϟ'����C�����A/+   xzMo��ڊ��ń�\Z]]�����u  L�  ���ۋ,˒�}���H�Mq   �:}ϋ�,�L�6T*����J^  ��	�  �C���1??�����F����������w    �����k�����f����V+y]   �'�  pO���R�w���H�Mq�~   �i4��Z��7�|��#��  �;w  �{jrr2�����]XX���ݡ�
��{y	   ��WE����]��eLNN&�����F4���u  ��;  �=���Y�%������V�C��v�W~o�;   ��u~~��l��l��ׯwt95~ss3y]   �'�  p�������r�SSSqrr2���(�Nk��z��    DQqqq�w�ݻw�LQ��ڊF���.   �p  ��vvv�RI����۷#�d�d~   �q:;;�;�}zz:���wQ��b}}=y]   F#�  pϵZ�XYYI^��lƛ7o��?(�.�   �t�y>pz����Z�&�����v����u  ��;  ����S�K��/_������Mq�   ��rvv�wmqq1vvvvs��h��  �@�  < �f3��֒׭T*��ݻ��_7Žߵ�    <�^/:�N��>$�擲H   0:w  �b{{;j�Z����1???��n��w�_�   ��a������h��	��466�����  �e�  �z�^�5ʣN���zW~o�;   ����v�?�T*���&�����NT*�   �_p   ���V����uWVVbccc���^�o��_�   ��m�����㘝�M�ͥ���XYYI^  �/'�  ���j����*���F�t�/�^E�y~[m   p\\\�=��������]��ݍ,�J�  ��p  x`666bll,y����888z��}���   <EQ����͛h�Z	;�455�v;y]   nF�  ���T*���[J�o��&���������E�w�    ���y�A�����]eX   ���;  ��������뎏�Ǜ7o��_E�i�&�   �0�y���}�?|��Z-aG��ٳg��  ps�   TYS�_�~333C�4��w   ���������R)gXY����^�   �w  �j~~>�?��n�R����wC�/��o�}Єw    �^��N�ʵ,����O�ѥ��՘��,�6   7'�  �����Rwkk+��ֆ�?hR��;   ��tzz�w���(vs�Z����N�   �w  �ljj*VVVJ�����G�2���AS��   �:�N�3�F��޽K�ѥ���h6���  �v�  <p{{{Q�V�ם���������z�(��ʵ<�4��    IDAT��   p�Eggg}׿��O�ѥF������  p��  �f�����~��]����ФvS�   �������ʵQ�"ܦ��ݨ�j��  ���  <����h4��m6�����Ф��(��   �~��<�������wQ���"������j�   �>w  �G�V����v)����baaa���n�;   ��vvv�wmss���"˲Rj  p��  ����O^7˲����?hR{Q���n�5    nQ�ۍN�s�Z�R�>$������H   ���  �,�boo����v;vww�����(n�-    nѠ��^�������\ʲ,�����  ���  <"KKK1;;[J�>D�Vz��I�   �/}�lZ�V�y�&qG����J	�  pw�  ����Ȳ,y݉���^d�z���ڋ��<�o�5    n�(����?|��F#aG�*�Ji7  pw�  ����XZZ*���W�bjjj���n��ڠ <    霝��=�Y\\�����]��܌V�UJm   ;  �#tpp�j5y�Z�?~z�u��Mq   (W�׋���+ײ,�,�65�����.�6   wK�  �*����zlmm�����]��\�   �D���}�^�x���	����   �=w  �Gjss3���K�����G�^joQ׆�   H�������x�{�.qG�fffbii���   �=w  �G�R����~)�'''��۷C���zQŕk��   �}EQ���Y����>�F>9<<�,�J�  ��p  x������~���H�����/    ��;;;�{���;;;�;����333��   w  �G���V�J%~�ᇡ��yy��]7�    �^�W�U�Ց�|nS�V����Rj  ���;  �#711kkk��n��qxx8��A!��(��   8==����_�6A}ww7��f)�  HG�  �	��ۋz�^J�>����P{���y��jl    n��������L�~�:qG����K�   @Z�   O@�V����Rj7��x�����{����)�    w�(�8;;����ǨV�	;����0*  ����?  �'buu5���J�}tt+++C�b/�"�<���    ����Ӿ����buu5qG�b~~���   �'�  �DdYGGG�eY)��ᇡ�l�y>0�~ݔw    F��v���\��h4�Ç�;�T�T��ࠔ�   �C�  �	�������Rj����˗/����v���   p;�����Ӿ��߿����}���QZm   �!�  ��E�Z-���w�bjjj���B��My   `8���}�Y���8qG��Floo�R  ���  <1�f3���J�]����z��QE��^�7p   ��z�^���_��eY��㏑eY�.D�V+�6   �p  x����bbb���;;;C�4�="Lq   ����Ӿk�^�������|277�v���   �K�  �	�T*q||\����?����P{���^��w=�s!w   �/pqq���eff&޽{���Ke�]  P.w  �'jnn.���J�=66>|z�׋�(�x   �_��<�������1j�Z>���,��A   �'�  ��F�^/����Alnn����0�   `ggg}������j�.������v)�  ��  ��F�����������y>0�~�:    �:�Nt:�+���������;����(��ji�  (��;  ����333�Ԟ���i�������N    �(�8==�����h4	;�dqq1J�  ��!�  @E�e��>99�v�=���B   �wzz�w@���^lmm�m���j�R  ��E�  ��������RjgY?��S�j����y>0�~�:   �S��v���\�666�}�]�>��ۋ�����  p�  ����l6K�=33o߾z�׻v��$2   ���(�8==�����G��J��'������^Jm   �w   "��胃���z�*����[ŵ!wS�   >9;;�{^���{{{�;����8�,+�>   ���;   �Y��:d~�*�J�����Je����Mi��\�    .�Q...�\k4�����}��������  ��p  �W��߶gϞ��ׯ����v�_�   x
~���k����brr2a7����R'�  p?	�  �+��㱵�UZ��o�����P{���^�7p�u�    ����Y�[����8qG�D�^/�>   ���;   �������ԮV��O��O�e�P����>L   �1��zq~~~�Z�V��~�)qG�������ri�  ���  ��J�'''C��o���R�z�j���nw�z��C�    ���?��w�Ç1==���O*�J�v�  ��&�  �����buu����|�M<{�l���Li7�   xJ���"��+�VWW���$qG�������Di�  ���  ���� ��f)���j���Je����^o���aB�    �A�׋���+��F���O�;�djj*677K�  ��'�  @_�j��i^ϟ?��o�����\����2   �������?���d�n>ɲ,NNN"˲R�  �0�  0���|�����y�&��;̔��&�   <dggg}��kk+���w�����ӥ�  �ap  �ZGGG�h4J�]�T��c�����`7�   x�z�^���_�666?��c�>������  �p�  p�z�����՟���o��v���nw�z���Nz   xH���������?��V+aG���W_E�"�   ���z  `(�v;K���ŋX[[joQ���<�v�;   �Cqvv��ֺ������N��'���1;;[Z}   w   �vtt�Z���?��S4�͡��z�k즸   �A�Ӊ���+�&&&�Ç�;�dll,���J�  ��#�  �К�f�Vbb"���w�݁��Lz   �ϊ����Ӿ��'''�L   ��p  `$+++������}�vQ׆��<�{}7   �}wzz���/^���Z�>)�	  ��I�  ��dY���Q�VK����V�5��a�^��`   �����":�Εk��������}�h4J�	  ��K�  ���Z����-����X���C�n�{�e�   ���<��ή\�T*����>j�Z�>9>>�z�^Z}   .w   ����f��ΖVkkk�)`ׅ܋�r   ���Ӿ7�}��ױ�����OJ�  ��&�  �;>>�J����?~:d��y�y~�=    e;??�����v;޾}���O��z�V  ��O�  �/699����կ�j��?�q�}���;���<�v   @Yz�^���]��h4��CdY���O�����l�V  ��O�  ���ڊ��������Ƿ�~;��~����(
S�  �{�(��������1���v�k�v;��vi�  x�  �����*j�Zi�_�zkkkC�-�"z���=y�_�    �������tt{{{�;���l���Qi�  x<�  ��V������ϲ,���?D��j�׋�(�����=    �t:�����rmzz:����}�eY���D�^/�   w   n���Z��ϗV��j������w��k���   �y�����k�J%���?�._]]-�\  ��E�  �[S�������ꫯ��[ŵ!��(��  �ҝ����i����������Oʾ�  ��G�  �[�l6����g�Ξ�ʷ�`����)40H F!@B�T�P�Uԩ����u���v����8G��o}c;�5����(7���;�s�[��^jg�{�ۥf��obrr���<�#��3J�   @Y���}Hff&�޽��D�s�N�j�R3   �eQp  ���������Ү_�V�ٳg]��������   �eY{{{mφ���ɓ'��W�^����f   �ˣ�  �'w���,�������7�t=��-��Ex   �O�(����9������h4z��]###1;;[��  �r)�  ������s�N$IRZ�����z�jW�EQD�e=   �����F�����r�J��?I����bT**   |z�6  �,&''czz���?�S�Nu5�e١?���   ����A�Z��g�����D�����R3   ��Rp  ೹}�v�v����x��Iכ�)��yޱ   p\Y����n۳Z�/^��Z���T����h�o�  ��Pp  ೩V����Xj�.���ZW�EQD���,��(>6   �;������C�>|ccc=L��j�KKK]/   ��Pp  ��+W���aee%.]���l��]mr�f   �(vww}s���|ܼy�ǉ�577�F��   |��  �����btt���'IϞ=�S�Nu5�͆��(��  �O��� Z�V۳������o{��]gΜ����R3   �uPp  �K�$����V���app0^�x�Jw��i�v��v�;   ��dY{{{m���z�x���U�Ν;�$Ii   �z(�  ��F#nݺUj�s�����fW�EQt]r��   �0EQ���Ρ�/<y�$���z��]���100Pj   �
�   �̅bjj��w�ލk׮u5��y�y�q.�2%w   �Xvww��aii���1>��W����d�   ��(�  �S�oߎ���R3<~�8FGG��MӴcy�(�Ȳ�SD   �"�j�ڞ�;w.�߿��D�����R3   ��Qp  ����z,--E�$�e���>j�ZW�i�v�Qr   �"˲���m{688ϟ?�J������j,--��  ���;Q   znll���kONN�7�|��lQ]���<Wr   :*�"vvv=��q4��&z��۷��h��  ����;   ��������R3,,,���\W�ݖ��<�<�?6   ����=�������z�jo�����ǅJ�   ��K�  ��,..F�^/5�Ç�.�gYEQ|�9   �볿��V�����t����8ѻcaa��   |��  (���P��ϗ��^�ǋ/�V�u5����m�   ��%M����k{6<<ϟ?�J����$��w�v�=	   |
�   �����q���R3����Ç����^��;   �<�cgg��Y�$����h4=N�����+5   (�  P�[�n���H�n޼w���j���z��J�   @DD���DQm��߿.\�q�w����իWK�    
�   �j�������;"��o�����f�,�<�;��y��   �����=�!�k׮�ݻw{��]�z=�ܹI���   "�  ����177Wj�J�/^��z�|���n^�ײ,�j   ��Z�888h{611O�>�q�w%I1<<\j   xK�  ��q�ҥ8�|�����իWQ�պ�OӴ��ö�   _�,�bww�����`�|���� >�K�.Źs�J�    ���;   }��ưF�Qj�3g�ģG���-����{QJ�   �)�"vvvھ�-I�x��Y�������9}�t�o�  ����  @_��jq��ݨTʽe��������f�<�<ϻ�Sr  �����Ρ�lnnƥK�z��]�z�/��  ���N  ���l6�֭[eǈ���tW�i�����ה�  �˷��w�߮]�����q��---���P�1   �=
�   ��������K�R�/^���HW�V��{7�  ����j���~۳���x��i���ڵk199Yv   hK�  ��5??�u��s���>��jW�mg�kY�uU�   N�,�bww�����`�|�2j�Z�S�k||<fggK�    ��  @ߪV����\���Ν�G�u5[��;   |����������I��ӧOctt��d����@,--E�$��   �Qp  ��5����/;Fܼy3����<�,�8WEWs   @���ى<�۞mll��˗{��}���188Xv   � w   ����T��̔#<x���]�fYv�����;   �|��������ի�����D�q�FLNN�   :Rp  �D�u�V��T*�����j>MӶ�%�k�n|   ����A�=�����O��8��Μ9׮]+;   tE�  ��R����R�j�Rs4�x��U�9�����<�j�;   �?�4���ݶgCCC���˨��=N�����X\\,5   ��;   'F�ш���H���gΜ��O�v��(��K�Y�)�  �	��y���=�T*���ߗ�6�$I��ݻ���  �(�  8QΞ=�.]*;F\�v-��׻���<�,�j6˲(��c�   �YQ���s�=��Ǐczz�ǩ�777ccce�   �#Qp  �Ĺy�f����#VVVbnn��٣lgWr  �����s���G���s:w�\\�|��   pd
�   �8o_�=44Tv�#mdKӴ��zQ]o|   zkoo/�4m{v�7�}N�f3#I���   ��)�  p"Ľ{��R)�ֶR�������]���_Sr  ��spp���m�Μ9O�>-�T^���޽{Q�VK�   ǥ�  ��5::eǈ���x��Ut�-�"Z�VW��繒;   �4Mcww��Y�шW�^E�V�q��---���p�1   ���  8Ѧ��cff��1>>/^��j�|Q]orWr  ���y;;;m�j�Z�|�2FFFz��}sssq�̙�c   �GQp  �Ļ}�v����#fff����]�����   �)�"����(���?�s���8��Ν;W�\);   |4w   N�$I��ݻ144Tv�XZZ�����f�,�<ϻ����Y   �����9��|ss3fgg{��}###���I��   >��;   _����XZZ�J��[��ŋ��MӴ��z�e�n�   >����HӴ��͛7cyy�ǉ�W��byy9��j�Q   ��(�W   �D��ƺޞ�9U*�x��E�>}���4M�.�e   8����888h{655�=�q�������h�   >w   �(���133Sv��~�!�����?l\;6�  ���j�boo�����h�|��/6����ř3gʎ   ���;   _�۷o���x�1������?F�V�8[E�Z��>�(�Ȳ�c�   m�i;;;mφ����������ܹsq�ʕ�c   �'��  �'I��{�n�%Ξ=/^��$I:�E��&w%w   ���<?��^���իWq����z���H,..v�}   �4
�   |���ݻQ���{���x��aW�y�w]\?�,   �aEQ���vE��Y�$��ٳ8�|	��U��byy9��j�Q   �(�W~   �L�������eǈ������w�^W�Y�E��]�*�  ��{[n?�~��o���W��6TI����R4���   �g��  ���ŋq���cDD������͛]ͦi��   =���{����r,..�8Q{7oތ3gΔ   >+w   �x�n݊�gϖ#""�����j6MӶ�EoG�   �gww7Z�V۳�������q��.\��7�  ���  �Waqq1��f�1�R�ċ/brr��y%w   �|�������م�ɓ'�t���񘟟/;   �;   _�Z���݋��������@���q�ԩ��EQD��]v������  ��B�Պ����g������˨V�=N��F����Q��y  ���;`   ����q�޽��A��hď?��U�(�C_��N�eJ�   �i����N۳�ܳn�z=VVV�V��   z��_�  ������Ν;�$I�Q��ܳ,��(>&   |��,;��~���}nI��ݻw��h�   zJ�  �����T\�z��q�x��IW��<ϏTrO�T�   ��<�c{{����ѭ    IDAT�r�R�/^���d	��w��혘�(;   ���;   _���٘��*;FD�K�����f�<�,˺�l��  �_|����ɓ����q���\��7Y   ���  �*%Iw�܉��Ѳ�DD���rܽ{���,�"��f��Pr  �WE���z?��7�č7z���3g����\�1   �4
�   |�*�J,//���`�Q"�_~L�}�vW�i�*�  @ޖ�{#���j��n###���I��   J��  �Wmpp0VVV�Z��%""=zׯ_�j6MӮK�J�   |�vww#MӶg�����D����XYY�Z�Vv   (��;   _�f����eǈ��$I�ٳg133��|��Rr  �C���F��j{v�ƍ�����'j�R����J�   J��   q�ܹ�q�F�1"�_~�~��e�?��y��  �}{{{qpp��lff&�<yI��8���$�;w���ӧˎ   }A�   �׮]�K�.�#""j�Z�z�*���;�Eq���ϲ�c�  @_��ߏ����g�ϟ��/_F��?�߸q#���ʎ   }�?��  �Oܺu+Ν;Wv����ׯ_G���8[š�\?l�(�x   8)boo�����D���Q��z����/�իWˎ   }E�   ��$Ibii�o^>22?��S4���J�   |�bww�����h�~�:{����g����|�1   ��(�  �_�T*����U������;   _�V�uh��(����ӧcii)�$);
   �w   h�^����j�%"��
���֋��,�>&   �*M����i{644�_��f���T����rT�ղ�   @_Rp  �C����ϟ��/_F���v>��#���<Wr  �DJ�4���۞�j�x��U����8U{��@=   �#w   ��~{e���L<y�<G-��   e˲����J%^�|�ϟ�q��*�J���D��(;
   �5w   ���ٳ1??_v��ݸq#>|��l�eG*�E��  ���eYlooGQ�U*�����cff��d�K�$�������eG  ����   ]�x�b\�z�����������Y%w   �4*�'IO�>�+W�����[�nŹs�ʎ   '��;   t�ƍ1==]v��ݾ};���ۮf�,�<ϻ�l%w   �U�����%$k�ڵkq�ҥ�c   ����   ]J�$�ܹeG����R|��7]ͦi��  ��֩���ɓ�q�F	�ڛ��ꫲ=   �
�   pI����r4�Ͳ����ݻ����լ�;   '��r�a��>�����:���xܹs'�$);
   �(
�   pD�j5���cpp��(�[[[�����f��  8i���Xn����q��5��X^^�J�O�   pT�  ����b}}=ʎ򻍍�X^^�jV�  ���S����������T�������jeG  �I�   ���h���j������nss3�ݻ���qK�EQ7   ��r{�emϏr��������Wo}  ��F�   >B�ٌ{����+Ǐ���8%�,˔�  ��:����׻~�Y/���XYY���Უ   ���?��  �	5>>w�ލ$Iʎ����|W�J�   ��N�����X]]�q��U��X^^�f�Yv   8��  �8{�lܹs���x��Qܾ}��Y%w   �E�r���R����8��*�Jܻw/���ʎ   _w   �D����.��ʣG��ƍ]ͦiz�º�;   �Z�r���b|��=Nu�$Ibqq1&''ˎ   _w   ��.]�ׯ_/;��$��O����\W�V��%���  ��N�����x��A�S.I�������ϗ   �(
�   �����ƕ+Wʎ�$I�ɓ'q��ͮ�Zr�����y�'   t,�߻w/>|��T677/^,;   |q�  �3����.��woK�]���e��;   Gܾ֩������q��v�Z_=�   _w   ��$����8w�\�Q�����X\\�j��j����  �Qt*�������f�S}؅bvv��   ��Rp  ��$I�XZZ���񲣼��������l���*�VL   ��:��766bmm�ǩ>�ܹs���I��   �X
�   �U*�XYY���Ѳ����o����ծf�Sr��\�  �Cu*�������T699KKK��   �)�  �gV�Vcee%FFFʎ�����7�)�  �t*���c�2>>��݋J�O�   ��  ������+�������fW�J�   |�<�ckk��{Ň���b�S}���X,//G�Z-;
   |�  �Gbuu5���ˎ�����~W�J�   W�籽����2I�x��I,,,���p�f3����V��   �
�   �CCCC����w%�{���Ç��=n�=M��D  ��M���͛%$;\�ٌ������eG  ����;   ����`����]�}aa!=zI�t�M���[ً��4M�(��F  �ʲ,���ږ�+�J�x�"���JHv����X]]Un  �(�  @	���cuu5ˎ�����K�Y���e��;  �W"˲���n{X�V��ￏk׮���p�F#���b``��(   �URp  ��4�X__ﻒ��۷�ٳgQ�t���%�4M�n�  �ˑ����Z��^��+W����p�z�   _w   (Q����W����Ə?��U�������;  ��)M����i[n��~�)fffJHv����X[[Sn  ��)�  @�N�:kkk}Wr�x�b���O144�q6˲H����8n9  ���j����h4�����ϗ��p��������=0   �y)�  @h6�����Z��(�8w�\�����h4:��y~��{��J�   _�������i{6::���KLLL�8Շ���Z�   w   ��f3VVV���>>>o޼���ю�J�   _�������m{611���KW���400���122Rv   ����   }dll,VVV�Z����f��-{y�G��:�5��  N�������k{655���KWo륷�ە�  ��(�  @�����+�7��������g��8v�=M�(��8  (���n���=�|�r�~�:z�����z���ƩS�ʎ   �w   �C����Z��(���~�)fff:ξ-���^EdY��  p������A۳7n�˗/�������f�Yv   �w   �S��㱲��w��k�Z���q�����SrO�4�<?nL   >��(b{{�зw-,,�ӧO�R鯟���  ���׷	   �;���b}}=��z�Q�Q�T����q����Sr��Ȳ,�,;��  ���-��i��|yy9>|I��8ه���z�:u��(   �(�  @������+�'I�}�]ܻw���V�u���y�+�  �<�ckk����o��&677{��������؈�����    (�  �	�l6cmm-ʎ�����7�|��l��J�   'T�e�������R�ĳg���ݻ%$�����X__�F�Qv   �
�   pB4��X__���������ݻ����G�Z�8�����y�G��Q�q"  ��4�����d�z=~�ᇸq�F	�>��h���z�   蒂;   � ###}[r�v�Z��������Y�E��G�FQ�e��;  @Zno4��/����L	�>�m����T   �(�  �	�h4bss�/�ϝ?>~���8u�T�ٷُ�(�H�4�<?ND   �`?vww۞���ǯ�����=N�Y??    |��;   �@CCC���֗%���3g�t���<Z�ֱ��eYdYv��  ��������k{v�x��MW8�Z�ٌ���v   8��  ������h4eGyO�ш��9.]��q�(�h�Zm_u�I��J�   �XQ���mϯ_�?��c�8Yg�������z��(   �1)�  �	644122Rv�����x��Uܾ}���ǖ��4=��  ���4M۞/..���ϣZ��8Yg��������   '��;   �p���ޗ%�J��}�]���u5�j�"��#_�(�ȲL�  �#�y[[[mߔ�$I����M<x� �$)!݇�����   _w   ����F���������x��qT*���HӴm����("M�c�  �vY����V�{�j�ϟ?�;w�����XYY�Z�Vv   �Pp  �/D�^���՘��(;J[�n݊~���mzY�����  �5j�Z������X�����O?����KH����T���F�Z-;
   ��(�  ��Z����J�?��(m��������8�eY�iz���y��  Ѕ������i{6::o޼���������L,--E�$eG   >!w   ��T*�XZZ�.����g�ƛ7ob||��l���j��u�<�#MӶ  ���ى����gSSS�믿���X�Su��ի1??_v   �3Pp  �/P�$���W�\);J[����믿��˗;�E�V�XE��("M����81  �HEQ����������ׯchh���:K�$n޼ssseG   >w   �B�����z=^�z���gߖ܏[Tϲ,�,;��  |I�<����HӴ����Z<�<j�Z��u�$I�������   ����J    ��իW�V�������(�I�$677��l��O��c�=MӨV�Q�V�|���}��  ��i;;;mߐU�V����q�ƍ�uV�Tbii)Ν;Wv   �3Sp  �����L�j��o��-2�m~~>FGG�o��o������Y�EQ��&��yE�j5�$9n\  ���� vww۞5�x��U�={�ǩ�S�V�޽{199Yv   �*e    zcjj*����R�ϯ.^����[���u���<�4=�u���4M;n�  �R���Zn����_��o��Z-��֔�  �+ҟ�h   �ř3gbuu�X��{������͛�p�B��<ϣ�j{#}�e�eٱ�  �$(�"vvvb����k��͛7q�ԩ'����`�����ӧˎ   ���;   |e���ccc#ˎ����`�~�::�E�Q%�������   �*����ڊV���|qq1^�xѷ@���F4�Ͳ�    =��   _�S�N���z���J�>�D�$�[�V�y~�kEY�)�  _�4Mckk��}R�Z�'O�t}�U�f����1<<\v   �
�   �j4q���-;ʡ�~������i�F�eǺNQ��   ���� ����>�;44�_���7o���;�����}    �eRp  �����@���Ǚ3gʎr�K�.��?��N��8�eY�iz�k�y��  �X{{{�����lbb"~�����q��MOO���j�j���    %Rp  ��\�Z����x�b�Q599���ʘ�y�Z���
���y�iz�  赢(b{{;���۞_�r%~��h6�=Nֽ˗/ǝ;w"I���    %Sp   "I�XXX������jhh(~���X^^�8[E�Z����X�*�"�4=��  �J�e���u�۬����իW100��d�I�$����֭[��   @DDx�   �W����@��/���J%677cbb"�������[i�F�Z�j�z��eYEQ��  >�V����m����ӧq�ʕ�u�Z����R�={��(   @Qp   �q����_�kdYVv��nܸ������ݿ������ےz�v��A�<���n�   �/���b�����D�|�2FGG{��{�z=���cll��(   @���    �?������eG9���d���oq��Ŏ�y�G��:�V��("M����X  �E��ۇ�ۯ_����k_�ۇ��cssS�   hK�   h��l���F�����PCCC����X^^�8[E�Z��*�gYַ[� �/_�e���i��w�$IlnnƋ/���^8}�tlnnF��(;
   Ч�  �C���F�����PoKϞ=�đ��G���<�4M��  �8Z�Vloo�}hwpp0~��Ǯ�-�ٳgcmm-ʎ   �1w   ����z�������ˎ�A7n܈7o�D���8�eYۍ��*�"�4��m�   ���ۋ�����NLL�o��333%$��ŋ�޽{Q�Vˎ   �9w   ��J�KKKq�ʕ��|���d���oq��Ŏ�y�G����M�Y�}�6x  ���<���b�����l���1::��d�K�$�_��$I�q   �@�   �J�$q��͸y�f_�������ױ���q�(�h�Z��=��H�����   -M����j�Pm�$���ϟ?�Z�VB��T*�X\\���ٲ�    'H�~�   ��+W����H����4Mˎ��۲���d����}�Z�Χi�j5��걮WE�i�J�؟  ����A���=��ϟǅz��hcyy����   ��w   ��Μ9144Tv�����?��111�q6˲�E�N�<�,�ls  ��(����9��>==�ӟ����l6cccC�   8w   �XN�:�|�M�����N�>���[���w�-�">��������?  ��dY[[[�>x���?��S4�';��D�   8��  �c��뱺����eG��j��=�'O�D�V�8�j�"˲c_�(�Ȳ�>  �z�Z����n�����P��������T����˗/���JT�ղ�    'X�_t   >�R����b���������8t���8w�\����m����>8�eYE�U!�0y�GQQ�V#I�c  �e*�"��������ٳg�ŋ�l6{��h*�J���ǅʎ   |��   �ĸ|�rܽ{��7����ů�����g�<�V�EQ�zEQD����  ���<���-����Ǜ7o������^��   ��b�;   �ɜ?>�F����_b��8��������t�R��?�C�iz�lQ�j��Z�~Ty?����͆�� �׭�j���nۇi��z|��w]=�[�F�+++�h4ʎ   |Alp   >�f���ߏ��Ѳ�tt�����_�ʚe������<�,���  |}vwwcgg�m�}rr2���?��r���Dlnn*�   ���;   �����FLMM���3g����Ǹ~�z��<ϣ�j�-�t�(�Ȳ,�,;�g   'O�籵�m�����͛7'�a�/���j�����    _ w   ೨T*���ׯ_�$Iʎ�A��ŋx��AT*���(�h�Z��=��H�����  ���j�bkk�탮�Z-���x��i�j��u/I�����������   N����   8ђ$����h4���K����b�={6����.�������i�F�R��JQ�N�Z=��   ��(���ݍV���|rr2�?ccc=Nvt�z=�޽eG   �p6�   ����tlnn���p�Q::�|��O������y���  ��eYlmmZn����7oޜ�r{�ٌ���+�   =��   ���B���d�Q:��O�Ɠ'O�^�p���,�>ꚟ�s  �����Vۇa����~�G�}��z���󱱱q"X   ����	   �Ũ�뱲�����������tt��͘�������������g�,�<ϣV�E�$Ǿf��QET�Տ�  ��������HӴ��ŋ��ӧ�h4z���$�7nĕ+Wܛ    =e�;   �SI����\,--E�Z-;NG�f3~���X[[�X�(�"Z�V�-�Ga�;  �<i����V�r{�R����x����(����X]]��W�*�   =g�;   P����������ݲ�|��2���t����b{{���i�F�R�Z��z��  N�������k{666Ϟ=�3g��8��4�͸w�^�   �J��   ���l����cbb��(]�p�B��O�+W�t���<Z�VE�Q�|���c��T���    IDAT  �^�籵�uh�}nn.~��Sn�������v   �T
�   @���z����իWOĖ򡡡x��U<y����(��jE�e}�,�"Mӏ.�  �F�Պ������ĳg���ӧQ��KHw4I����\,--E�Z-;   ����d   |o��f3��|�B��v���8{�l�����������,ˢ(����N�ns�T*J'  P��(bww7Z�V��s��ųg�btt��Ɏ�^����RLNN�    "�  �>255###�������[v�������_�����s��/��l��qpp�Z-*��{�^��QET����  �i����N�7+U*�XYY�����z�ٌ{�����p�Q    ~�q��   |b�f3�߿eG�J�V����ׯcdd��|�����G_��6����  N��(boo/���ۖ�GGG��C�����r���Tlll(�   }G�   �;�z=VWW����eG����L���oc~~��l���j�"��n�瑦�'�,  �}Y����V���=�����o�MLMM�8��T*��u�V,--E�Z-;   �{je    h'I�����������eG�h`` =z/^�������Cg�n`�T*Q�}�W4EQD�eQ��
  |B�����_�ԩx��q\�x�ǩ�ohh(���bll��(    �Rp   ����Dܿ?���?�������8]�~�zLOO����1���郳o���j�H�䣮��yE�J%*/� ����<vvv"��ػӧ��4o�߳�H�,$$!#	b1�'N�=�����t�t����;[�O��t�xc��+����H�m��Б��T���/��q@�n���
]�xQ�p�œ}�D"�cǎ)
=
     ���    @ۋD":w�nܸ������Ho�F�������7�|�j���Y��U�VeY�Go`g�;   �q*��J�Ҏ���Fu��E������������Ƃ     ���    ��`�&&&���믿�V�=�;)����iyyyϳ����ms�<O�i�   ���<mmm����lV���o������>\8։'�ł     ���Z�     ��$	}��g���z�w��ݭ�����x�l{�}�m��6�=�S�V눭�   @P*��^�x�c��8�.^�����������}��g��     ���     t�h4�s��i~~^���A��Φ���N������Z[[��l3�����Z��6w   �5o�ڞ�d�w�w���n�d�0�r9�����K      ��     t$�4599���~]�|y� ���b1���/���?����<o׳�m�e5%L�<O���4M�&/�  �íR��T*��jG�m�̙3:y�dGE�PH������A�     ���    @GRww�~��g�x�"�qމi�:uꔎ=�����֣G��<��m��6B�N�u   �fx�����a����Uooo�'�8���:~����pУ      |Vu    ����եO?�T�L&�Q�K<׿������o��^���nSn��<�j��}<   �T*�x�bǸ�q}������~�Qq�a�f�:{�,q;     8��     �4533���>]�~�c���6�B����������盹�]z�׷��&�   p0�mk{6��_|����O�qB���;�D"�(      MC�     �L&���~]�tIϞ=z�w��۫�����z�����[U��]�ַ�[��������}��+�����   �vR�TT*����ׅ�a�?^���L�q4;;��v     p��    ����K�ϟ׭[�t�֭��y/���:z�����WKKK{�ݏm���4MBw   t<�u�����;
}���D"-�������Q���=
     �� p     �aS,��˗U.���������t��-}���*�J���os7MS�ݜ�z<ϓ��2MS�i6�c   �T.�w���ե/��B�|��C5A$�����ł     `��    �mppP�}���\�������y/�BA�tZ�~������<�y��ժ,�jJ����\�m����   �7�u���)��v�~bbB�����p�'�x�tZ��Ӽ�     8��    ���8�N�<���e]�vm�إE�Q}��*
��믵����Y��U�՚����<��IH  �����J��*�ʎ������ŋ�d2-���Y����i���G     h	w     p(��L&���>]�tI/^�z�����N���w���ի{��<O�JE�m7e�{�cַ�7�c   �P�մ����Y���Ԕ.\�д'��Roo�N�8�h4�(      -�y��      |���n}�駚�����b���qt����6��O��y�V��0ٶ-�0>��}ߗ��<O�e5�c   ��<�J%U���O$�x���x�'k�l6�b���n     p��    �C�4MMNN���_W�\�5�iW�LF����+W����W�V������V��,K�e5��}�W�Vkls'�  @�U*�J%����u���ܹs:v�XG�W��:~������      �     ��R__�.]��Ǐ=�{1MS����f���ot���=�o߼n�fSf�<O���4ͦ��   �^\���֖\����l6��/�ȑ#-��9���433�P(�(      �!p     �Z8�ٳgu��ݼys����W�������}��7z��Ůg�o^���=,�y�|�olt   ���}�J%U*������_|��G��x��,K�b�c�     h&w     p�����Q%	���z��y�#��\.�L&��Q���<�����y�T*�,�i��}�eK�aM��   @�V���֎�qm��ɓ'u�ԩ�}U���>��Ϊ��+�Q      ��;     �����֧�~�[�n������ݶm�?^ccc��믵�����z�n�vӂ��[�M�$t  ��<O[[[��j;^?<<�/��B�X�œ5G����B���      ��     lc�������믿jss3��������?hnnN�~��J�Үg}�W�Z�i����=T�y�<ϓi��I   ��}_�Je���]]]:����b�'k���n��Ϊ��'�Q      ��;     ����t�������ݻ��]��Ţr�����{]�zuϳ��Z�ʲ,��ٴ�  �>j������y������)}��r'��>�a��rk��n     ����     `�ijrrR�x\W�\�sz�
�úx�������_�ɓ'���}_�ZM�aȶm�Ѵ9<ϓ��2M��   o�<O[[[��j;^?44�/��B�x�œ5O4���b�XУ      �5w     ��ԅ477�{��=�ֿ������������}�W�Z�i����=|���\ו�y�,��=   :����T*��?����ٳg555ձ�����&''yU#     �w@�     �l����Lc�{�Zz��f�����U(����E�/_������<O�JE�e55ĩo��os��P	   �Z��T*��7�3MS333:w��	`��D":v��     �c�     ����!�b1]�rEkkkA��A��>��s�E��O���ʞ��[�m�nj��y�<�#t  hS�W�i6�uU*�T��v�>���7���b�X�o���ɤfff���H      ���      �'�qt��)����ʕ+��9�.��_��_����o��F/^�������V�2M���;  @{��?k��2��U.�U.�w����O.\P6�m���8������PУ      t$w     ��L&��ק+W��ѣGA���r��2��~��g����{���R�Ȳ��o�$t  �����d��z�R��T*���7��?��ĉ2M�i��T*���I9��(      ��     �#D"�9sF����z����j�#}۶u��YMMM���������]ו�y�,����н�=   ��z��L�ZM�RI��q�a�g�}�h4���n�p8���)��     4�;     @$�I����ڵkZ]]z�v��}�嗚��ԟ��'����z��}�j�F�����   �k?�v��T*�v}��А>�����hlm�BA�     p �     4��8:q����t��U���G�`���������y}��*�J�����v�n�<O���4ͦo�  8��3l�}_�ry���G��'�|�b����n�h4���=
     ��B�     �d�DB�XL���Z^^���A��A�P�XT.���?��K�.�u�]�{��J�"˲��q��}��+����  ���3l��J��R����_۶5;;�ӧO�M�LF����7     ��      � 
iffF�tZW�\���f�#}�p8����kffF��_u�ڵ=�}�u���5B{�"  ���ﰽV�ikkkǏo��&''u��Yuuu���Rww��;���ޠG     8��     �Q�>��3ݺuK��]z�\�xQSSS��ﴼ������M�l�,�?GBw  ���w�J��j�ڎ�g2]�pA�r��d�r����ƚ~�      �"p     �g�eibbBCCC�|��666��$	����׽{�����������g}�W�V�a�m[�a4u�z�^�Bw  ���=�S�\V�R���D"��>�L�tz_n��b���������(      ��;     @�����ZXX�͛7�-8j�L&�?�񏚟��������]����j�*�4e��������  F�����r��r�������:w���~������1�r��?Q      �#p     h!�0���588��W���ӧA��Q�P�XT�PЯ����~�i�M���m��JE�e�[�N�  �V��JE�r��
:ۅ�a�<yRǏ?0��5==�h4�(      ��;     @ zzzt��yݿ_ׯ_W�Zz��b۶N�:���)��㏺r�ʞ���r]��  �#�w�.���t�ijffF�Ν��8�6C+��aMLL(�N=
     ��E�     �t:���A���ieeeǍ��$����?�������;-..�y�u]y�'�4[���)�0��v   Z�a��2n��6�����>��uww�����d499ɓ#     F�     0�q4;;�L&��W�jcc#�>Z����+=x�@?����ݻ��Y����eY2Ms_f���;  �T��}��Y���d2}�駊���:C+���hffF���A�      �     ����~]�pAw��Ս7v��:��А~���ieeE?����߿�����	�  ��]�����+�H���d۶���422�}B     �6B�     �F�P6�U"�еk����àGj�T*���ֽ{���w���y��cw  �v⺮|�4lO&���O4<<��3�Z"���Ԕ"�HУ      �5�      m(�����Z[[�իWU.���)2������M���������m���U����O�  ڂ��<o�o��FD�����9sF�Ba��h���.MNN*�=
      vA�     ����t��--,,����V��r�f��}�����{={�l׳��Z��4MY��o3� � ��/������u�������|>���Q��     �9w     �6gY�&&&�J�t��U=}�4葚�0
��y]�~]?���666v=_��G�����=�k���u[   ������ԩS���:p�}455�#G�=
      ��;     @�������絴��7n�Z�=RS�����iMNN������_�����]��j5=}�T�HD����N���.�;  h��O�k�m��www���Ӛ��<p����&''�L&�      ��     ��=zT�TJ�o����bK�}�B=tׯ���K�.�T*�z�T*�T*)+�,t���   ���C�^��~��ۘ��l6�B� ˲�      ��     �ٶ���	e2]�vM�=
z��	�B:}���?�k׮駟~�s�{�\V�\��8
���1�c�z$F0  ޅ�������ĉ���>��e��&''�F�      ��     ��uuu�̙3Z[[���׵���HMc۶fgg5==���9��������|�RQ�RiY�.I�Z����0�}�=  Й<�k��������^�<yR���nc�$9rD�bQ�x<�Q      ��     �D"���A---��͛��jA��4�eizzZ����q�~��G={�l��ݥ���뺄�  ����}��|�no�����_'O�������m���ؘFFF�     p@�     �i*��*�Lj~~^+++-��Z�4M�E����ƍ�駟��ɓ]��C�P(�H$���]Ҿ�  h/�M���.���ĉ���8��a�����	z      4�;     ��5;;��������w�z�>11�۷o����c�ZU�ZU(R8�m��Cb���V��� �C����]����A�>}Z�B�e������Ţzzz�      ���     ������'�|����knnN�J%葚�0
���jqqQ��_����]Ϸ:t�^��^�� @����s�
�S��N�<�\.ײyZ-kbbB�t:�Q      ���     �t:���!ݹsGw��i�v�V0C�\N�\Nw���_��W����z>��}{ �Vw  :S=lo��)�u���e2�>}Z���-���,�R.����(O     8�     ˲466�t:���y=x� ��E>�W>���ʊ~��'-..�z��[��p8�P(���y=pg�;  ����r[��{�n�FFFt���t�V2C�tZ���
��A�     �!p     8D���t��I=}�T���z��q�#�T*����JO�>��˗u���]�������M���H$Ғ�]zs��eY�~�  ����]�=l�m[:q����Z>W+jbbB===A�     �#p     8����t��9���innN���A��/���������Ӻr�~��W����z����Q8nY�.I�Z���  �������/�uw�Ѩffft��1E"����j��ݚ��P<z      ��     �K$���Z^^֍7T�T�i_D�Q�={V'N�������/��ŋ;��<O�RI�R���j���[�M�lId �aWڃ�־W���۫��YMMMɶ���"��
�������     p��G�      �V�a(��(�J�Ν;�s�N qW+�B!���jffF7n��/������]�W*U*�B!��ᖅe���u]�� �O�A��'����yr]w�ێ�㚝����ā��-�R.����(�w       ��      �ǲ,���)���֭[Z^^$�j�4U,U,�����~�I������V��V��m[���q���Z��<�k��=t `?���~�;��ahddDǏW&�	d�V2C���o�}+      �?w      �"�hffF�\Nsssz��a�#�T*����Jkkk��_t���]��Z��Z��r��p8�P(�������Vw��  ��Ճ� _��u�F\��mۚ��������������Ţ����      m��      ;:r�N�>�G�i~~^ϟ?z�}�H$���������ܜ._�����Ϻ����M���H$H�.���hlv  S��믆�u�����������;�H$�d���קb�xhB~      |w      �ippP���n޼�R��H����K�N�҉'t��]�tI���;��<O����$�q�[�U��y�G� �Ԉڃ��^Օ�fH�R���U>�?4߳���5>>�D"�(      � �      x+�04<<�t:���eݼyS�r9���i�*
*
z��^�����7�JR�RQ"��y    IDAT�R�m�r��[ݥ����-��i�|  ��Q{}�u��oY�
��N�<������k�H$�B����a�      ���     ����L&�t:�����ƍ�T*A�����.^���g�jnnN�/_���Ǝgk��j��L�llu"t�$�u�M� 8h�A{�Q��{���ե��i;vL�H$��Z/kll��      ��      ��4Me2�R)ݽ{W�o�V�Vz�}��եS�N�ĉ�s�.]������z��R��R���-�j��o��a�4͖� @3ԣ��X�,;��K*�����������8�r�������     �\�      �`�e)����ѣZZZҭ[�v���4U(T(���C]�tI7o��u�l�RQ�R�eY
��
�B�l3�ǀ��� :F;E��y\�}���eY*
:y��.�PH�|^###�<�      �;      >�m�����d2�s�w���x<�/��R�~�����t��5={�lǳ��jssS�i6���K�� ���nQ��ƶ����b*����R$	h�`X�������ʶ��#      ��G�      �4�PH�����M���եS�N��ɓZ^^�իWu�Ν?��T*�T*��8��	4
#v ��v���3��
5�e)��izzZ�L&��cY�2��FGG�8N��      ��!p     @�E"MNN*������Z^^n�Pm���L&�L&���-]�~}ϭ�JE�JE�e)+
��]"v �V;F���'��/��m�d���������      �;      �M4��̌r��n߾��������[4}���jssS�a�q�B�@��K�� ��ѮQ����q}��þ�]z�g2���C�     ���     ��9���Y���kaaAKKK;F���lu�}_�rY�rY�e�q9��V��\�� ���Q�����}�þ�]z���v6�     �U�     �2�HD�����r�2t�����֖����{�[ݥ7cw��fנ#| @{i�]b[�^�a����	z      2��4      �N=t���޽+�u���^��~��]�~]���;��T*�T*m��]R#
t]�� ����	l�mkO�R������ء�m��ѣG���
��      ��;      �8�&&&���t��]-..�V�=V�E�Q?~\Ǐ��Ǐ5??��ׯkkk덳��]z5v�^F��a�4� � ��v�v�ڥ���9rD���T___��/
iddD�l��      �k��|     �PsGccc�f�Z\\<���$���������O������9ݾ}{�?��Vw�4�{;��ۃ�z�^�  :W�k{��|��<�q��,K�\N�f���{��8���e=       ��      m$
illL�\N��˺}��*�J�c�0e2e2��7��͛75??����7�z��R��R��P(Ը�S��=����vw �ۃ�v������m�a(�LjbbB���l(�˰=��)���      m��      mǶme�YkiiI�6t�^Fh��Ӛ��֓'Ot��M�������o��V��V�2C��(
ɶ��a�zp�vw h_������<���ʬ�����Ԕz{{��}D�Q��y�     �m��O�      �ml�V>�W6����n߾������
T,�ٳgu��---i~~^w��Q�V{���*��*�˲,K�PH��e��vw �����=�;�}_��2��8*
*�J�RN�^zzz���J�x2      ��;      ڞi�J��J�RZ__�ݻw����X�2C###Q�Vӽ{����a��r]W�RI�P�qi��m����˿�8/ t���;aK�����٥�O�V�PP�Ph�W.	R,S>�W"�z      ���      :�a��ࠞ={���E���tL��_l�V.�S.�S�Rѝ;wt��----��W�UU�UIj��]�[���+��� ��۾��S���գ��ܖe)�ɨP(httT�P(�	ۇi�J&�������z      ��     �#���jvvVcccZ\\Խ{��n�c�q�E�E��e-,,h~~^���o<����P($۶;"v��%x��ur�.����T*�B����qE"��'l/�M��\�?      t4w      t�h4���I�����ݻ�{�ncC�a����Ɔn߾�[�niee�s��R��R��09�����^��i��� A�}�q�Ġ]z�9���c�>66�h4����q=zT�l�M�      8��'T      �;rGccc���nݺ���͠�jG����fgg���ݹsGsssz���+�|�W�\V�\�i�rG�m�}�.��{�G���;A������_����_�BA�bQ===N׾�����f�N��>     ���*      ��4�N��J�������E=}�4��Jwww#v���n߾�;w��{��R�$I�K{�� t��!{'���>����~cS{>����(Q����500��2      H��(      �=�C�T*�gϞiiiI����� �������߯3g�46�/,,��g�鱻�j�.�-t���D� ������K��)jO&�*
*
���
zĶe���ɤ�������      �W���'      ����jffF���Z^^�����r�c����K��u��-ݻwO��6���[��Q��N����M�j4 ��Aڥ7�v۶522�B��|>/�q�����ae2e�Y�B���      Z��      ���8����f�Z[[��⢞<y�Xm)��X,�X,�V��޽{�u�T�T���a(
ɶm�B���������9��@����Wy=j�i���j��X,�l6���!��      ��!p     ��c���ɤ�ɤ�={���%ݿ����b۶r��r��\���ʊt��-mnn6����J���C�P�ҩq���}�-�D� �E=�����lg����=�46������~�$�˩��'�q      ���     �P�����̌��ǵ�����E����j[�e)��(���ZYY�ݻw�������W�V�UU�UIjlv�m[�e1z����a����1{��M$Q6�U"�x�α}�=��      w      @��8�����٬��ִ���'O�=V[3C�tZ�tZ�ϟ���V#v_ZZjlr�^��M�T(�eY��};�w�p��������[�=ϓm��d2�W����
z���Ŕ�f544��      `w      `�4�L&�L&���Sݽ{W������]4U�XT�X��yz�������Ǐ7�y��ʖ�P(���n�f�E���5�������?�z���۫l6�\.�t:}��n��m�J�R:z��zzz�      hK�      �.�����ק���F���ŋ����i*�J)�J����z���ݻ���ݻwO��6����۽Ĳ�h?�C���%�V���6�G�e)�J)��)�ϫ��;��:Roo��=�d2)���s      �^x      x�P(�L&�L&�gϞiiiI+++�D��[oo�z{{5==�Z����%ݽ{WKKKz��y��N��mۖeY:d�;�Z��=��0���)���ѣ�f�J�Ӳ,+��:�m�J&�:z��z{{�      ��'B      �>�����̌&&&���ݽ{��@og۶������$5��߻wO���*�J���ow�m[�m���{�m�u����v
�sľ��-�HDG�U&����[�?R}[{*���      � p      > [ݛg�vw�����ݻ����<U*U*I/��P($˲E�^�S���wf�vB�����<ϓi�J&��d2:z����x��u<��      �C�      |��V�b����U�������yZ__��Ғ�ݻ������<I/��r����,˒mۇ.x�n������و�?��y�?����Ɩ�t:-�4��``[;      �|�      @�ض������cݻwO���� ��4M��q��q�:uJ�JE��ˍ�O�<i�u]����н��������}����Z���9��}�W�{R:��m�#�f�m[�TJG�UOOO��       �f      ����_��������ښ�߿���ub͏�8�������$ikkK<���VVV�����
^�MӔmۍۋ�f���n�Н-�x�����~��Sڥ��wR��R������D�����bf[;      ���     �}d۶����J��VVV��������G;�Ѩr��r��$�Z����ZYYi\ꑻ�y�T*�T*�^����}�B!��a��=�"o�^�;��׃�wy�>^=h�,KJ�RJ&�J��r'���#G�(�L*���      �E�     ��D"���O�<���VWWU�Ղ���B�d2�d2�^F������޽{*�ˍ�J��J�R㟷m[�pX�pX�m�q����W����w���k�H�]�Ѐ��y�|ߗmۊ���d2J�R�	9�(
ihhH�������k      �b�      @ b��b��������������ÇģMf������fgg���=z��WWW����8_��T���3C�pX��4��[�ԧs�����n׿Oh���{�������C�������z����)�J)�J���?��<�0400�t:���!��      "p      d���ɤ�ɤJ�Rc����fУH�a��K���������C���iuu��������G"9�#۶
�ؤ�B�f{�'�u�z���wB���B!�b1�R)%�I)�=ޡq��kxxX��=       �      m#�(��+����ӧ���VWWU�V��@���R.�S.�k��ٳgZYY�Ç�{=���jz���+ö�Ɩ���w���AD�����zzz1{"�`;{ �Q*����zzz�      �k�     �6c�b��b��&''���#���jmmM�Z-�����^����X,Jz�	|}}]+++�m�?n���jo��y=z�B�m��z����"���ɤR������,�
z�C)
)�+�L*���+7       �?M      ژi�J$J$�<��?x�Q��4M��q�����J�������ѣ���ӧ�-�;E�e)7b��[BK�3�Cv�0��۫��jppP�DB��=�f���N��H$xe      �C�      b{�^�մ�����U=|��U�u"��FFF422�x��yz��ic��Ç���#U�UI�����|�cm��n�v#~'|����\ו�y�<O��M�XL������o<��Whh��=�Ljhh���      @��V      �ٶ�t:�t:M��FL�lD��b������F�����'O��ٳg��w��.��=
)
ɲ,�w`���j�ڈ�]�U8V<����b����b����0��ק��a�R)�v      ���      n{�^.�������U=}��ؽMtuu)��)��5޷�����u=~�XO�<��Ǐ���c�J�ƙJ��J���ǫ�e������[�k����pc+{�������p��b�XL�dR�TJ��=      �&!p      �p8�l6�l6���-���jmm�ؽE�Qe2e2�W�_.����s����ɓ'��ϟ?o�;�m��j��8�lۖm�l4ơS�=�k��pX}}}�WZ���������h�������~ihh�'        �;      p@E�Q��y��yU*=z�H���z��<�z<�"++����j����������_���[�n�B�P#v�m[�iʲ���N���|�W�V������9��6�X,�X,���d���������      <�      ��(�N+�N�V��ѣGZ[[Ӄ�n����B!%	%�7�+��z���?~��ϟ�ٳg�K�R��2�T*���d���z��=�7c�>?`7�p��Ư-�R4Uoo�z{{����x������gY��L&544�+P       ��;      p�ض�d2�d2)������ڞ�3�W8V*�R*�z�r��J�^��������s���8����:�0^	����MӔi���y���}_����B!E"�#���ޠGF��B!��q%�I�u      8��     �C�4��Vp�����S���juuU�r9����pX�pX�x���j���?���mll�ŋz���+��V����5��^��m7B�������۶���(���rCw$QWW��9���.uww���[]]]���ak�!�F�H$��500��       ��      ��0����499�'O�hmmM>ԋ/����m�������3�J���������j��J�������eY2C�a46:o����q���4Muuu��www7�vww˶���a��۫x<���!���=      �6�#�       vT��'&&������u=z�H�=z�o���q�=#x�uU.�U.�������U*�Ư��r��/^�hl�o��P������{�'�u��Ƴ9~o�G�PH��(
)�*�(�(���K]]]
��:r��	z|�˲400�����	      @�#p      �V�hT�LF�LF������Z__��ښ666��,�9���mmm�T*ikkK[[[� �������0���}����s�#�ݶ���7.��-
ɶmٶ�P(Ԉ��y%Z�D"�F��xo�h�����7^}       ��;      ��b��588��v���5=z�h���F��F���oW��v߫ժ*��|�W�R�뺪�j��jr]W�jU���z�R��x{�c��7�o�|����}�6l�~�v뿯��e5��8�L�l��P�q��[˲>jV`7�i���_�x\�DB�h4���ٻ�����<�ϩ��&��֊��hn�����^)�#!k˾p4���F�1�F�'��#@�6�#� �cc�N��A����@"8���
'�fe�w��,������]=;Cv��"��
�:u��}8=��S�   �;L�    x)�Ow��:���y�w�}-��|��GΧ���k������z��r��{�/į��E��r��i��v/�;/����|����;��:w�`0���Q>|��}�c��    ���;    pm����t��������Y�<y��O�����}b�����2����������g�M|�     Qp    nHQ������^>�O�i������ӧ��i6�p�3���(GGG9<<L���t,    ���    ܊�(�������|��H]�9>>�(����*�l�`0���Q>|��}�ci�ۛ�    ���   ��h��y��a>|�$Y,y��Y�<y�'O�d6�m8!�����rpppQh��z��    ��    l�������ky�ג$UU��ӧy��I����\.7��n��z9<<���a>|��`��H     ��    l��h��h�����L�L���ٳg9>>NUUN���Arxx�d4�(�M�    �P
�    ��02��<I2��s|||���N�9EQd8^����7    ���   �;�����^�k���$��:���y���E�}�^o8%��(�"{{{9::�(�w:��    p��M'    p/���<|�0>L�����I�={�������,���x1;;;y��A<x��������jm:    ��Sp    �v�����]\���9>>���n�;��Χ�d?{{{�F)�b��     n��;    ����zy����k�%I��IUU����q&�I���pR�U2.�����   �W��;    ��*�"�������w|�w$I�����Ť����,�'�^�w1�}?�v���    �5�   ��W;    IDAT ��n�spp�����k��4�����9;;�x<�|>�`J`�E�~���������~z�ަ�    l5w    ��02�m��m�V��E����,UUe<g�^o0)�	EQd8f?����F���7�    �(�    ��N��I�MӤ�����^�ޏ���\.7��N�n���~^f���M���t4    �{A�    ��E���������t:���i�����Y&�I��J]�J
|�v�}Q^?�����~���h     ���;    ��>��/&����e6����4��b)����t2�Wf���)�b��     ^9
�     ����������w]_�V�*�WU��d��t���p�u:�w�G�Q���~�    ��Qp    �2�N'988x���r��tzQv��|>�PZ��[�yq��1��n�7    �KPp    �#��n��n������z��|>�d2�l6�(�O��TU���7��W��J���p8L��W�]�    �~Pp    �Z��E������(����g�Y��yf�Yf�Y���Rû�������G��{�$�^���(6    ���    p�EqQ�V�;����|��ju���oΧ��?���}    ��M�    �� n�X\��ϟ/�,�����,�ˋ�M��bz6�(�t�����|��yy���n:.     w��;     �r^X���������(���}^�?��Z��D��J��I������Ey���]�>/���.�bӱ    �G�    �VEQ\��/���V��������r�L]�Y.��z�Z��^�S��+_�/�"�v�����v��v�n������~~���Vk��     �8w     6��n��n����>��뺾x�^�/&�?��y��k��{-�ˏ�\~^8�N����?/�?��þ����	     w��x    po(z    ����          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(�          ��          �

�           lw           ���;           [A�          ����          �VPp          `+(��s��"�ժ��          �2��)�E���tnPg��~M�d:�f2�d�\fooO�         �;m�^�ɓ'�t:�i����o��SUU&��O�          p/�V��������������n:�D���k�&��<��$��|�q          ���f��f�t�݋��EQl:/A�����:��,UU���M�         ��Y.�999�x<�`0�h4J��*}�S�cΧ��f�MG         ���4M&�I&�Iz�^��a����cq
�w�z��t:5�          .i>�g>���je0dww7�Vkӱ�
�[l�\^|��eE���H          ��V�y�u��:UU�����������(���5Pp�2M�d6����,���K/���c         ��d6�e6���ng4e0��eܷD]ש�*��4��z�q          �ު�:��8�������F�v���E�7�i����L&����;����wf��Wo�kTU��;��/o:         �}���}m����6�㲚�Y&�ׯy�L��L��t�������<�+Rp߀��3��RUU꺾��>}�]I����&~(          ܼw�y�{����qYEQ<�����eNNNrzz��`��h�v�}�G��o�����l��(          �X�ש�*UU���e8���o:�+C������L��[��          \��|��|�V���p��h�V���X����Y,�L&�N���1O򗊢�W���d          x)����R�7��6�^��9;;KUU������ٹ���FM�d:��w�ɓ'O6Yn�j��8ɿX�姚�1:         ���)��ǒ��$o&��[�;�'O���=UU� ��e��5��:UUe:�f�^o*�:��\����ղ,W�
          7�,�q�/&���?��߻^�?��G�to3�j��x<���i�AF�Q:����j�&��<��$��|�Q���J�_(��o2          ܦG��z�-��OE�G������K���i�L&�L&�t�݌F��یp�(�_Q]י�f��*u]o2ʯ��<��˲�l2          lRY��,ɟ)��g��kI>������c�\���8���b�{�ݾ�w���%�Ok��f��1K�V���=��          ۦ,�u�/'�rY�ߕ�}���6s���TU������2�������վ�����!��u���6Lk������M��RY�O7          ,'�[_��?{��4M�$��m�����i���F���B��,��L&�L��4M��u�_K�eY��$          wէ?��y�/%���?��߻^�,�J2��u]g<����]S�y7�oj�&��,UUe�\n2�?M�+�N�x����           p�<z��ד��3?�3j6��p��$y�63���g�Y��n��a���������NUU�N�Y�כ��w����o��o�+o���F�          p����['I���ʲ�}I~,������2'''���F�t^��+��7M��|��d��|��('I�b���£G�~s�A          �Ԕe��$_.���E񇛦�I��VC4M&�I&�Iz�^��a���mF��T�����f�TU���7�ד|q4���}�s�&�           IY����ϔe��EQ�@�4?���%)n3�|>�|>O��N���h4J�ݾ��J�ϧ��f��eh�&��,��������܏o,          �-�e�H�$_��g>�f�����p�V�u�9�NUU�꾳����վ������z}1�}�Zm,�j������u������          .m2�|�(�������gww7�n�V3�ڞ�fi���F����~�
���2��$��4M�l,��S�7�          x9M�d:�f:�fgg'��0����K�u]g<���4�� ��(�����ߋ���S	ggg��^�u��i��J]��          ܌�b��b��x��p��px�%�i2�L2�L��v/r�w��Z�.������X,��ʴv          xE��뜝����,�^/��0�~�֧�/�˜���k�{�ݾ����ܛ��|>�d2�|>�X��z��l����\.7�          ج�|��|�v�}1M��K���:UU���w��;Sp����P^���r�O���ʴv          �B]�9==���Y��~��az�ޭ�x�p?�2�j�n=ǋ��������l��M�d6�m|j<          �����t:�t:M�۽��^ŭ��:��8��x�����ʂ�z���־Z�6����i���zc9          ��i�\���$��8�� ��(�n��s�f��f����`0����elU�}�\f2�d:��i���8�?�N7�          �?���d2�d2�����J�T��t��V��$M�d6����l�����u��i���R���r           ��b��b��x<�p8�p8������n��������[��A6Vp_�VS�����bd�Xl��x          �ղ^�svv�����z��F��z��Lu��YZ���T�v�}���j��i����L&�����<�}9��i���r��X          �$������t:S�[�֭fX�ש�*UU���g8fgg�V��Rp��:��,ggg��~>5~2�l4          �Y�V��9==M���h4���έ��f��f���`p+��-��Ok��f7ẏ:�_U�F��          \V�4�N��N�����p8L�߿����-����ӹ����^�3��RUUV��uoiu]g:�����u��           /c�Xd�X��j]Lu�v������}�۽��^ŵ�sm��r��d��t��i�k�+[,��*��tc           ��z��d2�d2I�׻(�߶�r�������f0d4��n_��/Upo�&��,ggg�������r��           �a>�g>�g<_{�����u��JUU��~��R{�P����TU��d��i����bZ�&s           lB]�9;;KUU������z���p�n�3�2Sŕ��R�}�Z���,����]��i2�N3�L�X,6�          `[�����i��n�����_F]���9==�h4�h4J�պ��K���u���6:�}�Ze2�d2�d�^o$          ��[.�999�x<N�����n���fh��b��p8���ޥ��Zp?o���ۛ��|>OUU���~>          �]��T�������[���4M���l6���~������-�u]���8����C~��z��d���R����          p�,�,����f0d4��n���u]�ٳg���y��AZ�������|�gϞ�����bq�����x          ����뜝����,�^�b��m��fY,988H��{���+��������V�%�9>�}�Z�ڹ           ���|��|���Ӌ��mLu_��y��i���3����E��i��������$����nZ;          �f�V���㜞����g8~�t��6�S�u���/�]�o���4M��i&�I�ō�          ������i��nF�Q�A����3��JQ���K�͂�t:��r{]יL&�L&�����          ��-�����$�� ��(�n�F�:;;K��M��Og�^����F��穪*���F�          ��4Ms1���e4���]�T�������svv��i�u��j�������k�          �͘�����v�988�։���:UU�5�ͮ��>�L���]�          �Z.�y�wRUյ�;���V]ד�ڰ��_�Dx           �G�4999�����Z�f�$��:6�����ױ           w���i���um�OZI����^�Mn          x����������Z��_~�]&��u          �Y��9;;���~���ѣ���_f��dra           ������n�ώ����V�&ɟ}�]��j�z�0           �Q��:����E�����o���$��"-��          ��P���.����/���$eYN����u          �ղ^�_t�ʲ���7�I�4�/'���Tŋ�           ��x�n��^����/.
�eY�����Uwk��/          �{���\yMQ��'~������o>~��L򗮲a��Vr          x�E�n�{�e��{��{���Z｣���x��U���          �����)��*K�$��7ި�������o����(>{�����Un          ��FW]�seY���^|_�=I?~����ew�t:/          �;���ggg�*K~+ɣz��I�$,��/{���^:��UB          p����\e�"ɏ�e9��7�U�=eY�n��7����j���0�ַ�          �{�����ϕe��}�7?t��,�Z����I�n7���)��
�           �k������+��?��>�*����d��v�{��UG�          p����g8^e�?���8I�a7}d���7ި�|*��\���`������          �1����{�%O��[o����G����$)��i������/�`ww7��買          ���A<xp�%�$?T���_���$�=���(�`��e����g0\�v           �T������U�4I���,��e\���$�?�EQ��$���_E����r           [������0EQ\zMQ�QY��r�s�TpO�Ǐ��$��B���0;;;W=
          ��t:9::J�u����<~���z֕�IR��K�^���(rtt�N��"�          ��v;GGGi��WY�ʲ��9�
�IR��[I��K�j��ÇWm�          �/8��H�G�4/r�˴͛���o&���.h��J�           [����v���M��eY�^�ܗj�����$�N���k��nS��          �988H�׻ʒ�I��eY��̹/=J�,�I�H�.��������e�          �����g0\e��&�7ʲ��/{�Kܓ�,�w:���&��e��<x��:�          ����eww�*K�I��,���:ο��{�����_I��$�.�f4]��          ��ë��I~�,����2\[�=Iʲ�?Z��&�]v���^���u�           �
��~R�e���|�,�/_g�k-�'ɣG��VQ?�����EQ�������          ����������.��,����r��$y���_M�'/{Q9<<����M�          �t���պR���eY~�&��H�=Iʲ��$���E����t�ݛ�          �7���)��RY��o*Ӎܓ�,˷���e�o�Z9::J�ݾ�T           ���n��I��EJr��$�믿�f�_���            �PE�����v����F�)�ruS���/��7ި���?���^vM�����Q����d           ���(rxx�����,��$����}���XneL�g?������$��ˮ��������          x�<x� �~�*K���eY>��H�r+�$�ɟ��'I�7�W.���������B          �"���3���$�(�����>�VpO��,��V����<���p����L r �e    IDAT         p��F����^e�4���e�o(��Ղ{�<z��7���$�ˮ����h4��P           ��`0ȃ���.��SeY�������z�=Iʲ��I~8��k<x�~�s�           �^������,i��x���ǿzS�>�F
�IR����O\e���az��%          �?��nS�U������_��Lec�$)��I����_E�����vo0          ����trtt�V�J��_,��O�T���h�=Iʲ|��?����%�v�}��           �v��"������ɛ�tY/�'�믿�&�˗���n��ÇW�4          ��v>P���\e��L�#o��F}3�.o+�o��F��������ˮ9�_�&          �����n�*�~#��e9��XW��$��g?;���ߟ�^v���N���n0          ��ppp�^�w�%�w���7˲<��LW�5�$y뭷N:��'����]���rppp��           ����~��U���n��O��O�ӛ��"����$o���W�|2��ˮ���߿�P           [jww7���WY2i�Z�����2���+�'IY��g���d��k^�          �N���ۻʒe�z���߻�H/e+�I�����������{��^�\7��9C&��"�4KcEQlZȀm��$�ٹ9�Pl-��VTP����z�"�Q�x1�H"�M�&xם�q33�������n���=gv�׼�k�����,��L�\��;]�}c�;�����m?V          �D��fY,�nӓ{I��Z��g�.e�$Y�����o��}�uY,��fC�          x�vvv�X,����=���f��Q:pO��z�c]׵M߿��}?�*          �Gc2�d�Ze4�*���z������ܓd�^�/�n�~4e�Ze2��
          �x���9sf۸�g�\h�Cu"���=��o����          �������m�>�Z���Z�;Ԯ��������ߒ�76��          �A�uY�V��~��'y��n4�;Q�wk�f�'�|tӛ��\.�u�p�           �u]�Evvv�9�Ӿ���Z�1Ԯ!���=IZkג�5�'7��N�Y,Í          ���Qvww�9yv<?q���g��4��'Ik����\��fww7GGG�          x��������$_}���4iP'2pO����'�<�����~�          �<@��B�w��>2Ф����=IZk������f>�o�           �jww7GGGۜ�M�-���4�X���=I���/'yg�{���.GGG��f�          x ��4��b۳�j���{�Ӊܓ����]�]��}�uY.����r          �V���r�L�uۜ������8���=I����$����.��*}��
          `3��8gΜ�h�U��ӭ�KCm:n�&p��;��ܦ�G�QV�U���           ^����I���������v7�7'��Mo��qV�ն�           ��>�{2�ls�����oh��jףp����Iޑ��6���>��*]�7          ��t]��r���9�x�'���<?ЬG���I�Z����?H�Movvv�\.�          �E�E���6'=�L��Z�:ԦG�T�Ir��ſI��$����fY,Í          ����(���ۜ|f4��ҥK�jӣvj�$i����h��$76�����|>p          ����������h4z�ʕ+jS�:pO�+W��n��M�¦7�          `#���988���Ů��ʕ+�9Ԧ*N}��$��_��'��������          �f�Y��e�������X�׿0�2��=I���N���ﻮ�b��t:p          �����b���뺶^�p�I�<6�{��־7ɿ��}�uY.���~�U          �i7�L�Z�2m�p��z�~�P�*z��$i�}W������h��j��x<�*          ������$�t�Ie=v�{�{�Ν�'I޿��x<Ι3g��          <�^����d����|ck��@��z,���������}G��lz3�LD�          �ƺ��j�J��ۜ��t:}kk�C�챭��z��;;;_�����}��b1�*          �4�.��";;;ۜ��d2y��}������6pO���~���x�D�g6���fY.��          N�������ns����-�.]���6��u��$�/_��$oKrcӛ�������F          '�|>����6'��Fo�|����x��$i�}8�ۓ���f>����`�Q          �������i��䛮\���M:Q����>�u�;�����~�          8�vwwstt��ɽ$�j���@�N���Y��?��M�w]����L��W          �M��,��n����Z��&�H�/�Z��$߿����Z������          ��&�I��e�����G����j�I%p�Zk�N�S���.��2��x�U          @5��(��*��Vi�K���t�	ܿ�{Iޕ�W7=�L&Y,���          p�-��L&�mN>�Z����vw�M'�����^H�5I>���t:�|>n          P�|>�t:�����|݅n4�������g�<��O6�����l6n          ��M��ls��I��Z{n�I����5��>��$�g��]�e�Xd4�         ��h4e�X��MO>5��h�m�$?�T�h��Y��J��OK��          8}���2�7}��$O^�|���tj�7�Z�X��O��&�g�Y����          ��l����M����k[kpҩ"p�Bk�ג|k����?<<��'3          �º�������u]�������t�ܷ�Z��I��&oG�Q�����          ��0��3�L6}���z�SC�9������I��&o��������          �!M&����o���Zk�?��J���ZkO%��M��          �|>O�u�<�/I�xΩ%pp�Ν;w>ɯ��Ý��L��c�          <l}�g6�m���;w���������ϟ����|������          ����&����I�q�1�	�_��ڍ$_��#��ngg'}��(          ��Ǜ|z��$y�����A���֞����I��������"          �a���{�Oo���d������t�	���/>�����|��L��t��          @����O�K�.��1�9���ŋ�&�W&��/���<���*          �AL��E������}���O�SO����֞[�VoI���ק���<	          x �W��/�f���x��3�:�1�J�p^�.�J�/Zk�����{�k{{{}d�          �������ݻw?�o=�u�����Gզ��'�����I����N�[I��l6��G�
          ����Ə%��$L�/���rq��|���Zkג����          �������G��q��          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�<� �Jn޼��ׯ�ڵk�~�znܸ��7o�Ν;�y�f��֭[�s�N����Ͻ{�^��L&��fI��t�����go?]�e?���~�}���       ����_����_�u�ƍ\�v-Ir�ƍ$ɝ;wr�֭$y���|�������w}�g>���� ��<���/���� �۷o��g��իW���=������۷�}�t:}9v?<<�r��ٳgs��ټ�o�ٳg�Z�2�CP       �W���|&W�^}��x�g��O����v�Z>������h�����o#^����ٻ��:�������#��f[�ٖ�)iI>)�d���L�L�L:�N�_2��	�f��%� �HXLk�=8	ƀ��1���}_�~t�s�H�+ɖ������c���[��#ٺ���z w �-�٬FGG��۫��>���̼��+&��D"�D"����y�q:�����y�khhкu�v�ZUTT,�j          �R�F����Soo�g�cccJ&�K��9e�Y�A���>W\\���ڙ��ڵk�v�Z555�L� �j�	 �i�hT���P�������=s4�J��d4::����Y��^�֬Y���&�Y�F���jnnfG3           �\6�����L6b:'188����nV8V8VGG�ק�655���u&+���$�0�h� ����; �d2�����x�.^����ɥ^VΈF��p�.\�0s�0555���M�7oV[[����p�           �Z��.^�8�����T*�Z�e�?x��ə�EEEڴi�LFbÆr�\K�R �rD� pU�x\===3��.(�.����4��߯��~<xP���8�    IDATTZZ�6���U�7o֖-[�����+          `����W�#���W�dv�D"�:uJ�N���I����ڼy�6oެ��vUUU-�* ���; �
�lV�.]ҙ3gt��i^�lu��ə]�.�K[�lѭ�ު[o�UK�B           V�p8��g�����:{�����R/i��d2�����P�����|�֭[�� ���; @�PH}��N�8�S�N)�,��f�����Y��N�$)/��9��k�C�lV�^���9�NK�C�?�J��5��RH&�:{��Ξ=���~Z555ڱc�v�ء[n�EK�6           V�4��ݭs����?�G}�L&��˚1W>b:1���a\���CMӜ�Ed2���l6�t:�t:�T*�d29��KixxX���ڿ�\.�6oެ�۷kǎjmm]ҵ rw X���������������Y�)�n�[�g���VAA�\.�\.�Ǣ�e:��H$���ǕH$���ǕL&���ؘ<��*??f��wܡ���EY           �]"��ɓ'u��	�={V�PhI֑���������t>��v��r̈́��t~:1WFb���dR�Νӹs�g������[o��߮m۶-jn �;��*��߯��{O��������������UQQ�
UXX(�0uW�p8�v��v�URR2�i������Ԕ�Ѩ"���Ѩ�ɤ��J�R3/s�w�VSS���N��_��***l�          �r�J�t��Y���{:~�������v:�*,,��FL��bد�0��	����s>�H$f�SSS�D"��b��mttTЁTTT��n�Mw�q�n��V9�N�� rC���	 ��t�������g^^�JJJf~*??Qz��0���~uu���t:�h4�p8�P(�P(�T*e�:�g��ݻWmmm��;t�w���ܶ�           �?�����6CEEE3���+�ǓS��n���?�g��L>"+ںy ��ȑ#:r䈊��u�8����nc�; �p�`���:t萎=���~����nϼ���������Sii�JKKg����{(R4���i��p�.\��ݻwk�֭���;u�w��v[�          �\b��>��:tHǏ��Ԕ���N�L>���T��ūj��t����H������� �(�d$LӴ�w8�	�WTT�3������/�����^ ���z҇��Ν;?��m�ױP�hT�����z��c��>��C<xPǏW&������Tii����T^^���B�z��dR�@@>�O~�_�tڶ^��g?�/}�Kjmm��           K!�����k�����>[{���B���*))YU�nD&�Q0�����u»$����K_�������x<��V����L0���v��v��Y�ԋ����v ��l~�_��o����q�����B���*--��&���P(4v�c�����V�y睺��;��zm�          �ݺ����o�ȑ#J&������SYY�LF��r��g��F�3a�p8�l6kK�7��;rU�R/  p�L��ɓ'��o�̙3�~�_YY���j��c52C���*--UKK���&''5>>�P(di���.uuu闿��>�����_�2/r          �e#
�w���<���Q[z8�N������JUUU�������USS�2��|>�������d��e}b��<��j��������}�sr�ݖ�  ,� ���R)����ׯ~�+�����̼���Wr��jhhPCC�b��&&&466���)�z��q���[z뭷�y�f�������/�B�ò           XettT����[o��D"ay}��qE�������t���Z���J�R�����Ą���a���Nuvv������^_���TQQaY} ����2������
�Ö����SMM�jjj�/����Y�Fk֬Q$��ؘFGG�N�-�q��]�pAuuu��W��/~��          �	]]]z��Wu��Q[N�/--U}}=�ڗX~~����TWW�D"1����b�����������o�3�������i�ڵ�� ؇?�W��;w~(i�R�c��Ѩ>��O/�2��022��^{MT2���~qq����U]]��;�M�T&�Q:�����d$I�lvf���?�p8d�Ø���p8���wů\~i5MSV0��~ii����/�+_�
           ��4M�<yR���.^�hy���|��Ԩ��^�׷�t>��f$��M������6cV>"��!�`P�������e���͛���}M��ԧr:+,����L0�Դ�k���;wV.�"`/&�@����/���'OZz���i����*,,����0MS�dR�DB�d�_�/jv���_ӡw��)��%��%�ۭ��|��n�\�%{�3c戮X,������*�JYR?�^Я�k}�_�׿�u���[R          ��d2:tH���FGG-�_VV���zUVV.y��4M���Y��D"1k؟��4����?g>��tھ���VVV���2�_�^###�t�����---��7���o�}�?7  ��;�*�w`�����/��cǎYl�x<jhhP}}���M�T<��Ԕ��b����e!�Ő��'�ۭ��y<���,��l6���1X�"'�a���wީ��Keee��          �4M;vL���/5<<lim�0TSS���Fy�^Kk/T2��"�ǕL&-ς���p��v���p&#QPP�$�w�4���o˩�k׮�7��M��_�%Aw�JLpG�b�; ���A����:z����ʋ����Դ���M�T,S4U4U<W"�X6/j��1�F���v���x��zUXX(��k�k�á��:������i``@�PȒکTJ�;Ｃ/|���7����RKj          V/�4u��I=�����v^^�������(��ei�I&��D"����	�/�I�v�f���b�����_��(**�}(�a*//Wyy��ᰆ��4>>nY���O=��6mڤ����ן���[R ps�r�
0��]���z��u��!ˏ����PSSӢ�3��L�=�(�-����a�


��z��zUTT��<����B!jbb�Һ�G�7����K��          ���;wN{��QWW��u�n�̉�vO�Ӂӡ��tr�


f�-��x<���A���X�Oټy���.m۶l�v�Ma�;r�U��;�{����}�Y[�����Z�n����-���L�T<W8V0�5����n���T��ŶNx���R__����-�[TT�o|���W��(�}          ������g�Qgg��u�����Ԥ��F[�L&�g~Y��Xi���U\\�������:�=�J���_��Ö�o����?��֮]ki] �pG�"�
prG&��믿��{NSSS��.++Ӛ5kTVVfi�i�LF�pX�PH�`����p8��zU\\���R��n[���a���krr�Һuuu���G�q���          ����ڻw��y���iY���|566���і�i��D"�D"
�B��b��X-Ð��QYY�JJJTPP`K�d2���~�'����}�s���g���ZV�%ܑ���܁�p��9=��S��nII�֮]���rK�JR:�V ���gJ��


TVV���2[��PH���
��ݶm���_����          ��DB���Ӿ}��L&-��t:��ب��&9�N��J���a�����r���Teee�z��׏����Ȉ��*�^����������oY] pG�"�
p���Аv�ޭS�NYZ��񨵵U����YM�}i���\eeer�\����|���tw����_��_�[���JJJ,�          X^L�Աc���3�hbb²��a���Ak׮U^^�eu�C�~�_�P�P�"s��*++Syy�<����Ѩ������-�[__�o}�[�x���;r�U��;�4�Ѩ�}�Y��曖�9�N555i͚52k~7MS�@@����D"����+,,TEE�***,;V�4M���_�tڒ��TTT���K_��m9          ��:::��O���˖�-++����UXXhYͩ�)MNN*j��g&a�&���Iuww[:P�n��V�˿��,�,��U�W���;q�~�����YV�0UWW���Ų�މDB>�O������a-�á��UVV���ؒ��tZ}}}��X���f�����Z[[-�	          �M�DB/���~��_+��ZV��񨹹Y��Ֆ��f��������<������"UVV���Ԓ���ijxxX����fc�N���կꮻ�4�,6��U��
 
z�'t��1K�k������MӜ	�OMMY�:�-��*(���@���7=�=//O������Qgg�B��%k����w��}��_�?��?(??ߒ�          ��r��=��������Ԛ5k���dI�9��Lk�2�{���p8�p8,��5�����ajhhPUU�zzz466f� �L&�W^yE�N�ҷ��mmڴ�k �ȹ���>�����j�z�J���ظ�� ��i�:r���>uuuYV��tjݺuڴi��n�M��d2WOO���R��E��bJ��
�BW2���㹩��.�Kuuu�x<
��ę��.��ѣZ�v�jj��A          �k�F�zꩧ�{�nK땕����]���7n�B������b���'�cqd2E"���kjjJn�����N�S���*))Q8�l�{0ԡC�������� @,;�P�L$I%K���{���_�E�^�WFGG���_���o�L&-�[ZZ��[�����^ܒɤFFF��۫p8̎��4M�b1MLLhjjJ.�K.������F�X̲�آѨ�9���������           K���Ӯ]���'�XV��t���E6l��p�i����TOO�&&&���$	MNN*��t��v�p���񨮮nfZ�U���t��Q566���β����#W���W X�L�Ծ}�����[�R����������T�=�htt��oƑ�B��B���^�jjjTZZzCu�n����5>>���NK>��O78�����o��n��          ������ӟ�T�N���nee�6l�pS������511�L&c��k�Ѩ�Ѩ<����UQQqC��á��UVV���S�HĒ����k׮]����+�ۿ���^�%u`5b��*�w�z���������[oY:���B۶mSii���#���1[VN�G�K�R

���ϗ�㹡:^�W������'��������i�����c�          ,Ǐ�=�ܣ��^�j��婭�M�֭��yc�t:���a���)��4M�ևܖN�
�����p8TPPpC9��m�4���^���;jmmUuu�eu;0�����*@��ֱc�t��jppв�N�S���jmm�����Ԕ���5<<�1[�\:��	�����P���t���Z
��E@WW���}������ܒ�           �%�I=��3z�g�H$,�[ZZ��۷���Ʋ��LF������%ؾ�e2�������2���)
)�N[��X,�Ç+�h���r8���F�����*@��F,ӓO>�={�X:���P������ݤ�x\����t�=
)??_n���kx�^UUU)[�y����o��t����O+           أ��O�v�҉',�i�����q�����f5>>����B!��1t�r8�x<םEp�ݪ��U2���{I�|��Μ9���v[V�
w�*� w��utt����u��9�j����:mݺ���ǩTJ������W<�l]XyR���~��Ѩ
��/
���U[[+�á@ `ɚ�٬>��C]�pA۷oWAA�%u          7�4M���k����/��oY]�ǣm۶������Ǧi��󩻻[�`�`;�N�
�TPP ��u]�p8TYY���Be�YK������[o���@7n��&`��U�W���3MS/���{�1��a�����k���jjj�����Q���Z�c+_2����2�������s�0������L>�ϲ����1>|XMMMjhh��&          ����~���z�7,���$���i۶m74�/����ҟSc�K����|����z�r:�/&YXX���jKO��d2:s�����g�g���B�����*@��1�XL?���x�Kw�i���7t�P `G2n��Ԕ&''�p8TPPp]Aw�ǣ����a%	K֓L&���*�Lj۶m׽�          ps.\����[}}}��4C���jnn��'�I���kxxX�tڲ5au��㚜�T6���뽮�ü�<���(�J)�Z����A;vL���*++��.p��#Wp_�ׯ��W;w�ԥK�,�[[[��[�*??��>.����[����d2��	�S6�U(R(��㹮��N�S���J�Ӗ�lp��utt��nc�2          ,���?����Ȼ�nm۶MUUU��q�ijxxX�����㖭��i��F���|���WAA��?�0UVV��rY:�2��СC���Tss�%5�E�����*@��>G����߯`0hYM�0��Ң�����j�������۫T*e�z�i��r%�I��p,���PEE�


,{�ѻﾫ͛7����          ��R���q����f���-))����UXXx]�D��եP(d�Z�i�lV�`PSSS***�ӹ��dQQ����,;Q ���>����-�ܲ�`5��U�W���d2����ݻ-���r���ޮ����2�~q���O,�������Y��y�^������[�u355�#G����\---��          ���Ą���<y�Һ���ڼy�����1�LF�T{�.�H�����t^�&�ۭ��jE�QKO����G}�[o�����V!��\E�} �\[ н�ޫ�G�ZZ���jǎ�z���l6���!��E��f�{����VMM�����ɤek9q���v���Ne          �ș3gt��wkddĲ��ahÆZ�v�u�l��եh4j�Z�k1MS�PH�PH^�w�2�N�jjj�H$,�����Б#G���z�4��E�����*@�����>�ܹS}}}�֭��P{{�\.ׂ?&
���S�p�ҵ �cz����Z��`��9�S9�Y����}��G�����v�-�          �������c�)�HXV��tj�֭���^�Ǥ�i���httT�lֲ� �#�JirrR�C���ڜa�***$�!�c�D"�w�}W���jnn��.p-ܑ���܁��;wN�v�R0��nMM����<�4M���h``�7��4��U\\��	��C����d2�nҘ������u�-����ز�          �Zd�Y=���z�d��eu].��mۦ���L8VWW���Ӏ���U\\����a*++������k*���>�i�ںu�u�� �(��U�W���~�����V2����aZ�f�֯_��@�$��quuu)X��*�x\�@@:��0���+??_~�߲uD"=zTmmm�����.          �t�DB?��t��aK�jǎ*,,\��ijhh���I�T�O��z�*))����s��?��ؘn��珀E�����*@���i�z��{�nKw%���7���i�;(�����ӣT*e�: �e2������]��wqq��^�&''-[G2��ѣGU__�5k�XV          V�@ �]�v�����-++ӎ;������c��:;;
�,]`������JJJ���x<*++���W&��l-����x�n���$nw�*� w��R��~����^�����P[[�jj����d��ݭ��	K��)�(���dAGr�������l6���_�i����    IDAT���ݲ�          ��h�Ν��nyy��m۶������Q:��t�]�O�/**Z�&�˥��
�|>K?����t��	}�S���뵬.��#Wq~�U#��{����y�K�:�Nm޼Y���z>��ҥK
�Ö�XSSS�x��?+**�}���j����z��S          `�8����?�C���֭��R{{��&[�����>�],;�DB�.]Z���ڱc�
-]������勉��Һ ���X���v�ܩ.XZw:�^YY���}>�._��D"a�:�ŔN���ե���=_ZZ�m۶)//��u�߿_�<�G|         �rw��)�{ｊF��֭����͛nO&��t�|>��k �i����W__߂6i��nm߾]EEE��#�?��?��ZZ rw +^ ����=���XZ7//O[�nUEE�5�5MS������S6��t�R0MS������Z��tII�v�ر�����ѣG���*�JYZ          ��'N��T2���n]]����n�B�x�b���k ����ӥK��Mp�\ڶm����-]C"��}�ݧ3g�XZ rw +�������絛��Һ������k>�N�u��eˏ�rA(ҥK�t*�������-��~��	=����          ,'v����ƍnQWW'qcŉ�b�x�"��5���Ϸ5�����[Z rw +��А����jdd�ҺN�S�7oVii�5����t钦��,]�K�?��7rw:�������ڵk           �J�#�<by����Z�ׯ��s�i������K��:;;511q�g������.��k�z�!���ۖ��\C���400��;wjrr�Һ�Cmmm*//���pX�/_f�4V�L&���N�|�k>[TT�m۶Yr����_��_
�Ö�         �\v��=���2M�Һ���jkk����L&�����~K���4Mhpp��NOr/,,�t�lV?��u��K�@.!�`�����w��]�_��ЦM�TYYy�g'''9r��i��������5�-))і-[t��������w�M�         ����/�'��<�^^^����&�I]�|Y�h���@�WOO�5��\.������x,�o���|�I�߿�Һ �+�XQ����k�.E"K���6�����ώ�������G`�V__�5��"׫��[�����          +�o�[=��s��---U{{�5�;55�K�.)�[�`9���� L�ǣm۶��v[��4M=���z���-� ���;�cxxؖ�͆a���EuuuW}�4M���jxx����r������u͐{ee�6l�`y����s�=�E
         ����ڽ{��u����m۶k�ۃ��:::�N�-_��D�Q]�|��_ڲe����,�o���x�	���[����F���011���[�@���uuujll��3�i���G~�����r�u���k�T���Ӛ5k,���%�w�}J�R��         �����o��'������V{{���G��~�zzz��f-_���q]�tI�d������_c��4M=���z��w-� K��;�e���i�Ν��vUU�֯_�gL�TWW��������njjjA�q577�������ϟ����O�         ��p��1���?��i����tj�֭r�\W}nrrR�������d2�˗/_����
���^���f�裏�ĉ����B���
�t��wktt������ڴi�U��4MS���
�Ö�V�X,���6nܨ��R���9sF?����         �\v��	=��Ö���0mٲEEEEW}nbbB�����V�T*����b��>W__���F��g2}���י3g,� ���;�ekjjJ�v������=��l�"��9�3�lV�/_V$��?����q]�|���q���[����������~�0E          ��t��9=��C��Z�~���˯���ؘ-�`�I���������U�knnVMM�-�|�A}��'����D����N���������yyyںu��n���L�ۯ��(�?J$���P*������<���+//����֞={,�          v�������՟�ި��&���_����QY�X�2��:;;��+2C7nTII�������>6� X��XvL��O~��?�����<z�ޫ�����qB fK&����P:������mٲŖ����Ӂl�          V��|�����H$,�]^^����>311���a�{+�t��j�"�á͛7_u獊F���{,� ���;�eg�޽:r�-�TUU5�}�4��եh4jK`5H$�����yeeeZ�n�-��z�)�8q�          `�X,�{�G>�����G�7o�a�>399�h�&L�ܯ�A��vkӦMr8��r�����{�e� ؍�;�e�w���^y�[j������e���i���[�pؖ��j����ѡl6;�3k׮Uee�彳٬y����X^          ���d����������S�����}��󩿿����j�N���ѡd29�3�C ����Fuuu顇�j> rw ��������ܖ��Gmmm�~�h�����
�l��F�XL���2Ms�g���TPP`K�{�G�����         ����O�ܹs��޸q�����	�J�R���P*������FUWW���ԩSz�gl� v!�`Y���׃>�t:mym�áM�6��r�������~�彁�.����{ސ���Ԗ-[�t:-�����k�.MMMY^          nԋ/��7�|Ӗ������~8VOO�U��~�dR����NR7C6l��뵥���������R �@�@Λ�F�Q�k����f��������S��B!�{���j����������?�Q\          r�;Ｃ�ޖ�EEEjmm��~<'��(�����C ���l(I�w�։'l� V#� �e2=��ö�������0��@ ���![z����	����{�����Sn��ӧ����R          ���G?���l	�;����0�9��iuuu)��X��E"����{������ٖ��lV?��500`K} �w 9�駟��lKm�˥6����F��% k����{���r�ݶ�~�Wt��1[j         ��D"=���J$��ommUaa��L�TWW��ɤ-�\���kddd����������w<�<�X,fK} �
w 9��ѣ:p��-��І��&�Iuww+����������F缗�����6[������G�R         ��L��#�<���Q[�WVV���~��===�����7���������y�0mܸѶ!�CCCz��Gm9- �B�@N����O�S����֪��r�{�lV���J�Ӷ�0�l6���n�R�9����і��R         ��}�Y�>}ږ�.�K7n����А���-�\]�"�Ȝ�\.�֯_/�0l����7���-��
��h4�x��c��^�Z[[����c[o זN����5�Nᖖ��{hhH�=���         ,�'N�W���m�7mڤ���9��|>�������M��0����J�����Ϟ=:{��m��fp�S�>v��p���UN�s��###
�B���p�XL}}}s�3Cmmm��R>~�8��         �nxxX�>��m����U^^>�x<���[�X�t:����,((��w6���C����R nw 9套^ҩS�l�_[[����9�B!���������������^aa�m�w�^}��Ƕ�         ��%	=����������Rss��2�������fm���LMMippp�{N�S---�����~�t:mK} �Q�䌎���⋶��x<󾼥R�y�EX:����F�s�knn�m�r&��#�<�H$bK}          ���ݻ���o[����+//o�{===J$��p�&&&4999���J����ֻ��C�=��m��Fp���y�e2[������9_�L�TWW;�d��zzz���4C�6m�����~����V         ��t��i<xж�UUU����������m�ܸ���yOuhii��岭��}�t��y����"� '������m����TYY9罁��b1�z�9�TJ���s�+))Q]]�m��;���~۶�          V�`0���G2MӖ�N�S���s�����/����f��۫l6;�^~~����e�-�M�ԣ�>� 9��;�%w��1>|ض�.�K---s���� w��aMLL�y���E�����~�'l݀         `u0MS?��m����*��=�z&�Q__�m}X#�Hh```�{555*//������{ 9��;�%599i�7FMMMs����i������u��g]��˛w���y�e2�z          X�^{�5�:uʶ�EEE�����^__�R��m�X������Ϻn�Z[[�p��|���u��!���Bp�dL��c�=�H$b[�׫���9����)�N����L�TOOϜG���֪��ض�z饗l�         `e���מ={l����*�0f]����uj< �̹)���@���{ ���;�%�o�>�?޶��ahݺus�ZW(��7 {��q�y������/���.^�hk          +O*���?�d2i[���j���κ�H$��+�ܕ�d��f���n�z'	N����X���z���m�Q^^����Yׯ����۠RRR���j��f�Y���?��>          �套^R__�m��ZZZf]�>%;�����}�Ѩ���g]���Ӛ5kl���ѡ���7�� ��!�`љ�����'��D���������;��F �G��	���"��i[ߡ�!���˶�         �����i߾}��hjj�s���ؘb�����kxxX�Db����:����^��Ȉ�= `>�,�7�|S�|�=�����zg]�����XR�Ԝ'1��n566���W���zzzl�         `�3MS�?����m=�n������T`0Ms� �Pss�ð�w2��O~��X�,*�߯�{���#??_MMM���R)���♘�P4�u���I������d2���~�1~          ���W_�ŋm�n�:9�#`}}}�R�"�jbbb����r�������?֡C�l� s!�`Q����3�j����9�����#�
�0�����R��t�>Ž��C��         ��k||\�=���=<�jjjf]�oX��kxxX�Tj��5k��:�]�v��-��gk ���X4����u��q[{��竡�a����I��a[{X|�x\������=�]���ݫ��1[{          X��q��q[{�[�nV���큕)�ɨ������UTT��{jjJO?���= ��"�`Q,�7:r�\W\�d2��+�������К5kl�H$�_���          ��Ç�̙3��(,,Tuu�������d2���4B������k׮�}��{�g�`S �S�,�={������#??_�����)�N����1Ms�]�smx���ӧ������         ���F��3���g�@k(R(��7��344$�4��VTT���*�{?�䓳�]�������z�-��466*??��k�XL>���� �V$Q0��aZ�v��y��R)��          �}�?���!s��;+�j�����l�`�%�I���ͺ�f�9��A'''�o�>[{ �4� l���O�~��|��g�Z�2͵K�����)�cccz��Wm�          ����_���\��'&&��m�`鍎�����zUYYi{�}��i||��> @����?��g��ާ��VyyyW\�D"�����&&&��f�l���K/�����         @�ڽ{�� �n��k&���Ȉ�}�l6;�����6�X-�Lj�޽��  ��; ��i������}�N���ijxx��� r��Ȉ��������t:m���y�         V�S�N���Ӷ�ijj�`�=X ���~E��+����������G��'�|b{ �w �y��W%d^UU%��sŵ��q%	�{�-�Lf��;yyy�������Ç���a{          �%��,� ��~������l� �κ��Դ(��z�)���(� �N��"��_�����5�=��jll��� r��盵��������i�         �BP��}����p\��g��*555�@ pŵ��
�޻��[����Ջ�; [<�쳚�����\G댍�)�N��@n2MS###W\�x<�������K���{���         @n��z�l��p8f����R(��7��5::zſ��(C %i�޽������C���FFFt��!���1kz{&�������@ 0k�{cc��~��g��d�         ����+�(��ާ��Z.��k��ö���b���~��jjjf�~a�߯�������D�����E	wz<UTT\qmll�`) ��9�/sJJJ��zm�=<<�w�y��>          �V �믿�(��� �h4�p8�(�䶑���9��N�S��Ջ��׿���l���p`���a��ҫ��V�a��;����@ ����{m�����;���s�hF	�$	$��8B`L�P�8�]qR��A*/���4�]�`[
`��E�F
 #a$!���{�z�g���tO���t��ޟ��=X�*z�����~���l��n(e�?��?��pX�Z      @����o�����q�Сmߙ�L�z�S�/�U������7���� ͣ������S���}_gjj*�?��'O��6P'O�����믏v{�/Μ9���w�}       ����x��GKY��A^������V��@5\<�}��1����F������
���y�����/e�k��&6?�F�8w�\)kձ���nw����ti����?�������      ������Jy�n�������Ń� ����)�e�����׿��R��C��3��?��m'�K�Պ'Nl���ٳ���:}����e��---ŷ���R�      �s�̙����]�ZǏ�����ϝN'���KY��3g�l�|������������\�Z@3(�{�瞋��ۿ-e����8z����(��ٳ��T���R��χ�����_���^�W�Z      @9����,��a)k�x��>�:u��u���t:�����yjj*�?^�ڽ^/���塞4��;�'���/�Lo���������u���m�U��v;s�[ ����R<��#��      쿓'O�_��_�����|>|x��`00!xC����j���_��_���R)k���\��_~9�x�R�j�Z;N^�z���={v�!�뮻�����o�h4*m=      `�|�k_+�����_����ӧK>T���jt:�������R���o~�����Sp��׾���n�������WVV��햲6P]��(Ν;��y~~~�^��Ν;���wKY      �?+++�W�W���u �x<�����l��0�������Q�z@})�Weyy9{���;v�ض���\����2������?LR      ���_��E��/e�������s���x<.em�ږ��b8n~>~�����~�t:��o����zSp��7������n��رc����~�����6P}�^o۞Q�	�^x!~����      ���A��_�ei�]<���ٳ��T[Qq�������������?���F��ԓ�;p�z�^<��#��0�    IDAT�7??����[��ںo�����ÇK[��_�zik      {�;��N,//���ց]kkk���J[���{U[���3g���?^�z@=)�W����v�Է�.�Ⓠ �byyy�)�2��?����/��      �7���?��?/m����8p���g�ہ�u�[���U������PO
��)���jŵ�^��yee%�Ai��p��2O(E���7K[      ��w/��ri�m}�9�J����)�1??_���=�\<��S��ԏ�;pE�����q����֛����n~v:�R[o����caa���{�1�|     ����׿^�z[ �?>��(u}�.~��5�\S��e�@�(�W�G)u�k��f�59�� ���J]��n���뛟��rh������]�z      ��y����?�qi�MOOo �u����-�e�#""����Ǚ3gJ]�wಝ;w.~�����ѣG7�����t2pU���m�_��裏��      �"y�R��]{� 766��햶6P?[�G�������.��@��)����G��x\�zSSSq�ȑ��KKK���Ӆ6	u�ȑh�˻$:u�T����}i�      Wf8�c�=V� ��N'z�^D���:|�p���[�*�gԇ�;pY��q|�;�)u���Ř�����^��N������F����v{�!�2<�裥�      \��<VVVJ]sk��������2e���ܹs��O��&P
��e����gϞ-uM7o�~غ�\{�����}o�`      �����]�z������X__��`P��@=m�G=z4Z�V�뗽����\��/8Z�ֶ��
��^Y^^��(""J��>J�!      p�N�:O=�T�k^s�5�֏ �J�ۍn�1;;[���w�m�<��Pp.���R<����955��������锺>P_��h�u������������      \�Gyds`VY ��dOi�Zq���R��F�W�W��	T��;pɾ��o�h4*u����tD��|����K�C�����/�?��OJ]      xs��(������u'�,���b0��>P_[{We�#"}���զ�\��{��5�^P-//��>Po+++�7Pe�#��      �{��'K·������ɛ��J�׋^�i��N��g�y��u��Rp.��~��x��K_wRp���tJ_���h��ue��w�[��1      �7���~��5�>�Tp��do9x�`LOO��~���.w������M�kNMM���#���VWW#�ʭV�ԵWVV��?�q�k      �o0����ߖ��d `�ߏn�[��@�M�W�Vk��U�������x\��@5)��$E�}vv6���"B��?����n����9�      �x�'6�]�C�E�~���֢(���塚2]�p!�~�����I�xS�=�\��ꫥ�;�y+�"���J_h�N���0"���=���1�J_      ������S��SSSq����Pp�OQ�o�O1 0"�T��;�RLo��͛������)�~���h��iuu5~����.      �]�׋�������� �oҏX\\�V�U��� �J�xS�
����A��2�g&�Nپ���&Y      �������vK_w2Iymm-��q���1�G������T�믬��SO=U��@�(�o�?�i�:u��u��v,,,D��;��&SRܿ���yS      $�j0��M����I������`0�V���#�j�*P-
�������d���队���(���$� 4�`0��`�v;���K_}}=~����.      �^�O<�D��'%��`.��49L39\S��}�{�V�)w���y[XX�V��N�P��Sܟ|��$�      O=�T�z�$k/..FQ����d}�Y&�T�������O�dm�:܁׵��/��b��'P^��%���;      ��j ���|LMM �f2 0���t{.P
���z�'�(�$kO.�܁��.�����q�ԩ$k     @ӥH5�G�������x<�D���Bj �f܁ו����\D(���t:1�6��������     ��z��W��ɓI�^XX��_NT�oEQ���zLOO'+�?�쳱���dm�܁]�F����d�V�sss���c0$� 4���z���'[�+�      �|)�����F��@�666��j%�HEa ��܁]��'?Iv��n�cvv�뷀�u:����IvB��?���=      P������������R����'�L�6�?w`W)oަ��bff&��n�@3u:���d'�{�^<���I�     �&������8������)ʒ��Z��(�d�ySpv����d�8�l��5�o�      �r<��S�����?77g  P�~���8i?buu5�}��d�ySpvX__����g��_XX��p����EQ��P
?�я��      M���0�����1==m  �D��IZp����~�t} _
���<�L�׿���FQIOH�TEt�ݘ��M��^p�      J���O'[�:���>��3�<�t} _
��)o�"^+�oll$� 4W�Ӊ���d�F�����d�     @S���x��瓭? h �B�ۍ���h�Z�2��
�K��!�ɸ�����d��n҂{D�}      ��?�i��d����D��S���t:��������<��@�܁mF�Q<��I3LOOG��O�h�
�ߤ      M�����̌��@2�^/�����N[#5؍�;����?�^/i�������1==�4�O~���I3      @ݥ.UNOO�`0H�h��pEQ$�H�>l�I��&�C��2�H���%����t��_L�      �(���O~�4��̌�@R9t$R6��l���A�Hm29��j%͑��      ��K/�kkkI3����G I�����S�N���R�@~܁mr(��Z��FIs �������+�~      u���8 ��r(�G�'yQp6]�p!�i�V���0i�~�SSSI3<���I�     �:{��gSG�v���$�����N_#}��RG 2�~g���/����H���G��J���W_�     �>y��SG��x��8u��z�^�~DD>�5 
���nަ��b0��4\'���q���KI3      @E�EG���r�GD(�;�ߙ�l�p��j������,n�rؗ     �nN�<�n7u��F�# 7����~�ܹX[[K�H����N�)�9�Y���/     @���n<�� 4\. #��cg��F��K/���v�	e ��h����7      �{�<�SpR�i�eo򐾹d�W^��`�:F��m܁�r)���g?K      j�w�_�e/�eo򐾹d!�p�VK�Hn8F��J#VVVbyy9u      ��\J��p� ��{.�5 
�@D�u��Hm<��     ��v�q����1"" ���^��/FQ�c �Pp""��ɓ�#DDDQ�\4͖�^t�ԩ�      �6N�<�M�� @ ��E�n7.\��:�	w ""Μ9�:¦\�&͖�^���      ������R*�-�~DD^{4���;�\�rJ ��\�g      ������H 9ȥ�����D�ߏ����1""�&��rُܼ     �������;��\�y��@Z
�@�>}:���\r ��y     ��s�̙�6�T*�+�~D���K
�@Vnހ\�-//G��K      jAG`�����!i)�n� v��~�      �FN��rz&	4�h4JaSN=6 -w���E���
.      ������t:�clґ r��^t��٬� �(�Y']� 9Pp     �����������h�ϟOȀ�;.\HaSN�R��rۋ���SG      ��˭4��sI��rۋr۫�4܁X]]Ma��.����mZYYI      *O?`������j w ����.����mZ[[K      *O? ���@
��pEQ���z�۸�R�mr�      W/��n�=��)��(��HC�ncc#F�Q���v�4�x<Na7o      p�r{��VEv{Qn{5���;4\��K��q�      ���s7� ������@
��p+++�#��H-�}(ǽ      �&��d��R�9r�GD�W�Sp��[[[Ka7o@j��C�� z�^�      Pi9�ʱ\
4G�{��;�����`��(�+�G��     ����37	 %� W
��p�n7u�ܼ)��_     @�t:��vȱ\
4G�������(�C����v�H%Ǜ����`�:      T�h4��h�:��>��!�=(�>P.wh�\/r�x�!�6
�      p��# vʱ#�D(�C��zA�H%ǩ���      � ��m�@*��8˂{��5P.wh�\/r-����/�rݯ     �
r}�VE�S���#��)�C��zA��P��?���      P���>�@ �\�EQ�wh�\��^@���Rοp     �����MGH!�'�=(��;4\�EQd}�S��N��5      TA� #�~N	�W�C s޳�r(�C��|1�([��N��5      �.�R9�L��ʹ#���C�.盤�/��z�yO�9      �.��m�@�r�wܡᦧ�SGx]9�\���\��5      ��λ&�#�)�=GG����w9_�~!��x<��(R�x]333�#      @e���MG(S�{NΝ6�
��p9_E��4e�^ܼ     @}���-��@����g�O��	e���߸y     �+��*�}����;4\�I7p@Y��a�o��      \���U(���{��j���T�@b
��p����~A�CQQE�o(��      rV��m:@r�k�����j��$�����x<ξt
T_�7o&�     ��ȽQ��@����G 
��xU� ��# 5W�}�
�p     �\U�y[�[�VE��*����Sp���B�=��*������*��      �����h�Z�c���(b<���XzX
��*�"uؕ�;4܁RGxSU(��5�+q�����:      TV�Պ����1ޔ������T��V'U���L
��p�J�MU��8@uU��-"�����#      @�U�#Q��@5Ua���^�?wh��\(���
7o^�      W�
��hd�.�/���Ta����;4\U.�P@��*o���^      9��s�*<���*{KU�꺨¡�I��*U9AT��7      h��<w3�U�[��WׅN�Rp'K6��������L���*Y@u��.��7      �zUy�쵪��>�:{u]�j�+w�4�SGh����pI�RD���      4KU��U�Y&PU�]Ue����h�J�v��N�\�����é#\��h���g����y     ��W��nU*���қ!��W�AU�34��;YRp/W�.
�t��J���>      ���s7�`�T�Uګ�@��\)����x�:B�\s�5�#\�*R�|EQ�_=z4u      ��*�#��L�W��VUګ�@W�\)���*���믿>u�K6���Z�~T�}      ru�uץ�pY��\�S���V�ǎK�Qt�ȕ�;YRp/WՊ�U;U�J7o�ۧ      Gǎ�����1.Y՞k��Ǖ��]{�133�:F�T��fQp'K
���	e?�ըګ�����      ���v?~<u�KV��pU��� X��x�:�J��,U�xX'N�H�T�d!���ݼ]{�1==�:      �B�ʓU{�	�j{H���:�F��`7
�dI��\Ǐ�v�Z�A�.��|Tm�p�      {�jo��F��Wd8FQ�c\���j��j5Zi����njj*�=�:�e����p8��/ܼ     �ީ��7=�JTq��]uU���
�dɩ��8q"u��R���U��j$       gU,OV�9'�VU�UUܣ�N��\)���*��ZuU,P��.��7      �����>�ҩj���{t�)��+w�SE����1�-oyK��m4�h4J���޼�x㍩#      @mT���.p9�ؑ����cǎ���(��H��l)��%����SG�"~V�KU����jUv     �9r$�9�:�e3�T������n�)�m��2U�KCs��R��K�q������pE��a%/Ȁr�(�"u��v������B�      P+U�H("�����#�;�����~%�44��;�)���E�*;~�x,..��qE��o���DU�      9�j��@��T�m:�����j�Rǀ])����x��0u�Fi�Zq�M7��qE�á���/y���5      �Y�K�U����� #t$R�o
9Sp';EQD�ղy&PՋ����ݸy      ���s��`` ������ᣪ��z�Q!K
�d��nO6OJT勄~��ءʯފ���      ��馛bjj*u�+b �z�< �ȑ#q�ȑ�1���W�WC�)���v��n7u�Ʃ�	e7p�n�|�6;;7�pC�      P;333q�7��q�.6�+ݝ2 0�n������N�Z��	�	���o�V��:�sl5�*�꭛n�)�m�j      ��\�,���þ��W�=��{r�u���F
wdIk�,�Z-�XXX���`S܁��~P��xG�      P[U7"����#"n�������x<Nv��N��ӹ�;RG�*���Mo�F�c\����=�#      @m�~��#\S܁�� �БHar0�wr��N���p�Anު�     @����w���L�W�@`<�p8L�=z4����1���FQ1�CB���RQ
�T}�{��pA����Oo��k�ĉ�c      @m���ĭ�ޚ:�U3�� MoOc����z�vdI��,M^Q��eU����%:�:�U1���7ou8l      ���[���~����1�F�Q-�uu؋�hRp�v��!K
�di�o��I��yZ�V�v�m�c\57p�L�����     `���\����.��W���FDD�����N��ɒ�{Zu�h��2��(��ܼ9�      ��;�V��:�U����\��`��(u��677o��S�h�I7scc���$�%w����#◧�(W]��uypi��~E������;���1      ��:7�pC�{�.���7W����v[LMM���H�n��ꪂ;YRp'K�����z�$���w�3���S��u����x<��������w�y     ����-�uzf
��� ���\E[
���a�v��Ҥ�>y嚝���w7p�u:����/u      h���+u�=S��+���u�����i0�p8�����v��� K
�diuu5"�S��>�:���1{�
��p8��p�:ƞ���SG      �Ƹ��j���'����p0`�:�_XX0�=��������I��)�������x���h�8M3թ���(��v��c�Ç�;���1      �1���n2������~�{߫`����zDD��*���O'Y�p�BD�V\�l����o�cǎ���g��a��1�=���j���|���      UQ�!��{�
�s�g���*�t2��q�$�����p8���鈈X[[K�������������A��F��\���SG      �Ʃ[�r<G��O�Cu�=�H�3�d*��3w�5y���{:u����IFhu    IDAT�n��:j�Z���/u      h�w���q�С�1�T�ߏ�h�:���a� �|��q����1k2��n?Wԋ�;�j�Z��͔�����<hP�� ��a��U��z�;E��w�;>�:      4N�ݎ�����c칺�&��@O����F��t""6�r��N�&�HMpOgaa!n����1�\�ۭ�+{�IF�Q-_���      ҩ�[�#"��q-���$u Q�=�*�^]]M�ޘ�;ٚ�{��W&%��~0u�=W�S�PQu����      ҹ��j��������T�p8��`�:ƞ[XX�;�#u���Zp_ZZJ�ޘ�;���؈��ʌ+++��4�=��S���^ B���d������|g�      �X�\sM��=�Ic_t:o����� �_��_�����1kk����	��Sp'[[7R��H��믏[o�5u�}Qע,��`0�����~���<L      Ur�=����/�\���������U1�b��m��ɚ�;�:����Ӻ��{SG�n�:��q�z��1���7      H��{���1��7�Cu����F�c����x��ߟ:FcE���4E��)���3g�l�Y�=�_��_��d��hT��,�E�ۭ���'N��M      P%�����=�c�o���ս��+��+133�:Fcu�����wș�P�����yJhmm�vBǎ�w��ݩc�~���7��^�Wۓ��"      �P��wEQD�ө�p1���(�������V�������ȝ�;Y�܋������i��{�Ia_u�]�( C�� ��~����      ����pLMM���o��q��PUu�/-..�]wݕ:F����n����$LoN���m�{��!�w�=�D��Jc�8���ǵ~�VD�[��ָ��S�       ~�СC����7u�}5k?h�����~��=�ܳ9�4���w�3��n��j��q)�x�����?��&�{��f�zyy9����%��tǎ��o�=�~���Q������B�(�xM9tr����       \�{�'�|2u�}�����n+�B�r��{�I�ъ��6��̙3�n����(����D�ժ�_ܛ�?����x��j~~�?==���צ�9r$"".\��2q�}�պ��������Q����ڭ��V����R�       .�|$������t�ۍD��Nk2���ڸ��;S�h������_}���?����K�	ވ��v����?w:�m,���G?ڈ��Mx��)��θ��S�       .r���FLnʛ�!WM�;x������T��������������H�ޜ�;Y�zJ�(�m�,囟��{�7u�Rt���F�c@��F�v+"���D�      ��h��L��u:�ڿ�>�7�����c4ޅ6�<==�0	\w�v���m����r�4DD��o�F�����l�E$�b86�'���éc       ��;n�)u�R4�Y-�I�7����ŉ'R�h�����p�0	\w�����w��]q�-���Q�&�Rk�T����133�:      �x���JӤ�mCj�^/�A��i�@՜��X__����ϐ+w������Ғ�q�����J��N'u���(bcc�Q�{��Q      ���Q���V���v��СC���?N��.\����s�̙�i��(������F�Q���$LC�k�����R�(�h4j�di(S���~{c^e      Uv�С���?�:F���n�F��1����a�:H���
�jiii��W^y%Q�t
�d��ٳ�>_��R�4�n04��[Q��tb<��R*��     �:��|���(���F��tR�(�<�:����v�m�;���N�^z�m��n���O}*u�����z�c@m4�"�{�7u      ��y��ַ�5u�RM��5�y.엦������9�F�����yff&��H�.��;�;s�LLOOo~Vp��m����~{��������Sǀ�k�/C>��O���\�      �%j�Z��|&u��5��ܰ���qt:�F�z������[��&�u�&w*ak�}0���j�4L4�"���)��U�t:1S�(���L#�~      Uw�}��5�\�:F銢���%w�B��8666Yn�[���R� v�:�r��N%�z�m�ϟ?�(	[���j�x㍩c$��W���������q����1      ��433���'S�H�$w�2M.�GD|�s��V��:��k�ꫯ&J�G��JXZZ����ٳ���U�Պ|0u�d����4�����     @]��o�V��ͥ��Ĥ��������#G��G?���1���`��˛�[�V<���	��Sp�^z�m�/\��9����J#�^����v��M-�GD|������m�c       W����q�}����LQ�����(u��h4jt�="�������1��o�Y����n��0\:w*��_��������8.\��0sss�O}*u�������u(��桇J      �J���g��nn�j��W�v7����4��>77����:�p�ܹm����I�4���J��;Nu�={6Q.��O������;\�/7^s뭷Ɲwޙ:      p�N�8�ЇR�Hʐ3��p8l�����O|�q�С�1������뉒��Sp�2������ϟO���9r$~��=u���At:��1 �����~���SG       ���>����Sr��t�^355���gR��:�Ύ��W^y%Q�|
�T�ŧ����L�����Ř��M#9�1����x�:Jr7�|s|�#I      �#��v[�}�ݩcd����X	M���u�~��뮻.u~��ٳ�>�Z�x��g��˧�Ne<����>E���N:G��x u�,�F#�^�!��~��h�Z�c       {�K_��瀿����{i�n��^/u�,��������1�����̌7P)
�T�+��333۾;s�L�4��w~�wbnn.u�,L&X�F��Q�4�Wn)����[o�}�C�c       {̳��<+�i���N��� u�l��o�f;v,u~a4����w|U��N����dϝ;g���ѣG㓟�d��(�"666\��N��dj      ԗ�9o�m�4�d��p8L%�����}.u�8w�\���m�]\x��)�S)����>���XZZJ���|�󟏅���1���v��ɩ�~��:JVn������S�       ���7���GR���x<���u�*���h;��M��O:�����1��̙3;�{�$�+��N����+;��m3&�C�ŧ?���1�3�T�v&7nN%������       �/}�K155�:FV&o�7$������?������~���c�EQq�ܹm�MMM����D���(�S)�<�L���l����}.S���h4rR�ژ�p*y�;�#���1      �}v�7Ư�گ����^��NG�ʛ�پ�륎��|0�9�:[�����ym���c*G��J��z133�����D����⢓y��Ie���F��M#K�V+�򕯤�      ��w�wwtYx�p848�J���l�:=�P�\�ԩS;�[]]M����;��[�r�M��z衸�R��V�׋n��d�2�c}}=�A�(����>��v[�      @IN�8>�`�ٚ�=g�j����=��ñ���:9}���^x�I��(�S9���ʎ�N�:�(������򗿜:F�&£�(uxSn�����\|�K_J      (������ѣGS��VQ��v��������(���\�&n����'>�:Y]]�N���v��>�l�Dp�ܩ���~:Z�ֶ�ݮ�hd�#�H��}�K#k��ʽ^/uؕ�K���>�?�:      P����x��S���p8���u� ��h4�������d�_�jLMM���EN�:����i-�$w*��������w{��}�+_�v�V�f�����dǍۥ;v�X|�3�I      H����w��]�cd�(
� �Ҥ�c�ߛ���?l�i�v�P���%HWO�J��"w��G�w�-��<�:F%�F���؈~��:
7y=��K�{��{177�:      �H�Պ?��?�V��:J%L�Ħ���d��C�fzz:���/���.���b}}}���=�\�4p�ܩ�_|q�w���� o�������1*�(���z�����p�� u�ʸ����{�I      H��n���2L�z=��(��Εy衇��oL�]�<yr�wSSS
�T��;�����155��{S��t�ȑ����:F�8J�&S�;��_\�V�����sS      �����W�����cT�i�mr���硫R)G�����c���(v-��Z-8�,w*i8�����O�<�����O�I�z뭩cTN�ߏ��u7q��``j�����-{      �������/~1u���Ǳ���nW��}3�gj����W��c������t:;�?�|�4�7ܩ������z=�r��������w������u:��ɉd� �2Ǐ��~8u       3=��AYWh2��dm���W��`�{ｩc�:v����3ϔ����;�����~�z�5��r�-�����QY�����[O${;�����_8�      �`��)�"z�^����p8L���F���n��UXXX�?��?J��QE�:uj������~U��Ne��g?����ߟ>}ڔ�����n�8q"u�ʚ�ĭ��9Q����N$}�c�}(u       S� ^��x�N��"�����??W��_�r;v,u^����w�j�*U��N��6yx8��ӧ��R���ſ�W�*Z�V�(�f7�k�^��D�U:t�P����~�      @���?��q�7��Qy����n.�7 ��n�->��O���x��w���^(9	�-w*��?���߿��+%'�r�u�]q�}���Q��(666�y]��n��D���W�G�I      ����!�{h��rEwvS��ψ��{czz:��������`gΜ��}�ݎ��~:A"�;
�T��Ø����������$Hĥ����}�=����&?^ն������>�:      Pw�yg����c�����;~&�����x��ޖ:o��ɓ�����v��`�(�Si�� ���w|_E���	q�<�G�:F�(53v�'�������      �e�����8v�X��r�n���Ql�_��rK��o�v����_~y��w��U��N�={v��_o�&�������'RǨ��p��뱱���0uJ0b}}=:��b�>��?�ø��R�       *fqq1�ݿ�w�n�j�(���)97�x<���>�����o��g����Z�����ߞz꩒���s�D���?�u�n�ۍ���'H����?��x�[ޒ:Fm�F��t:����3549�����n���}��<>�я��      T�?�G�(>��Ϧ�Q[[��WO��(�ݮ��%��W�7�|s����^zi��gff�%�����N�---���ܮ���6q�177�'���>����vcmm�E~8�\�믿>�����c       ���ǻ����1jo8���Ft:o�������;���@��o�f����x�����mee��4�?ܩ��;qt�����z%��r�z���/~1u�F���krbٍ\�LnڜF.O�Պ�o�M,,,��      T���T�ɟ�I��ϧ����0:�N���E����ٻ��,�;��~.��2g0�9�1����ƉǁqH��g�v<���Ď�ĎI2US�������nmmm���TmM�&�L��E��/@ �� Y:��=����GVv@�x���y����*������.�ۼ=���c"fM�:U?��d��QpW�^�e�����N�w�����`�m[W�\q ���꯴f��c�n�7m�:p��V�^�t          9�;�ГO>�t��b۶��B����0� ]���1C����5u�T��`���o���~����2�H
��	===*((�鶶�6>�d�0���ϫ����(y���H$�D"����,�R<��a˖-�7���c          �1�w��֭[����L���0@��9/�L*�2��a�<�֯_�t�A0Եk�n��ܑ3nuю�b����pLČ3������A_�i��9#��ڹ�vVII�~�����:         @z��g5c��c��=e��3M�so����%K��;����10F���.I.\�` �(�#g�?�����.�p�-[���Gu:D�=n����{������={��Q          䨲�2���
NG�{�K?۶?�C	�ü��%JKK���/���;c�H$���y�m~���ۀlD�9���S7���קP(��D��'�xB�֭s:np�M7sg�����C�_K��ַ��k�          �ݝwީ�}�{N���8�n��mY��Ѳ�eYJ$�D"
�BWt!�0��/0 0�\�r�=�`0��4@zQpGN���鿷m[���N���x<|xr�/�̍܀p3ws�ir�E6lؠo|�N�          �'v�ء]�v97q�!v�d���M�ڣ����W4���b���wB�El�V[[�-�WUUe0�~ܑS*++e�M�uvv*�Hd8&���T���
��r�_!
������n��v���=���~w�q�:t˟#          ��<�-[�t���@�H$�����C��x^vnUhgHbv�򗿬}��9���ݭH$r�m~�_���N�w�k׮�����L�T{{{�a2��N=���N��8�X��������9Uz�,K�dR�X���n,����k6z饗TRR�t          y����W^є)S���q
��>�V�X,�D"�3���.�H�}��J�={͝;W�?�< �Lkk�-����g0	�^� 7��|�=�S�*��Eyy�
o�-
iѢE�p�"K�,Q�������	�m[�e�4M%�I��q%	%�I��)˲d۶lۖa����1���Z<W,�^ؿ�π�u��A�w�}N�          ������t�R}������,6RO&��;7�GHr]?���#�G�#=�ٯ��P���/4s�L��`�����g��r{EE�b�؄ֶm;
�~5�l@��� �Zee����{ӧ c�����t�w8���3Ϩ��C���NGA������t����x���f�F�������ߏܜ��eY<]�G��ۧ|��          �ܚ5k�������7�� �F� ��1���x�#	J���0:tH.t:
����˷����u�ڵ�2��;rN$����k~ZZZ4g�W=����~��'?��Ç����t�ٍ7P1����b˖-z�'��          ��GyD]]]z뭷���8Q�aЏ��=��ڴi��10N�HD]]]����֖�4@�x� �åK�n�-���/�i�
eee:|���N��t�܍��F�l�2=���<�         �U�~�iJ���={��Gq:&���˷�^�z�����p" 3(�#'�?^����Ғ�0H�9s���^��- ���ٳ��          p%�0��/h���NG�֯_�����w:& �����ۓɤ�D�C�9+�r����3���l�2��?`�2�	+--�          \-�'?��f͚�t Ylɒ%z饗��P�F����,��/\���4@fq�BΪ���}����A*mݺU���w�� �|>���˚7o��Q          `TӦM�믿����� �B�f��O�S�n��L�T{{�-���~���d.�aܑ����F�><<��DH����k���N� �E��~��Y���(  	w�    IDAT        0&,��/�,���t Y���D�����M��tLP[[���-����g0�yܑ����F���ܜ�$H�g�}V۶ms:�,�w�wھ}��1          `\������z�NG�


�ꫯj��NG����˗/�r���ѩS�2��<
��i�O��+W�^e�{�x<:t�6n��t .��O�/��/��          �y�f=��s2��( \����W^ѪU����IhooW<��v۶�3��<
��i�e)
��OSSS�� �^�^~�e�[���( \���ڿ��1          `Rv�ء�RrpS��r�i�jiiu����̄D�9���ӣ~����b�{�y�p���NG�2_��W���;          Rb�Νz��'���e<�:��7:����6��v�߯�>�,�� gPpG����U u�����A���^�ҥK���%|�A=���N�          ��z�Gt���c p	�0���}O۶ms:
&�4M]�|y�}zzz2�pw�K�.����ի
�J�t)**��Ç�h�"�� pؖ-[��s��j>          9���׾}����a�a�g�Ѯ]�������v�׫���&�C�y�ܹs*,,u^ۑ����_���;�Ƕo߮_|Qs          �'�xB_��ל��!�a詧��_��_8)�L&���2�>�Xl�<�K�N n���{<��


R���Y�4ں�pX���***J���Y���ھ}�jkk����t �{�n}��ߧ�          �����O�@@555N��A�G�޽{���ijj��f�N�:�p8���ڶ�B�J�@
��B�8~���~���466f(ҭ��D?��ϵf��� Ȑ�~X����d��Q           c��߯����q:��z�������;w:)�����6�>�G===J8��;�F<W,u���A���f(ҭ��P����֭[�t i��~=��3��         �}����g����9���륗^Ҏ;���jjjR2�u�����܁�;��ɓ'���מ)��@����6o��t i����'�p:          8j�޽:t萼^��Q �AAA�^{�5mڴ��(H�H$����Q���|�x�b��@�y��������\���D���Ǔ�@2CO?��8�t          p���_?��)�9���X?��ϴv�Z�� �eY֨��gD>�\���-�x<O���HDs��u���!-X���ޑ=��ƍ
���� �߯�^�v�r:
          ���d��>}Z�d��8 &���\?��ϵl�2�� �u�ҥQ��z����d�vZ2ض�B�J���$��E޹|��nW���b�|�r�!S<������駟�� �����g?���o��t          p����뗿��f̘�t ��h�"����ŋ����m[�.]�mq�����ށ\�w�J&&��(//u��А�͛'�ϗ�,Ȭ�˗�K_��*++e���q �Ü9s����Z�t��Q          �զN��m۶����t:�qZ�v�>��S�:i��ե���Q��x<:v�XZ;nLp�[1�y���N�����c��>��%B�mڴI����|� �������_�R���w:
          d��ӧ��韴~�z�� ��;w���_Wqq��Q��e������B!���$܇	�p�LNp/**RYY٨�k�̙�Dd޴i�xR��7o֫�������          @V��|ڶm��� ��3C���7��SO��a~q�jiiQww���x<}��GJ$i��w�w�J&�W�^�ڵk�L&G�/
i޼y2#홐yEEEڶm�o���3����������|NG         ��d�֯_�@ ����;�M��~���z�ᇝ��4�F�����mۣ���UWW��<��V��*�,�KRii�m�G�Q�v�;�W ���߯d2����� ����~<xP����!#          H��+Wj�ҥ:{�lڧ�3f���ú��{���4���U0u�0��'�(��=�eY�P(��i?0N���s�'�R���B�������ŋ������z��O�^P�� pkw�q���_�E=���Q           ��_�^��կ�h�"�� �t��w�_��_�l�2�� ����}����]���D����\a&��UF&���t�*eee���n��,��̙33�
NY�h�6oެ����>) =֯_�Çk֬YNG         ��TZZ��zH���jiiq:����������ϫ����8H3۶U]]}۩�a��O?U4�T����������@���D��ʕ+��{d���i���
J�L�2E;v�Е+W����t o�ܸ=��s\k          ͼ^�6mڤ��rUUUɶ�dJQQ�~���k_���p:2���]W�\��~�dR�ϟ�@�?�,+
�(��u(��U|>�b�02Zp���S�������k޼y|��~�_[�nU Ѕ��Ҭ��H/�����կr�         �Z�d�֬Y�����M�ټy��_�B�W�v:
2$���A"�0��'��v�{*ٶ�B�c�N�w���%���Ck׮U2�u�h4���BM�2%C��$�0�r�J�X�B555��ir�]w��?��V�X�t          �K3g�Զm���ܬ���� 9kǎz��WU^^�tdPmm����m�K$�p�B�7۶C��F��*N�%���`L����͟?_^/�>�bΜ9z��u�ʕ1�&��x<�۷O�RYY��q           �iǎ*--����eY�ӑ��Q\\������|>��q�A���jll��~�G}����xR�7˲�C����ѓc@C������H���ի���{o;�ݲ,��q͞=;C��ڶm��̙���j���t$ �͜9S?��O�k�.y<��           ����/_�\�ׯ��a ��뮻����Lw�}��Q�a�i���궝DI
�ê���@��3Ms(��?1p��*Nܥ?��������aM�6M���H7Y�x�6oެ�/j``��8@Vںu�^�u͟?��(          ���>}�v�ڥh4:��� ����Ձ�����f�<��g�������y�^����c*§�eY��p�����۠�W)��0������W��sϘ�sh��L�CS�L�Ν;e���꜎d���"=��s�����@ �t          �(�^���>-_�\555�F�NG���ٳ��k�iǎ����`0�.�i���A555�9�͙�9��WGN���;\�邻$E�Q͙3��%�I%�I͜93��6�Gw�}�V�Z���z�B!�#��v�Z>|X�W�v:
          `������r�:;;����az�����xL4�&˲TUU�X,v�}}>���}Y���d�4��p8��9rr`��*n(�j���c��144���re �h���ڽ{��^�d۶ӑ W)))�w��]=��S*))q:          `����}�v-Y�Duuu�D"NG\g�ܹz饗������9jjjRWWט��r����Ӝ�֒�do$�� �w��H�=���8����G�/SYy``@���w4/���zu��wk�ƍjnnV�ӑ Wذa�>��ﾛ�m         @�7o�v�ܩ��a577;p�׫}��饗^�ܹs����A]�paL�C�ϧ>��ѡ��i�D"��ñ �-Pp������D�dɒ1eH&�2MS3g��@2�ٴi���C���Luuu2M��H�#�O��C�����          �c��6nܨ��[/^T0t:��+V�?���o�.��:f��m[UUU�F�cڿ��V}}}iN5�d2y5����� n�+*\e���������֦U�V���<44���rf ����h���ڶm������� ��ݻw��^��ŋ��          H�Y�fi׮]�z�jhhpt1�i������jڴiNǁK������sL�z<?~<͉n/�wD������Qp�����>2�}�����͛7����p���R=���7o��D����ʕ+��+�hϞ=���N�          d�����w߭6���C===NG��0=��z��Wu�}��0�#�%���Ο??��}��ɓ'
�2�lt�D�-���N� ���;\e����z��������v�s�=J&���7�L*�Hh֬YH�l`�-Z�={����H�.]��% �����g��SO=���r��           0}�t=��CZ�d�]Q�Rm�ҥ�я~�GyDEEENǁ�X��3g�(��i�x<�s�Υ9���b��X,��8��"
�p������sE�ݶm%�I͘1cL��A������4�ɐM|>�V�\�|PCCCjmmu:0iz��G��K/iٲe<�          мy�w�^M�2EDN�>}��|�I=��?�M]�xQ���c�������s��1�5���s:�E��*7Np���NǑ$���i��ղ,kL�h޼y�z����i��ͺ����֦��>�#�a����?Ֆ-[\�0          �=<��/_�|P�HD���NG&$\��b�
������U__?��;;;]5 5�]������9�/��W)�{<��\w��U-Y�dL%w�4�u�wd �Qyy�v�ܩٳg���E�p��H���Z�J/�����߯����           \���H7n�}�ݧ��N���8	�0t�����?���l��A�p�d2���J��9��}>����4��h4z1�H���9�/�"�Jaa������Sii��q>g׮]***��+W��Ә��4M}�����o~���n�� 7�|�r=��cڸq��Q           Y���^����U[[�t��������o[�/v:���s����5��ϟ?�����'۶u�ڵ�
�Ï:��"
�p������UYY��q>���i����F�c����hӦM��s���ɤ>����7������q IҢE�t��mٲ��l          R�ܹs������F�� ׭]�VO<�,Y�td���v��Սy˲��o�1�����`0H��D[�2Rp�x<�2e��q�̪U��t��1�_\\�-[�����1rI"�бc����t:�Ԃ��o}�b;           mΝ;���WSS��Q��֮]����ֲe˜��,2<<���
��9���^��9�H$��d�L&5<<L��Dk�2Rp��iӦ9�����߯d29���ϟ�իW�1rQ4��o��7�x��;2��;������u�V��          ���m[Ǐ��������8��a��{�Ձ�b�
�� �X����
��1��٩���4���D"�P(D��D{�rc�}�ԩ�,X���jϞ=J$c>f�ڵ�3gNS!W%�I}��'������V�� G�\�R���ӆ\y�          ���z����ՙ3gd۶�q��|>���h߾}Z�h��q��jkk���1��=����?�����)�Õh��Un,�O�2E���D7���|E���c����j���*))Ic*�:n�Jܴ          ܨ��Uo����;6����顇�׿�u͘1��8�bW�^UMM͸�9y�zzzҔhr�Ѩ��(w�w�ʍ���R�|>��ځ�FǼii�6m�$�כ�T�---����O>�D�i:Y��6          @6�v��y����[v:�ЬY��w�^�ݻW���N�A���:y��䘏�|��P��D��(�Õ(��Un,�+8���fϞ��[���`<w�\�Y�&���O����������s�S~p�e˖i���ڶm�
��          ��D"}��Gz��w����t��aZ�n�v�ޭ�7���8	9 �L���B�Ph���|>��p� �P(�D"A��D��rc������%̝;w���U�Vi��iJ�|d۶jjjt��QUTT��C2���X_��W�w�^�y�N�          `R�������ѣLu�甗��О={4{�l�� ǜ?^����:���F�/_NS���2M��;\��;\�Ƃ{ p��a��c�=�X,6�c<����/kʔ)iL�|
�t��q���[jmmu:�d��ٳG���


��          @J%	�>}ZG�UMM�l�v:��x�f��޽[�6m���u:rPkk��uL4�ѣGӔ(u�]�&۶)�Õ(��Un,���~���8����Ν�M�6�kjvAA��l٢@ ��d�g�m���V}��***���4�;w��nݪ;vh޼yN�           #��������������u:2`ɒ%ڶm�v�ء�S�:9lppP����,k���|>���J$iL6y�m�ڵk�D��D��rc����d͔�={��{J�iӴa�y<�4��Ĳ,]�xQǏ�����!�#!EfΜ�M�6i�֭Z�b���          ����֦?�P~��������Z�`��nݪ�۷3���t��	���qW[[����4�J˲Fzd��J4��*7��Ț'�<�{�1E��q�p�B�\�2M��?gY�Ο?�cǎ�ԩS�D"NG�8͘1C�7o��          �-ض���?~\Ǐ����ӑ0#��m۶i���N�A�,K�N�� �X,�?��iJ�Z�dR���w��8�ʍwI�:uj֔7��m޼Y�i��իW��H$����ٳgUUU���n�#�&�В%K�n�:�_�^˗/Ϛ�"           N�,K������TUU���۝��[�z�Z�b�֭[��7j�NGB����UGGǸ���|z�7�H$Ҕ*�����D�.EC��ł{YY��^�����Д)S�u���ц4mڴ4�Ʀ��K555:w�Ξ=;�7 u��ʴf��]�V�ׯWyy�ӑ           �	������Vee����G
�p�ԩSu��j�ƍZ�v�JJJ���<��ڪ���qc������֖�T��D��$
�p)
�p�/܋��L4~���7F.�c����y�f�)0>�XL���:{��.\����6ٶ�t������t�R�]�V�֭Ӳe˘�          @�%�I��׫��J���jmm�eYN��i�뮻�n�:�[�N�-r:p]__�Ξ=;�T0Աc�Ҕ*=����D�.E{��ł{aa�
L4~ӦM�C=4�W������_���~���Dt��%��׫��Iuuu<�<	EEEZ�|�V�X��+WjժU|�          �h4������_�
����զM���K�j�ʕZ�r��.]JG�
�TQQ�d29��^�~���g���`0(�4%
�p)
�p�/������L417n�ܹs��Ck�̙Z�n���z�i���Y���jhhPss������Z&�|>-X�@w�y�V�Z�+Vh޼yN�           �a��ZZZ��Р��z566�����X���z�`��u�]Z�r�V�X�9s�8��x<���
E"�q��x��'����/M��gppp���J�h�*_,��|>���:�h����7�Ӹ̟?_�W�NC" ��ɤ:;;��Ԥ��v������Q׮]s:Z�L�>].Ԃ�d�-\�P.��c           rD$Qgg���ڮw$������Q%%%Z�p��~�HW"8˲t���	u��\��3gΤ!Uzٶ}㟗�;\��;\�w�04u�TM\ У�>�X,6�cW�X�E��!�y}}}jkkSgg������ӣ��nuwwg�k��O��ٳgk֬Y�={�fϞ��s��K_��JJJ��           2̶m�����������\7���G�D��RZZ���Ĝ9s�`�}�K_�ڡ������~�     IDAT�ի�>β,���iH�~�dR���#�H��D���ł�$M�:U���U,X�6Lh����ޫٳg�!��P��M]OO�544���a��뿆��'�}4V~�_eee�M�2���O���2;��          �Xٶ���Auuu]�H���khh��:�d2#�
��QVVv�1ғ(..�H�)jmm�q>�Oo�����hR�_<W8�G
�p��l#gݬ�^ZZ*���P��۱c�����}����}�ݧ���4��O8�����W�HD�iʲ,E"IR,���^AA�|>�ø~�d���������            n�D4<<�k׮)+��4Mٶ}�/����%�i����W �$���������Pҟ��@�zG�����~����v���M��s��M���h��r>w�R����7,�r:¤;vL�=����ceY�����i�&����)�=���y2           䬢�"i֬YNGrZww����Y]n����E ��q: p;�^p����zkB��ɤ*++��Ґ
             ��100����	�駟�0�3r����G���OE"�:uJ^�w���b1�={V�D"�              �}��ê���P������wߕm�iH�Yܑ(���r�b��ڪ���	UYYI�             �q�D":s�̄;xgΜQ$Iq��˅�����z�e��SOҟ^O2�)�ҟJ�UUU2M3ũ              �M�x\gΜQ,������jkkKq*g���a�>
��
�T�~뭷TXX8�c'��              �I"�Pee������7MS)N�\�b"�QpGVȥ�j<ױc����'t|__�Ν;�3S�             H5�4UUU����	��zu����rV.u1��(�#+$�I�#�TOO���L�[���G555��             �˲TUU����	��zu��1%�'swd
��
�xQ���յk�&||WW�jkkS�             ��fY�������?�5.\�0�r�[Y��P]d
��
�za=v�|>߄��r����S�             ��dY�Ν;����	���ק����r�d2�t`�(�#k��wIz�7TXX8�����t�ҥ&              �ض�s�Ω��g�k$�I?~<���#W;��Mܑ5r��H$���*Lx���555�0              ���,���L����z��?�1���%W;��Mܑ5r��:s�|>߄���Ϙ�             �+�e�ܹs����>�OG���x.�ِ{(�#k��ŵ��E���2cRkPr             ��4UUU5���a����
�B)L�.�iʶm�c cF�Yò�����9sF��ÓZ���Euuu9��             �D"�3gΨ��oR�444Lj�{6H&�NG ƅ�;�J>\d��}y<���looWCC%w             @Ή�㪬����������ŋS�ʽL�t:0.ܑU��"�_��_����Z���M.\��             �#��`08�u���u�ԩ�r�|.��B�Y%_.��e�7�PAA������Tuu�,�JQ2              ��Dt��)Oj�4u�ر�r7۶�"�PpGV1M3o&���q9rd�%����9s&o��             rO8֩S��'��a:r�H�t�e�0rwd۶���*Lj����>}Z�x<E�              ȌP(�ӧO+�Mj�׫#G��U1����ܑu��b��ӣ��j�|�I�344�ӧO+��(              �588�S�N�����{�Mz�l�H$�� �wd�|��~��gjhh����:�PH'O����P��             ���ݪ���to�����?V0LQ��oC��(�#���Ŷ��N����x&�m��u��i����(              ���ڪ��jY�5�u<�***��ח�d�#
#7PpGֱm[�d���8{�����eƤ�1MSUUU���HQ2              &϶m}��gjhh��Z�G������LA�쓯]Kd?
��J�:�]�N�8����I��m�V]]����d�v��             01�e���FMMM)Y���N�/_N�Zو�;�wd�|m��￯H$2�uF�t�����k\              ��D"�3gΨ��+%뵴��ҥK)Y+ٶ��Ä��(�#+����SǏ=�x<������TYY���              ���a�8qB�^�0�������)H���}�0�wd%۶yu��#G����>88��'O*�d=              n���O�N�R4��Z�a���]���)H���X"�QpG����'G��eY)Y+��ԩS���M�z              �Jkk�Ξ=��>`GG�Ξ=����Kd3
��Z�>㿽�曲m;%k����gϪ��9ek             0²,]�pA)����W��̙3)H��,�J��\�	ܑ�� �o���'�U]]�S\             ����b:}���\�����PGG�N�>���r���(�#�q����~;�_����<yR�P(ek             ����N�8�k׮�d=�0������/�[�lG�Y���{�w�DR�^8֩S���ۛ�5             ����M�O�V<O�z�G/^TMMMJ���m�4M�c �B�Y���ͽ�D"2#%�%	UUU���Q�m�dM             @�3MS555���OY��0�?^)Y/�$	z~�zܑ�l�f��-���LY�ݶm577���R�X,%k             rW8VEE��^���5=������Ԕ�5s	�J�
��z\�o�>RWW�<��}��ĉ���Oٚ             ��r��U�8qB���)[�������jmmMٚ�&�L:�4
��z�GWQQ�˗/����l�x<�3gΨ��%ek             ��eY���SMM�L�Lٺ^�W�~���\���5sM2��m�N� &��t `�l�V2����_�[���V4ժU�R�t�mۺt�����f��d]             @v
�B���Q0L�^�W�����R�n�a`0rܑ�(�^CC�������S�n�N�8���ޔ�             �:q�D����G����1�K�\A�9����477룏>RaaaJ׍�㪪�Rmm�,�J��              �2MS555i���#G���4����$�=�
��	�e)�L:#+�����7�TAAAJ׵m[������pJ�             �O�>��S]�z5�k���7�|S�h4�k�"#�PpG���<v�pX�������R�v0�ɓ'���"۶S�>             �Y�e�ҥK���LK=�wޑi�)_;WѡD.������y|�ɤ~��ߥ��~㇗H$���             θqj�����n���{�,+���*�4�z!�PpGΰ,K�d��YŶm����Ǔ�������?�+W��|m             @�ض���fUTThxx8����K�.���"�k�:#�x� ����-6㩉o��~
凶�6�|>͞=;�Oqٶ���]�vMӧO���K��             ��VUU�:;;e�v���x<:u�TZ���p8<��.�įS��,
�p���-�RAA��Ha����ӣ��A-^�X�i�|�H$���y�^M�:5��             R˶m]�|Y555�F�i9���ѻﾫ�������ɤb��D��W�8 H%۶�L&�����^��?��*((H���i���A����D"i9             `򆆆t��I]�tI�e���dRo���B�PZ���x��@�QpG��b=9�`P���o�2�}D��?���ִ��             01�i��ŋ���P0L�9�P��y���N�m�J$N� R��t �F>�o�aOMf۶UPP �0R�*�ض���F������4-%t۶��ק��������0��              �]oo�Ξ=��������񨾾^���i;G�H&��
|1�H�:Uy�T��WIE�]��^��^�zOV{{�b��,X�����x\���
�Ú>}:��              ������t�ҥ�NT�z������ё�s�h4*˲&�w���� @:��q�c䄖�j׮]��bi9�m����T�V�X�9s��<             ��f۶�����ؘ�b���i�o��v�ϓ/l��k��Ũd�J�&�[��@  �0R�
�hT���;��x�v�4��ե�������� m�            �|644���juttLv
���P�>�����'���q%��.�w�w�J�
�#�~���{�m���Q���*//O��h4���E�QM�6M^/�*             H�X,���z544(���\^�W���:�|Zϓ���l۞�2��J>� �H$TTT�t��SUU���Nm߾=�nl�VGG�zzz�l�2͟??m�            �\gY�Z[[���$�4�~>�0t��Q�B���+�$�I��#�N nTXX����|���JJJ��&>�O_���2�C���Lw�u����3r>         ���[�\�y��{�nv�����V;�}��r\e�ʩا��{�@Rɉ]�˻�$�m���4�ݫ{��@�yB��y��\W%r���!��� �U�R��7o�;�eY��Ew�ލ����8��<�|>�����y>���a��a���h�rQ��0_s2����']���o�gΜ���z��C�������q�޽�����        �3ܻw/�x�x����i�#��p���o㷿�푿�i�R:�.�u�������ܻ���dE��
�������?�.��֔eW�^��rgϞ���/c         Z,��[o�ŋ��j{����������?<��;������������^Y__��`0��!�f����K��� ���1666��ce��a�?>^~������         }U�u���K�.E�u����n݊_��W�֎�f{{{�y������?֋�aq��^9��m���ښ+�G,���^���W�r,��SJq��ݸz�jE;;;�:        �N�4�?�!~���Ɲ;w�-4��_�2.^�x,�w�5M���0_�wzI	J�������͘L&���|��������}/\��Ν�        +�뺸|�r�������}����l?��O��*��f�����;��;�r�#�_����i��ŋ���_���n���[�n����#"b{{[�        �����ڵk�?��?q���ck�""��a������k�ۥx�w�eY�˺�N/)?镣��q?v=�qܶ����?��>�o}}=����Źs�b0��        ��m�ʕ+��?�1��:����*~�dy��n�X�b�8�u��^��+G�O&����<���1����]�;w.��9����؈�_~Y�        �Hm���˗��������x뭷��ŋ���ܿ޾��{������^9���(���ى��}.�����(K�q�!�_|1��/�"F�Q�         ����t�R\�|9�β�����O��2��s���|>?����KJ_z�(�?�~���������׾��l_p�F�8w�\���˱���e        ��)�2.]�W�^��m�l���oĻﾛ�����������;�$p�W�:pwŽ?Μ9?�я�뺣�ؔ�2�ܹs��K/���V�         �vww�ҥK��d�""f�Y����{4M�m�5M����^^�N/�|镣�#"677c2��[���oķ����_�/})^~��x��g=         �[�n��˗����Yw�����׮]˺��o6�E]�G��wzI�I�G�>bgg�(߂'4�?�a���d�8�}���q�����W���0�        `u5M7n܈?��1�ϳn)�"nܸ�����^��㺮���ݣ|�;�$p�W�#p����ڊ�x|�o�z����?�ATU�{J�F�8w�\��⋱���{        �"����ʕ+��D�4��D�u�ӟ�4f�Y�)|�_o���Swz���p���G�6|N���w���#"vvv��_�^x!�A�9        �	�u]ܺu+�^��o��='"�}��7�w��=���.���������^��+��GD�9s&F��q���d2��������.������ܹs�կ~5677s�        zn:��իW����G}�����u�V���M�ş+�2���Q����^��+���F�8s��q�_�������~Ћ���WE�={6Ν;�?��%        �M������ڵk����{���u?���b:���#��bww����G��)�;�r��{D���v���z;��o~�������D������ǹs�⩧��=        � ��oߎ�ׯ�͛7{w}0�o~�r�J�)<��b���8�J�N/	������qlmm��q��o�6^z��|\σ����瞋�>���/�        ��tׯ_��ׯ��xg��������_?�k��c��!p�����q����D��8~�����V�m�{�Cmmm�/�_��Wbcc#�        ���f��~�z|��Q�e�95�ƍ��_��w��y�c��!p����J�����k{{;����>F�Q��.��ى�{.�{�9�       �	���7oތ�7o�t:�=�SE��,~�����<�v���#�����^��G��~�=������?���u�q�̙��}{{;�        �S����͛7�ƍ1��s��L��2~���:��ю�z{������+�wW�W�/������m�އ����O�3�<�>���,         ����Ν;��ƍ7N���(�i���/~w���=�/ ����;=%p�Wr��/k�F�o�!{饗�o��o���GD�Ã���g�����ܓ        `�-�����֭[��GE�u�'=��(���կ~�n��=�CP�e��*�����d�Xę3gr��\�t).]�/��b��꫑R�}�޶mܼy3n޼����3�x�        A۶q����裏⣏>����ܓ�HQ�R�_�����R:� �E1	�4M4M#$^!W�\�+W�������W_��msOzleY�իW��ի1��ٳ��3��SO=;;;1rO       ���.�ݻw�܉۷oǽ{�z,��4M��կ⣏>�=�C�X,rO�^Q��ʲ�����38d�/_�˗/�s�=���wc8������E��;w�Ν;q�)����x���K_�R<��S�        ���}oo��J��;wNT+�I�� ��e�򗿌�w����.���=z��= ������`�677c2���;{�l|�{ߋ���u���E;;;���gϞ��g����f�Y        p�RJQ�eܻw�෽��{��A�� ��i�����|�{Gh>����y>��S�7�O#p�W�������9�c�������cgg'��=�P����}{{;���c}}=�,        ��ʲ��t���������[��g8ƍ7�?��?�i��s8b]����n�	wzI�N��!p��>�����1�ꫯ����W�������ގ�����ގ3g����f���        �@�u1��b:��{{{+���F����o���J\���L���2��%�;�җ��(���ى��S䴹p�B|��ߎ�қU܂    IDAT��B�(���؈3g�������1�r�       `�5MeY���ߖeyjڝ����^�k׮��1k�&��i�wzI��R��b��p��{�x��⩧���~�������	�#�R��|������d2������؈�����܌���X__���5�        �H)�X.��X,b�Xt*eY�|>���rO�b0�ݻw���b6��C&eY� �%p�OQUUL&�������;w�_��_�(�����.\���Nœ���������ݻ�犢��d����q���X[[��d��D       �bRJm��ou]�b�8�˲���NUo�(EQ�`0��/��~�;���r��2ڶ�=zK��b�������S�(����z������s�ū�����+}��q���X.���cG��A�>�>����0�A�F�<�����        ���?iSJ�K�u?��h����뺎�i>�����x��a����o~�w�^�9�@J)�E��kwx��+�*Dܼy3��_�%��������o|�Ѷ��)?C�4�4���       �T(�"RJq���x�w�E|�b���|�.|��,c{{;�z$�o��V���[������j<���QUU�i        @&�� n޼�����B7ն����>C۶�\.cmm-�zhww7~�DDĹs��[��Vlmm�&        8��a���������|�{=�z;<�;<��b��$���=��v�Z\�v-���.�7����Fbw        X!�� �E����q��%�2�����:�8��RJQ�elnn��	�R�w�}7�}��(�"�����+����X�        '�p8<����}Q;O$���"�81�𘪪�������p�����ߎ��~;���W^y%��/�2&���        zl�R�ŋE�|!��2ڶ�=N�;<��|��۹gpB���wމw�y'�������׿��8s�L�m�`        Ȩ(��q�޽x뭷�ƍ����mc�\�'�����?h���rO�K)ťK��ҥK�����ַ��矏����        ���.�]�����b>��Ċ)�҃������E������Bvww��?�yD���������+��ٳg��k_�        �!�Ǳ����n\�t)���=�UUU4M�{�8wxB)�(�2���rOaEu]��~����������7�ܹs1�L����       ����X,��������>���=�S`�5���>�������ǹ�p
,�x����^�������p�B�?>677}�        �QUU\�v-�y睘��'q
�e)��3�D���T�e�F�(�"�N��,��7ߌ7�|3"�_x�W�^����H)E۶�W       �����W�\���?�μ�Ӯi�K�����u]�e�����p�-�x�7�7ވ���(��_�r|�k_�g�y&��֢m��.�R        ������`��"nݺ��^ܻwϕlz%�eY�'������b2��h���R��7o�͛7�o?z饗��g�����H)E�4�       ����H)�|>�[�nťK��޽{�<�{��"ڶ�=N4U.|A��<����(��S�S=,z��X__��~�������ٳgcmm-"B�       ���Q�eܽ{7�_�7n܈��2/�'�4M,���3�����u]�e������[,���ƻ�������3��W��xꩧ�̙31��(�h���:       �X��8��^UUL�Ӹ}�vܸq#�޽��5+c��/N������L&1�)�jh��������ǳ�>O?�t��������~��\�       Xq��(����R�uUU�l6�{����۷��ݻ�X,rτc�\.���3`%�q������ގ�(rO�#�X,�ʕ+q�ʕG���d���q�̙��ڊ���X__�����L&1c8�`0��8xZ�(��/��9�] ��4M�;   �G�Fv�)7b�}v]�EJ��a۶QUU,��X,Q�e�����ۋ�lUU�����4��9���W8$]��|>�����S�7���۷o��۷sO V�r����s�    ��d��$�  X9)����g�J� �d�cv         ��7�ϣ��3`��ᐕe�V         ����I�p�p�|�         ���봂pD�p����r�{         p��y��rπ�$p�#R�e4M�{         p���>�����'�         `u4M��"�Xiw8B]�EY��g          _PJ)��y����pĪ����r�          ���|]��+O�Ǡ,�h�6�         �sX,Q�u�p*����b6�EJ)�         �	4M��2�85�pL����|�{         �RJ1����c$p�cT׵��         ����f�u]�p��ᘕeM��         <�b���Aw��]         �_u]�b��=N%�;d�R��l)��S         �t]��,�8��I۶1��s�          �d��-���2�&         ���<ڶ�=N5�;d�X,�i��3         �T+�2��=N=�;��t:���r�         �S���X.��g !p�ޘN��R�=         N��i�,��3�?�COt]��L�         �D��#p��         ����zH�=SUU,��3         `e���m��|��zh�XDUU�g         �J����4M��Cܡ���y�u�{         ���b�σ�C�yB         �r���b�{�w豔R�f�h�6�         8�꺎�,s� >��z.���<RJ��         ���4M����3�� p��mۘN�"w         xB<8Y�pB�m���?`        �1�����!p��i�;         <���4wp	��i�&ʲ�=         z+���,���=xB���'WUUDDlnnf^         ��R���=q;�P.��	UUU����3         �7RJ1�N��p�	���        �}�q{۶�� _��N����,��3          ��l&n� p��\.c�X�         YL��h�&���aE,����g         ��I)��aŌr OUU����y	         ����m��S�C�;����b6��         GF��K�+��k�;         +������Ê�Êڏ�SJ��         ���.f�Yt]�{
pD��\r        `Ut]����vXqwXqM���ޞK�         �Xm���ޞ��p
���v         N*�^�t��)���,"w         N���b6��#�;�"]����^4M�{
         <�r���|�r;�2w8eRJ1�͢���S         �ʲ��,s� 2��)�R��|��"�         8�߷-���S�LF� �,�H)���F�)         �r)���f�4M�)@Fw8��e�m[[[QE�9         �Bm��|>��msO2� ��4M���E�u��         p�4M��T�D������boo�G�         pl����l)��S���RJ1�͢���S         XqeY�|>�#p>f?r�E         G!���4��e�)@�r �����.����(��s         Xm��l6���rOz�w�S5M{{{Ѷm�)         �pu]�t:��$p�뺘N�Q�u�)         �@)�(�2f�Y��r�zN�|��R�f���羸         �u]��,��e�)�	1�= 89����mckk+��         �隦q�xb
U���m���Q�u�)         ��r���t*n����\f�Y�e�         ��b:�FY��� '�(� ��Z.��4Mlnn�p8�=        ������|]���`.�_H۶���u]�        @)�X,1�N���&p�l6��|)��S         8&]��l6��b�{
�"F� ����h�&677c4��        �*���aT��)P�C�u]L��X[[����(�"�$         QJ)��y�u�{
�����X.�Q�ulmm�p8�=        �CP�u�e]���(�;pd>y�        ��)�eYFUU�� +N���R,�h�&677c0�        �p�8Nw�X4M{{{1�Lb}}=���=	        �Gp��A���R,�˃k���0�$         ��v �;p�ڶ��t�;        @�t]eYF]׹� ����b��{]ױ����_�         r��*��y��)�(��.��i�����؈�`�{        ��Ҷm�eM�� p����h�&���cmm-�        ���R��b��2��w�7RJQ�eTU1�%
        �(�u��<RJ�� |�z蝶mc:��x<�����'        ���m�,�h�&�����U�u4M���1�L�(�ܓ         N��R�eUU��Hw�����Z.������8�$        �#�UUEY��� <�;p"t]��,��alll�h�/        �G��*�Et]�{
�cS�'J۶1�Nc2����z�ܓ         z�i�(�2ڶ�=��	܁�����:���         "����bUU��	܁+�t��_t/�"�,        �c%lV��8�RJ�\.���X__��d"t        V��XEw`e���,�X,���kkkBw        `�t]wp4��{���+'���"�˥�        X�v�4�+K�        ���mc�\F]��v`�	܁��`�>�Lbmm-�A�Y         ���WU�{
����FJ�����x���Bw        �w��9��p�܁S'�UU��kkk1��        �'�u]�r���ms��F�	�ju]G]�1cmm-��qE�{        pJ��\.��u]�9 �	�"�mۘ��QEL&�X[[��`�{        ��ڶ������H)��w���b�\FUU1�c2��h�J        ��K)E]�QUU4M�{@/�6b�c����`kkk1�L�(���        ��뺨�:��et]�{@�	�>C�uQ�e,W�       �ǒR��i�����:��C�	���>b��`�{        �]��r����"��{��#p�ڶ��mc�X�h4��d��8���=        8f�l�6��M��5MM�DQ1�c<�h4�       �
K)E]�Q�u4M�Z;�!����,����h�Z        X)�h�� l�>�%�H)�r���r������8�4        �	�������}��x<��d��0���=        ����A��4���	���'c��h��8F�Q���        �����R�� �;@&>�1����p�y        ���R�m{��m�{ !p荦i�i�X,Q��ew��       �p�_io�&���=����PJ)��:�"z0\v��QE�        �m�F۶Q�u4M)�ܓ �w���X.�<b4D�.�       ��Φ��h�6�����rO�		�N�������p8��p��(�á+�        ���ibv�V��`t]w���c��+�w        N���A�޶mt]m�������m����K����`0��`�i!        ����ߺ��=�c"p8Ev�="b4����E��;        G"�t��7-���R�=��� D�4����F�~        <LJ� bO)�Y�.b����T��R�0���AE��~�K�        �e?P�dľ���jN ���\�������?������{D|�۔��Z�b< �(��    ��uݧ~�/ p:���O���o���O�> %�; G���� Ga0x    ���e,��3   �3���          �w           zA�          @/�          ��;           � p          ��           ��          �^�          �w           zA�          @/�          ��;           � p          ��           ��          �^�          �w           zA�          @/�          ��;           � p          ��           ��          �^�          �w           zA�          @/�          ��;           � p          ��           ��          �^�          �w           zA�          @/�          ��;           � p          ��           ��          �^�          �w           zA�          @/�          ��;           � p      �WE�	   �XF�   ����kkk�g    �VY��\.s�   ���;      ��ػ�ظ�;����)QCQTlY�����J��v`�M�C�ė8���=�����[�m�t�@�E��}��)�}�E�u��AV�S%�d�O�-��H���I�(�D�3�}����"����ן3��O    ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�        _V��    IDAT  @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           �0�z    ����zlll��   ��x<n=   �E�  @���       fC��            ��          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p'��z          ����C��k=n&p'�R�V�          {�񭭭}�G���d#p         �&&#�;��P         �~���z�L�N6w         �]���u��#p''�         �w�}W�I:wR�         ����fwR�q��F�          {���t����F�7          ��#b������T��憭7          ��MR����ꪋ%         ��Z�[�������G          ̲R�C�II�N65<         0U�V�;)	���         `�HLJw2Zi=          `�]m= nE�NFWZ          �e��&)	�I���^�          �L�IVw��D         �t�Z���$p'#L         �)��zzMR���'�          ����^�p+w�)��`         L���J�NFo�          0����[�7�������          f�^���Sku�         ��^���$%�;��         �jsee��#�V�s���7Zo          �aoEDm=nE�NF����z         ��z�� x?wR*���z         �������������          fԅ����I��"p         ��&i	��ʅ         `
J)Np'-�;Y	�         �����$-�;Y�p         L��7��NZwR��zw         �ɫ��믵�G�NJ׮]�qD��;          f̥���z��;Y�E��G          ̒R��i�nG�NZ.�          �Uk�g�����\@         &��r����;���         L�x<v 1�	�I�	�          �UJ�g�����J)���          0C���¹�#�vJ�p��`��          �������#�v��d6����z         ���~�p'w�s!         ��R�_�� w"p'�Z�)         ��Z<LzwR��zw         �	p�0] p'5O
         LD=p�����J�p��`5"�Z         ���GZ��;q�;�]���         �q�m= �C�Nz�VT         ���c�	w��         `g��t����j��z         @�	���;���FDm�         �����Z�����޻ﾻ�Z�          �(���w:���R�          �ä3�tş�          �E��;�!p�J)w         ��W���_��UZ�m�W#�@�!          rv8~���.'��7"�/[�          蘗Z��!p�3J)�z         @��/��;�1��G�          ]�����tJi= ��СC�mnn��          ؎����hD��C`���t���ʻq��         ������1w��[�          tA���Zo��%p�Sj�w         �m��z�K:�� wcqq�X����;          ��:��C�n8��NY[[{#"ζ�         �ܷB�N	��R�7[o          Ȭ֪����t�.         ����?i��Ei= ���`0x'"��         ����px���Np���J)/�         �����,�;�Tk�f�          �,�2�;]�ǭ          $�5??�_[��{%p������q��         �LJ)�^YYy���Ww��F��         ��� ;!p�˾�z          @&�}%�VZ�X�#b��         �����G�N8��.[����z         @��� �)�;]��          ��R��� ;UZ��X\\<Vk}-<�         �mW�����z�(�N[[[{#"^j�         ����vf���Ϋ��~�          ��)�	�� ة|��r>�}         ��Z��h4:�[o��r�;�7�.F�˭w          4�_B�Ό�3J)���         �F��z LJi= &aaa�Wz�ޏ��i         `����F�c1l�&�	�̄�ׯ�����         ��J)_q;3D��,���          vS)�w[o�I*���<x���x�ZD̷�         �������C`R���̸v����w          �R��#pg��R~��         ��0������z L��`0��Z         ��R�+kkkg"�����wf�ZD���#          ��k!ng	ܙ9�֯��          0E����zL����3�^����w          L���K�G�4ܙI���n�         `j�_k���� �0�Gą��k�         `�������C`���L��G�7Z�          ��Z�o���&pgf�R��z         ���x���#`��̬���o�R^i�         `B�t}}]�L�3�jDxJ	         �	�֯�� �VZ�iZZZ�kk�ՈXh� Z�q�Flmm��LX)%����z p�������z0a�����qlll��L���\��͵� ����p�+q���&wx̴���w�����_m� Z���x<n=  �$��  Ж�q�M��� `��f���z��.���          v�F����G�n�3�����b�          ����{����;`7��j�_n�         �^�R�Y��[��	���?Dď[�          ���o����z��;{�V)執         p7j�����Mw�����ߊ�k�w          lӹ�p���#`7	��3�\�r���w          l�?����#`7	��S���?����;          ���p�/[���&pgO�F�EĿn�         �vJ)_��Q�����9�~�Eĸ�         ���2??���#��;{���������z         ���Z�r�ʕ+�w@w��Z믷�          p�K)��z�"pgO�F�z         �M~k8^j=Z��g�Z�A�          ?g����G@Kw���h�RD�q�          ?���h�j��Ri= Z:p��'K)�i� v���V�Z������8t�P,--���\�z���i�����V�F�XYY�+W����ֶ������ �0�c<o�����e��n��������8 ����knn.>������Ômmm���f����իWcmmm�������Y�^k�kw�:?����F�����D��Zo�i��zwܗ����h�:u*<�Kˀ�mmmŅ����~����- `�R����`0��<N�>�~��ڊ����ٳg��ŋ��  ����RJ<���q�̙���?,����^����J�={6���m_[��=�9No�p�;8��=�������}�ⓟ�d�9sƛ��̥K�����v\�|�}_�� ����O<O>�d�����2�v�z�x����7�|�׸�n������Cŧ?��X^^��E��lnn�����x��css�)����%�k����o= Z���|u~~�q�� h���^x!>��zZZZ��{,��~\�t閯� �u�ȑ���'N��~�۵����b�9���:~�7n��� ��z����g>��ԧ>V����������#��ŋc}}��^#p`��Z�<�~����'&�����"�Q; �)'O���{.����z
p��8~�x=z4Ο?[[[��� @�<��C�/|!8�z
p���Ї>����t���q 膛�������??�p�E�v-,,ģ�>��N\�z�~O���������������zd p����ظ<??2"�j� v��ӧ㳟��S"�C�������������7��{N�8����cnn��`��ﾸ����ܹs��u�� �?�~ھ}��K_�R=z��"�n���8y�d���뱺��������_[[[���; 5�D���n)�oG�O�y<�@<��s�v蠥��XXX�.��k޼�n9|�p<����v�ÇG�ߏ�^{�g_s? �����������رc�w��'N����G�������'`�=��p8�h=�P4�Olnn^ݷo���[o�i���4���o=�GG�����x�w"BP ]����^�����S�{t�ر�|�r\�z5"܏@W�4p�g��k��Wsssq�����~�V�; 3����VVV�{��I�� Ȥ��kq�� ��O|�1Z� v��g��}���� ܥ�}�c����z���x��g��� t�}��O=�T��9r$N�:�z Lʹ�h�/Z��l��
?�ڵko�R�a� 0-�� >�񏷞L���B<���g  wa߾}���O��L���r<�裭g  w�駟��̈g�y&���Z� ����݈Xo����dmm��q�� ��'�|қ}0C������g  �t�̙ؿ���<��SQJi= ئ��#�<�z0!���q����3 `��3���zd$p�_�Qk���G ���R�w�0c�#�H� �6�>}��`������ѣ�g  �t��)����s6 W#����W�&w���h�o"���; `��9����`��{�,yz������\zF7.�[����0D��uL��%P�6�����kbS_7e;66�Ș�	�c�W8DVH��Kk,aVBBB�R�ЕEG3���=��s�O�ؙլ4םs����׫j��fvw��Tm�ӿ���� �&�I|��~���=��O��  � ��`��~��1�kg ��RJ�W9�w�2p��(�����( 6�m��V;8n���p�m��-6��� �RJ�����_��3 �����jG@���U�m{_D�S� ��S���	�	x�\; ���y�W;8Ozғj'  7�	OxB�F���	�z�5�ڶ�p��3w����_��O�� �㰷�W;8��8/� ��vwwk' '�� ����k' 'ğ���9�@��;+���i*���� p�N�)��o X��vp��a� ��N N��� ��y��;�<���mx2��w�յ[ �VL&�����kg  �V���u��X,j'  7��:�q�P;;;� �f�5���������]����`���j� ��5�b  ����L�ժv p���a3�d���8��];�Šv ���|��R��Y�         X;�p:��Z�X�p�F�ѫ#�v         �6�9����N��M�Ӄ���jw          �!��]1�����nB��GK)o��         ��=M��[;֍�;ܜ2��+"�C         ��:7�r�XG�p����E�kjw          ��R�����wjw�:2p��!�����         @���4Ϳ��������G�C         ��x���(�C`]����4�{#���          z�/�m�������䜿/">P�         ������Q�֝�;ܚ�ŏY�         ��]���!�����m�Έ���;         �j��|>����	��䜿/"�S�         ���l���Վ�Ma��c9_m�         ��|2���Qj���0p�c2�N�/��]�         8���j��kw�&1p�cԶ�G�[kw          '�G۶����i��x���wD�wc        ��z`2�|o��D�p̚�y(���Qj�          �n���`Z;6��;���i~6��kw          ǫ��Wrο\�6��;���i�jw          ��۶���������V��G�õC         �[���p�ʈ(�C`���	Z,*����         �-Yv]������vl:w8am۾!��C�;         ��'�t�|>{���p
���K��         �M{S�4�K���p:�J)���         ܰvww_�vlw8%m�~t0�,"V�[         ��G�Kϟ?�vlw8E���ߧ��F�         ��RJ:�����m��5M�RJo��         \Y)�������������i�3"�];        �W    IDAT x�Rʿk������ܡ���?��         <�7G���"bY;���;T2�������v         ���K���A��f�P�|>{D��v         l����i�_;���;T�s������         �m�R��m���v`���4��Fějw         ��M��@�����d2yyD�J�         �)���s���;��0p��888��R^���         ���r�h4���8��|��;�H۶N)�0".�n        ��ɮ�^r��C��2p��i������[#bQ�         6M)ex�X�z��s�C�f���R�3"J�         � G����rο\;�2w詶m<���jw         ��()�������C��3p�k���G��V�         6�_o��_Ԏ ���z.�����         ���p���Վ �������tD�?�C         `ݓs�����1p����9����s�C         `��9�WED��wX�3g^�T;         ���9�EĲvp��a�L�������n        ��J)�=��-����wX3���`0���         =t�����#���<wXC��쓃������-         �#���/:88��wXS���wRJ�/��_�         z�WF���p����!��g�k�i��"�#���-         P�����?���!��1p�5׶�G"⎈�`�         ��������t���!��3p��s�DJ���[         ത�޾�����tzP�8�!��yh0���         '���yѹs���w� ���w���7D���         '��m۾8"f�C��e���������X�         �[)��r�4"�[��g���s�/�����         �蟶m�ʈX�N��;l��s����j�         ��*��Ü�wEDW�89��������kk�         ��UJyM۶5"J��d���+M�|oD���!         p��Rʫ۶��vp:�a;���_��WEĲv         ܀E)��m۾�vpz�a���yJ�ť�i�         ���]׽�m���.w�2MӼ%�tgD�N�         ������a>��|������9�k�Z���x�v         \�=�i�W;�����b�x`4=����-         ?����9�O��1p�-����k��#�Gj�         ��RJ?�s��s��=\����X��\)���Վ        `�,#��5M�=a���;pQ۶���o��Y�         �¹�`��������xT��M���٥��k�         ����u�sf�������x��t�k���ϋ����        ��I)�������k� �c�|�s��=�s�֔��Qj�         �V)����yYD4�c�~2p��4M�Rʟ��Y�         �ڹ�ҋ��yM�x�w��ڶ}�p8|vD��v         k闻�{N�4��v���uM��_�9?/"�y�         �G)��9�;�����[��`�ܨ6�����+#��        @��J)�m�W��p܁��4�=�"»�         ����m��C��c�ܴ��'�ɳJ)?V�        ��(��>����l��k� ���x\�m�~GJ�1��        @UJ)�޶�+"���/w��4MsO�uό��j�         P�}]�}M۶�W�`���l>��f���R~ "��=         ������s�w���ߨlw��m�WJ)wD��c         89���#��s�'"V�{��a���mq2�|mD��v         ǮD��ڶ}v���j� ���8vӜ�])�?��        �������]�Ԏ6��;pb�����x�U�6w        ���Rz�p8�����l6w�D]�p���w�8">R�        ���)�6M���t���1��3pNE���www����^j�         pM%"^7�L��i��Ԏ���;pjΟ?!�|WJ��`�         >W)�����`������i�`����i��朿*"�/"�{         ���yD|_۶Ϛ��o�l'w��6���V��3K)��v        �6K)��p8�����
��U-�_o���?Dħj�         l��RJ/o�������c ܁>(9���OO)�PD�j        l�eD�n8~e�4��v�%�@o\�p�|�4ߓRzvJ��{         6Q)��RJ_�s�k:�~�v��܁�i��M�����p�        ���+۶�o��y��+1pz+����WF�ߎ��v        ���E���9?�i�{j� \��;�w���ߌ�/���EĪr        ���J)���/�9D��� ���X9���_?]�        ���M)}m۶��9�v��2p��l6�`����xO�        ������s�/h��Wj� �,w`-�&��{#�%���=         5�R�/��4��ܦi�R���2p�Y�9�9���R�K#���A         ���qW۶�l���Qj�
w`tm۾1���R�wG�Gk        ��G���s~z��u��p܁M�h���9?-��ʈ�P�         �c��Rʫsο'���G�a� ��d�l�æi��9�š���         n�o]�Y۶���y� ��`�l���C�g\��j�         ����)�W䜟~qؾ�p�܁mpi���R�����        p�/�9u�4�����A ����*m۾#��ͥ�;"�M��n        �����,�����9�7GD�p�܁�Զ�/��ۮ�^JyMD���        l�YD�n0|U��[ڶ���� j1p��|>�mۻ'�ɗD�]���k7        [�7RJw�F�/�9�5���s� ��F� ����`���6�L�9"�lD|cx#        p�������Oڶ}SD�j�;�cu9矌������]���奔?O�        ��OGĿ���f��Wn&���m?�4�kr�O+�����(��        ��QRJ?_J��9��s�w�\����m�7D�����:�T)��D��        ���K)���G�ů׎X'� 7�mۏF�k"�����>���"�L�2        ��EJ�M����&"��� �Ѡv ���ڶ}G�������"��ʈ��p(       �m���{#�U;;;�7M�Ҝ�Î�qs�;�-:w���qOD���'>��V��7�R�#"T�        8L)�SJ�'������s�&��`�p�~��sqq쾷��%�����R�hD|]��        XW%"ޕR���j����kl*w�2��+"~0"~�	Ox�t]��RʷE�#b\�        ��."~1����r�����A ����L�Ӄ�x��ٳg����R�7E�7F���        5�ֈ�7)��j��klw�S6��>�������oJ)}sD<�j        l�ߌ��D�O���9 �����U۶wD�ݻ��O�/��D��#��U�        `ÔR�)��+��u4�u:��_�	��0p��b��PD��x�v�g��^�R�C���E�^�B        X;G񮈸��{���/FĲr Wa��_��m��d2��.��;��        �َ"�}��{SJ�����Ο?�v 7��`},s�wG�k"b����{#�����J)_�e�B        8}���RJ�u]��m۾+"�~1�\���f�������gΜ����x^D<'"�6">�R        ��SJ���]q_D��mۏԎ���l��i��7]����_�RzVD|MD<��7�       �w���F�{J)���=�����(�� 8A� ��;T?o��wϞ=�����)��L)=����{"bX%       �mu>">(�|p0| "��G ���;�vZ�f�D�"⍗���ٳg��u��J)_�RzZD|iD<-"�8"�Z       Xo]D|���@J�C)�����`0x`�C�ځ �; ��_6|�l��dr{)�#��E���KJ)O���J)_�R�="�t��        T�#⡈���dD|$�����h�u�UJ��|>�xD]�n���JX� ܨ.�����u������/L)ݖR�®랜RzJJ�ɗ�u)�))�q)�lD�G�^D<!���p[<       �I*��}��r�R�ED�F���ҧK)�.�|z0���ן*�<4���u ���; �mѶ�G#����<�IO�=�'l��������m�;�����>�����w�jw  W���<�oF���� ����N3���v pm/zы�("~�vp��㎿s�}������Aw����; �F��.�r�Xg����vp2���O��-o���  �nooo^J����R�p���� ��}���k7 'coo�u& �<��           a�          @O�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �¨v   �V�U�j����N��1b4�h4��ҩ��  �7��2��婟�G�Q���<� `{�R=�w]��(����R��ң�Ǉ���~  ��yJ  =�u],�X,qxx�ժj�`0��x�������a>  �y  �Z.���ɏ��N퍦W3=����  N��;  T�\.�m�h۶���r�|��i������~����N �c�\.#��������l���1�Lb<�  �Q�E4M���'~K��X�V�s��s����ߏ�d�ͧ  pJ� ����׾��zJ)Ѷm�����ۋ3g��x<��  ��:�ǻ�s `��l6��bѫa���V���fѶm�9s&���c0�� ��f�  �l>��l6�����)7�������C|  �R)%��y4M�����d���y ���Z��m��9��S�n�j���t��"Ξ=;;;��  `c� �))�D�4k���r��/��8s�L�F^V  �]�=zk����g�Y,��8{���8  k���(����|��[ۯ����"V�գ���jg ����  NA�u��ۻ���s�.��u]�9s�M5  ��&����yDD�9s&��q�"  �������f��c��r���l��3r#w  8^�  p�6mLsɥQMJ)RJF5  ��&��۶�#w  �m�XD�yc�헬V��9GJ)&���;  �A�   �d���9oܘ�r��<rα\.k�  �cl�y|�Z�N ��qttm�nܸ��K#�M��  �w  8!�n8���;�����ٶm�Rj�  @D<rN],[s�9;� �+]�m�����rm����a�  ��  pB��e,�8::��r⺮{t<  }�\.c>�;� @%�.�ن7bnÛk �4�j  ��Z,�X,n��K)�`0��p)�G��RJt]]��j���?t8::������ى�pxB�  pcn�<>c0��y����y �Mqtt��"V��M�����1?N�����Ȼ���3�|>��h���* `{� �	�4.���ZRJ1�b<�����.��e��ױX,bwwנ ��n�<ޗ��j���r���y ���X,��������`��8F�Q�,�1��ǜ�od�Z����Й  ���;  �����zx�R�����ǽ�_n0���N����r������޶�Z�b�X���N/� ��t���K#�>�Ǉ�a����ݽ�����n�  ��j���S��a����hԯ�ʥ7��F�(����a]w�~��3p �[ӯW  �.=�ރ�K��u�\z��\.c>�_�k;::��je� @]�m�y���(��u����2���) �g\�d�kI)����Z�[/�����b����v�����S, ��cq  ���G�^�`0��d���*�F�8s��5oӹ��  '�뺍=����8s��5o���1  ��K��\ͥ���0n�\J)���b���%n��z  ��� ���V��>��1�L���ISJ���;;;W��K7� @��r������qw  j����������n4�d2�꧘^�5	  pc� ��E)�s~~4��������������  Բ\.�ǝ� ���r�q����Uߨ�n.}2ԕF�]�� �-2p �cv�������1c�Kvvv����ꊣ"  8iW�l�y  j���}ww7��q���s��N�4rw& �[c�  ����`�n��lW���+�� �4l�y|4=�纮�S  �(�|�Y�jo��W{��9  �w  8f���~o��l������Ƙ �Z��<����< @/|��{8���n���1>�kt& �[c�  ����;;;1+֜��R���=��<� ���G8� PەΩ�j<?擕�� ��� �	���W2c<��  ��p �.v����|�Ц�����O� �Ӳ=�$  �����{��M"  ��y  �I)m��t0<�w  ��3p ��R���=� ��� ��m|�i�7� �q1p ����#b+�D  ��h4r ����\:b8��  ��g�  '`�oM��1  ���c��q  ��1l�e�_�  �q��W  pBRJ[C�6� ��y�y ����<��G  �8l��
  8^�  P����  um�yt0D)�v  �57� �1��^���  �Z�E}  ��y��   n�5  3�}  ��Y��  �z�A��jgT�L  �Ɖ  �����  ��,�{  @=΢��}  �[c�          @/� �1s3�#|  ��9��  ����  �5�           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;           �`�          @/�          ��           �;      ��q�  IDAT     �`�          @/�          ��           �;  ����݄X��u �s?�VW�t�AFA%���
(�Bѝ�dT�Y:H�`�Ǥ�(�'c�iLd�va��H�.c��`�L�` &��N�Խ�.�[��tOWw�{�����A�t7��ץ�~�[��        ���          @�          ���;           UPp          �

�           TA� `}�� ������3  o��:�8�&�8 ,�����+*�t�t  fO� `}|�t `.n)�@�RJ��� ̅{m X�~���ȥs ��s6� � w �5�R�J��\|�t  �\�㰚�� �vww�#�J� f/�l& XA
�  k��.���o��L&�͆���� �s�����k�����!  �=w �5q�֭�F��s 3���  vxx�JD�G��l��>U: p>9g�h�z>{xx�{_  +H� `MM"��s 3ukss�J�  ��OK f�7n�C� ���YD�K� f'��> `E)� ����G"�-�����������,� 8��i~/"�K� f#����� X���,������d�'�C  0
�  k�������9��8n����! ������ψ���9�����~�t ��4M����VB��7�{�� �|(� ���үDĭ�9��I)�����+�s  g<�_+�������� �d�^��o)��s �Rz���}�t  �G� `����OED.�x4)��y���mo�%��s�}=��31)�xd�������! �G��������9�Gv��'www�K `~� �����'sοV:�H��4�O?��m�  ��988�TJ���s ���9�RJ�%���O���yOD|�t����wpp��9  �/w �5������|�������ǯ^����A ����ۻ�8,���'n� \������z���/����$������?. ��Sp XS)���������F��8B�r�=�����Y �����>����ҷJg�7o�|��g����A �ٸz��˛���J)�E�,���9�����K��  ��t   �{��ߑs�`D�;̈v||mۖ�Q���V���|5"~��͛tttԕ ��/����~���sa�0��)��̼�R����ݏ���q VP�9]�~��9�"�{K�Yvm���:�� 666J�X9"����={��՗K� `q�n p�����4Ms?��y��B�)���RJ�nܸ�;GGG�K� ���_|W���q:�J�YV��S�������oll��3�<�F�0 ������!"~>"~�t�e��~J���ވ��L)}hoo�s��  �xN� x���;���)�w朿/"�Dķ��u�E]L��T�B�k��"/8+)�o圿�s�jD|�������� �q���o�9?�s~gD|D\�9_I��Vn"�yA�������E^pVRJ���F��O����v������9�PD<���[�c=��\���O(��D�y��"��8���JJ�3����y�o� @A��  x(׮]�tD<���)Ԝ*P������/.�  ���^zi�����"�i?U`j�㋼   v�ڵE�᢮��~j����+{{{߳� ��5�           @��;           �Pp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�  f,�T:B|  �`=�s  �s�)�  \��;  �X��SJ� (�<n ���)�  \��  f��P��  �R̢>  �i�F�;��  pQ�*  `�\G��  XS�q�8  e��}  pQ
�  0c�~�7����  XS�qw  �Z���u�� `���  �d4��PL�ߏ^�W:  kl��q�" (i8��C��#  ��[�;
  �����H)��Q���f�  �9�8  ��RZۇN{���  0
�  0MӬe����;� �8�8  �5��r���K�JG  ���~w  � ��(z�^����}��9�I  XW�9�<n ���қ��u0�85� ��(� ��M�SJ���)�ckkk�
D  ��<  e��y�R�4o*���}  ̋�;  �؝�Yz��Zl��F1��~n;  ��� �������K�.�m5_U)�x���TjwF  ��  3v���p8����Bi�occ#�����k� (e����h��y��R  ,ʽΆ���W��>-���6%g�  p1
�  0c�:��o��
.]�tύ�� (e�����
�  ��Rz�<�R�����{�P�׋˗/G����� �b� `��wp=�ʕ+�<�^6M��c�=�����}��  ��u�=���`p��ɲy�<�S  J������V���ă���0._������� `� `ڶ��7M�/_�����=��Fq�ʕ�����  `Q�W�nX4� ���m{ߙ|8ƕ+Wbccc��f�i����yۢ���?   ��� �
�m{��-S��(666����q���(�lll�����~]� (�뺕��SJ1��  ,���ɛ�������܌���x�7����z�����{X��:oT �Pp �9�9�d2�~��#wJ)677c4�x<����899���{0�p8��pM��@�	 @��{�C��4�?�D3e ���#NK����q�ҥ�y|</(�5Msv>~�7(�M�  fC�  �dz���"�t�p8<�s��$ڶ=;_āxJ)���^��~�\��f[$  ��L&�4ͅ��E�SJ����i�8  K�<K`�����h����ϵm��3�yK)���aL�  .N�  �h2��{��T��{��L��   �0� @9ӇN��vЩ�R����K�� ��8�]  �к�[�C�u�: X.�2����	 �rI)�x<^�1۶]Ȧy  X
�  0gmۮt�$���t  ��U�Ǖ� ��d2Y���x<��mK�  ����  �����m�� �ު��]��x<^�  �/�'''+��}��eվ.  �A�t   X�W����H)��sa���V  �F۶�u]���h�����s��m��  ,��x�~?z�^�(6-�{�  �C�  ��899Y�C���V���  ��i	e���iY  ��d29{�t����� ��Qp ����{���kl� `ULK5�^oi����r �2�.�����0�O���  �|)� @!ӂʴ��4M�k��!۶�2  <�i1%�d ��U�%�g��◮��  H�  
��#"RJ�R:;�O)E�y!l���Ӄ���k��  ��t���w�j�s��g�;��i�>�l `-ܹ�γ�鏈���wne�s[;  P��;  TdZbqp  �5}��m��Q  `m9  ""�           �A�          �*(�          Pw           ���          @�          ���;           UPp          �

�           TA�          �*������r�=    IEND�B`�PK
     �9s[���7�  �  /   images/06c5fde6-b2c8-47bb-9830-971f0c5559bd.png�PNG

   IHDR   d   �   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��	�TE�ǳ�����j�kT�@�E�{V�p�@gE'tXdǝ	c���G�qu��X� D��tO��S��ꦻ��%�yT����z�/��DF]�^����}�e旙U�C���/����3]�t1�;t谽����G��;v�f���f����{��a�����o�5?�������޽{�nlll�^��k׮5��KBD���ݻwG؝E����������ܹs��4��������7\'�5	z�u��#$-�8q�-��w�����jH-!���BjkkS�a+�,y���`y���-d�Tޟ�g�z��F4Aj�~hR������������r!���_~'	Z��o�1>�BT+�����"�?I�7���^'��׈6�k�u�^�� I�H���D3�2{4�+��5�零xC6{چ=!�~$�!hN
�f	�k�|4 h1U6��;�����%'�=C�?J�M>d<A��p�V�*Dy�W�S�|l@�9LB6�a�U�H�bh?�r���.y�I�uuuF̚�.I�僆��4F�2I��a�;"�8&G������
��F!g�\�_R7y�?�O�mD"��[����a��h�4���{���H&!r:H��g��6�S�NZ�$��D�v��!�!m�tEX�v���BF:r���4H���lj�:�$�$M��n�t���a2\��@�T�C�u�����A���Yi�SB��yx/^'���@K���P�L�)�)��E[��ۆmY�n���8%�vS��ѻ{^�V2�ۏ�����n�s����N		z�]�1�cv:_�Ӏ�Wg��o?�<'ezT���;v8-�3Bz��m\_-��(��$�0��I?D��O��}u��d��y�]B�.ym�������9�CL�|��&JWpFB�ZX-f���`aex(<�<
!HG*��ђ_�|f��<h7y��Vb�t��F�v����].��҈��������K;���=-g��K^{�e���L��B�ܷ/�(������,�0I��'Bcz7n��	1GK��R�NMV�����F!\��=nv9��I=���D�@�euJ�������2%�D'���f�m�,��]�B�%�L�؇ zH�� !@J�ZB��DL�H�'
G�$Ưt�б�B�����f�;)���zU7�:T���F0��$�!4�0��BST3�W�,:M�'�9y-�3D�^�PtnDI�&���s����� $
s��:y���������xG�N\��h���w%FS @�	�Y�W����o<�KB�?k�#v?� ��du��IH��GxG�B��6�ꕵf��׆g(+<eVxK�dՔ0Ajz�UU-�Q��y�=}�ׄ�6e��~x1���NB%CH��jwJ%IȾ/���4{bּ ���#���Ю�C�h�2!��L�g(�\��@�p�ۜ��;�&+���\�uloI�FP\��vF��MMM��,^آ������|�3B�ٽ{�UUU;�k�����ټy��jtg�����|%�U�ׄ��T�oz�yyW{h9#$^�L:-)�z�27nt��3B�	�����s��;�v��MTt�3)oݚ5k�H�����]��߉]�$���%E#'��N����ӝ�5���G��\��!m	Q��X��^r�KrU�SB4�6}�W���.�I��<c���&�q�"B���R�Sa��f�2%]Ir&d��٦o߾�$LO�k+�y�s뭷6����?���6oٲ�i���f���9�+l���7�ׯ7�F��鿭���i�&[h29�3:|���U�)�RN���h1bD��/��B����
/5p�
��˨�%�\R3}����V�ʵ`��uuu�_x�F��nz���Y�z5���猄<�䓦��V@0ܭ[�D;.�ϛ;w�`y��L�d��K�R[*
�-[��z]�"�ef����=�0)�Kz�&L�/��1Om�v��~)��BMM�k׮]�i~�7�,.����?F2s�LK�}�ĉ�{�����߅�>hH[L��q��Gx�@zu�/M�T�@c�6n�xh[�=
�=V����[�N��'!�r�!��{�5�&Mj�HB`�1lذ���k�u��S�uq�n	��Ս��LWKA���q�2*��xg�g��\֔ /���ţ|��/��#����.����ÇOX�`A�СC#�ӂ1G�!�裏h��,5d<jMc��ߚ��%K���[�Z��N<�D�Z���n:���-��r�>q���}�/_n�~�m�b�
��2^w�GXو��fY�s�k���U��Ih��1�����~-�UF7E�c7l��3�@��/6Ҹن)lw�m��K/��#G��ڣA��/\kU��@G��e��Q[���uB� �̙c+lx�����l�:�(K�\�/�����u6�e:Zۧ�v�y��go�hh������[��3#�3f̰�q�tO�8^��rԅ����������y�S;�ͬY���?��?�����L�bd�*��.�`����[ܳ!���ꫯ~_��dm+}�Qk���=���w�q����י�+��A��^�{�:%0�$�	d����|2Ɇ
;m�4s�7��b>O}�W�l۶����� D."��fu@[�ړ(�JϜ�Q���GE[���m;�;�ͼy󬙢�h�ZL�W_}e=,�M�T��DƭxR���M��5B ���w�O_}�zȃg�YsZ�Fv�azS��2� $p+�������zs5�:x�\G�ò	���(yf�7����6;
�\��`6U6�uxuS�>}�쵾>B,*������E������]����gg�tөN�,��j�m�J���3�zZ���aZ{�z�h;z���>��Z?l�03d����d�ƃk��^xᅦgϞ�v	Z��cǎ5�V�2/��r*~�q��۱4��[+�eX��[n1+W����������r`������=�P�׿��|��שq��H�7�$��C������ok{�1�ӏ�J� -��?�����)�i�J�ѣG�3�<ӎ�Ц`7<�@۸��`{�LK�����`E���=���'h"�Cu�����R&K'��3td�6OJMV[d����6�e�D�Ԕ�x�2!��L�g(�ʄx���_QF�����T����!:6%���eB���&��H)B4r"��?\�<bQ�3�5�Ў^:t�m�(6��%���tB�x����PSFQ!��Ky���9��[�>��Rj{��(X�ǹ�{�:���1!�ZȺ�ey�2!��L�g(�ʄx�2!��L�g(�\��kJ	�b{�2��L�g(�ʄx�2!��L�gp��)#;��C�����B�t�^���:�R +�X[�[�N	ٰaCN}��/�����ņ3B0U.7����^���	;���ڦ;ӕ�
���/�]X�
g��G6�d���p�3�D�h�n���4��ڲeK�}A|Z��KT&W��:���J��2�\u��R\N�[�����CJ��:qF^J).�qyn�3Bx0z���)��2��+T=���M��g�4������(��?_
�PVʜm'��,u7^��>���Ν;���e��{K1��X
�;e���n�-m�Y4�H�s�8<�BU!B��xckjjz��b�9��m�֮]k|?���-�)s�6ekBz�v̓ק���A�+�ZP�bO�W���\��YЈ����F�EDOIWi.���QP��6������!g�c��pS�8��&Cf`͚5N��|�y����[Rf���:������Gm�m�Gy�-�k8%���Ɇ��-2�֭�NK�ڍc�=֖���Υ�w���=o�{�9�tV���I�)��ѫԼ�Ç�/��Ҟ��ː
���T�$�$b/�ux0l9��b&1i�t\O?�t[�vq�B{��92��ݤ:����gR&ʖ����UK�	�1���ϧΈr	�`�6Ƞ,�)ɭ���ќu�Y����ve�Sc�t� Q����O��D �~��Z�)�i,ֈ���M�q�)����уC'h���0��Y�A�3�Cw��3������썞���!@V�aj�;�c�z�-녅�.lT#��ob���o�kxC�3q;�b�M��O�11]�3u3uܔ �����c���	�q��7�"�0���ќ�!����ᑩ��g���=$p��Adl��p:�ʂFO����\�1�#���$l�r�5z$������«΋����E�8U�3���x%�~0I����gA��b�{BQ�}Ј�8a=��a	Q�E��P�J),5a���T�R��M�6m�t���~�J��}2_�~}����D�ϊ��DڽJkn� ��ܾ}�6!����h@[��� ��l�;�|u�ȼJP%�ʟ���bs+�U��ư��V�"pѭ�E�Dً3rOլY��u�ر]ĥ��RkC�����dM�9s���������7��(��S�L�
 �Fu�.]f>�F���-Z�0p���6n��K.*Wx@�[-��U�/�G[��D�녭�%e��b�v {<]�TU7�t����r�ȜQ��e��ʄx�2!��L�gȋz�|g��+h��!L�#�����L���I/Y��N,����U��N?qw�	3��W�Xag3��bb���|��s"�W�Zef̘a>��3;����L�25z�E٘��F
�Y�`�yꩧl�����42q�]v���eme���.w�y�]�ꧫi)�����}��g���jsꩧ��T�uP�͛g|�A[�eÀ��k� �L�bC�ZӔV	A�M�fV�^�"x-<�	�<�9�#�w	�N�ϬdD��\��L�>�\w�u��7+!h��Y�;5$�}��7��ѣ�ݗ���?��
f�ìA�H��V	Y�t�m3��hd����Q�F�}X �5W
���_X'([[I���۶m˹���ځ�Ϛ!z׷}�NW�h�Í�k��mG%�0�R�¯��<+ȶ)߫Fp��/�q����	�!iʆƋ+{7×&X�Äe�{Pی�C������p�� �th��O�����͛Y`���#��	�%>����0x��h7�c�s�9v���q�GJ�xXx�l�t�I�/B�?��ͬY���p��ցk��,�`�;��t	��2�p��H�|¦�R:�G����K/�����!�LUSԼ��^{�V��!TD��I�&�����6̕��(�p�*�4n�8+K<��?��,^���zއѢQgH����k6R\�o���SgA�kfdN�W^y��lhG=u�����2������?l�	w���A��M4��Ȗm� 1-�O�ss��1cƌ��q�k����1>��S�}*�����@c��X�@�_��׶���L�X���OE瓐)�G4�)�-��� �Q�_|�zVg�}�e�c�D�
m�v���q�gG�R�1@͹�1�
օ��rQ\[�Ǡ�p�ٳg�a��0 r3���r���*�C��b\+LTT%�4Y$���=C'�0L�I�$�ݩ}��c�)Ǭ�a��DZ�Hh��Bƞ:��gn���o���{/���P�[�����7d[}�ׯ����󪉋Bֱ,'���RW��^(�>'t�U�C2͆V��u���a������h�� '�����eCN3��bl���-+�-3�]@Wqq/d��!9�A���5�>�Z���"��1W��u'�4W�r���U��r���4@=\��PyRH<P����%��	���U$]��Q�&�4.�%IJ�����	Ɉ�h/BB�qֲUT��5B��g&Ym�(6"e�!���-��{��5Z��Њσ��w�~�4�������m͑!�LD�Q���5���.4�L��I'�.��"		�VIO������YT'KC0	9m��\@� ڜ>Y��<��6H�-C3������?��+�t�I��?�V�o��C6�<#�I�����䖉�B7���^f;}������X�AQπf� k�4�S��~lAn�n�'���]we>9�ʡ���8��u4��B�P��iD������_���r�3��@��U�hO�Cҁ��M.w*�K��3Iw���(yMᆼ-g�͔4Vҹ��y�G�u���py��;����F^W�6xq�_�E��������O�R��fE��$e�+�g���S�@Ü�� ��=�	��m���f3�!�N!b6I�$j_�%D�駟n��ϞU�߇��|�I'M9r��'O�[Xs��m~����)��C�+�������1a��x衇��ў e}8����gϞ_M�8���o�}�8{��#���F&r��ickj��l�����=w�-����"v��h��6�.�'EЍ��р�RF�hl�ܖ<��޽{*��vDOo�YP�p�	MD%�G�CD9���ܐp����ۨ�afTE ��7�l~��_�|��&d`�R�!�<�͕��xsm+��
�_�q�ʕ��??��c&.kp�z���]CS�$!��ޟUD�I�O�{�f��ԕ�h;6��*I�$u��օ���a��EfO�;V��_H-�n�֭�������C�m���+�ib���9yG�|_/ߍ�ڌ�
]�5G� !�"�g��}��Lɣ!�<Z�X�4X'�ޫ�8ks<'�Q�e��QP�G��M�NA��͊��믿޾�q��UJu�_C����UƙGx1mCpR ��<2��T��+���� %ޕ8ƽ�4�s�u<�1��Q ��    IEND�B`�PK
     �9s[�;� � /   images/31959ea2-aec5-42cb-a646-ec7cb3b6e41e.png�PNG

   IHDR  �  J   yp66   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���|ս����ٕd�w\ c���!���)��dUK)���8��I��.K�!=7�RoB
$�$�$�1�m���Μ��Jbp��ڝ����~��n�hV����j�9��r��Z                 ��                 "��;                 (�賄R2&Q(q�-�!�t:�}�>{�Sv��P��*G�&K\�}x�><�f/&�d|�o3��){�k���X���=�C�ً�>��{]���
e�db�J̜3D���n��2�o|��=هg�9���9�9͑�q�s�>4;͜�ҜcMH�8{�{�^�      �@G�@��pdΨYW?i{Qm_ʾ��=����]�B��0'/����d�g��Ϸ�$��z(��$c��/L����}���u������ε��{�����d�����dR�N�����5���WC�w���:���xE��J(�NH������ÐTN����w��*���q�o���C�!eo/�s��|M~�������Y�đ�{���      �`(�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�                "��;                 (�"G)5h��+-c���y�24��8D\�Jaޠ��}{�C<ߓ�];�m��eS�VY�k�lص���               �<�qe���2�p�y&#�˰�!�}��D�Nz�6�iOw��w�m�m�n�&ٰs��7S^J�>�,�cFM��#�ȴ�e���2iȸ��|�������^��[��3_��                ��s�r��i2�<��8\��$��N�.�e����X/�������*�nY-�6� ��A�Pp? ;��3CN��2m�ݮ؞)�k�/��8GN������7<'��{R�X�T��                ��vsg��.���%'�;N�y�$��֧�>'��8o�����-��c۫�����ן�'7>�*�@���mΚx��;���lK�a�8dl���i�u�U�^�߿����lj�*                �{5���'�O>]N�x��+�)u�ާ����xǌ+���G_��<�ʟ�ϯ�U:ҝ���.��)�g���.����dJ��c�뱣��~�q������/=$��s�`               �Ɩǯ�v�\pę�(�H��'�L>��a����������S����]�����UG]l�2z�(h���cft?�|�����G��R�n_'               @.���ە��v��r��i2ٲ�EG�����������ꇤ=�!q˂��!c�W�%Sϕ��������G]"WyQ��
���gݫ�               �dP���3{�Q����#%WL:N�|��t����~#?|��dkG��M�
�v����F.�v��ʑ\dWu?s���[p��߾�}�               ` K�Iy˔s����!#
�I�*L��g^ݽ2�/V�N���cUt�E�}H^��x����#/���o�۱���O_�A�㫏���-ym�z               � �ESΖ�f�SF!q����ێ�T.�z^w��������亜n{;Jɕ�/�[f]'C�
%�Κt��6���s��������:               ������Sn��GM���(��Nx�\>�����䑵�K.�ق��ᓤ���ʌæ�{��ws�\t�Y������<*               @���g�6y�1Wu/z��c��J�Ok���Ǿ*wm�\�swW9r��7�|���+؛�-Ç�)���I���l��)               @T�8v�T�q��<J�fgL<I�s��|��~/�&�
�c��3�ɱ������!�Fϐ�|U���c               ��.n}ñ��l�p�#ؿ���� �w�4<���Z�:g
�~���~�JNk-��n����'�F̐���'���               �lW8Z>x�B9r�A�l۶M�7)��	�r�Kߑg6=/�`��]��-����g^-�[n��e�֭�����H��ˤv՗es�V               �儱3�γ����a�ޱ�v��}_�oi����<:�i��s?��n@��j��q^��8�XAＱ���۞��G�O���噭/
               �io;�R�s�lq�#���}`�����.��#e�	�K�߿$��e������_$�G!����{t�w��㮑_��<��a               2���W�m'�K�{v��իW�Un��y��Y �yB����=�3�K�Yp_8F�\T���s�r{�t*%>UFN.�y�g               �'G))>�6�|����������HˇfΗ��(�;���Wp�2|�|�J5h��wz[n�����L�!G^'_z�{               􇤛��3�ʹ�O�ށVnߗ��N�<�����嵝d P��F-��B%
���r���*�}G�S���w               8�|���r��������o�j��H��_��;��@1`
��G!w�WJ����޳�2Nn�~�|��               D�I��YH�����r�u�wJ񔛥��/ˆ��2�������.�!y���9�r����&�uG\&����	               ��r����%轠+���-��y�|v�
ّ�)Q����A#���P��֟����wR��<~����?	               �[�N�YΜx���u��7J��;��#���rIy)��H�%��W������������e�ϖu��dՖ               8�wͼZ�>�bA�����o��H��Yw�g����_�?E�ஔ��3�ɴ�z'S���TJn��v��Ε��k�                �cWm�u�u������(�+�}�|���KTE��~��k�Ad��ޣsW�Tw�|��#|�               �3a�XYt�q�#�[n�}`��3��9��L�3'�,����DQ$�'�?^n:����V����{���/���                �.�Mʇ�-���`A�d��ޣ��K�w����e�ؾE�&r�a�Ce�wp�F/e�ܾg���9y�q����               �q��7����c��/��BwG7[v�퐊��'K�R+��|��/"Wp/;�}2�`����(��8�ä��ۤ����t�                ��?^�>�bAﴵ�u���Yn������3�ڶ��{��\�$R�˦�/gN<Ippa��Ǎ'�'ﾪf��7J���(               ���y���9���-�ە�}?�+�w�ۏ9F�ɤ�g�u���&k�^���L�ݮ�~���\T��֥Sϓ��I_��                ��8i��(&8�(�ۭ�����o�?��uv���D����[dH^����Tn��6O�U*~�1��R              ��9i�rɔs�r{��M����H~���(��8v��3�T���Yn?~�L�4i���p���+�O�H               /�rd��7v/���Z���-ǿC�ǟ��k��-�c�ܓoXT��=���V��K����6               ���#/�)�'	,��vkH^��<����W%l�ܯ�~� �^n��ܤ�:�R��J              @<&ˍǿ]p`Q.���b��r�s��W��&a
���t��c���@(�����3�{�~&/m{E               ���1�r�W(ؿ�Pn�\��ͳ�����Y�j�����"�!ط�Tn�3�o8��5               2���>�2���r{�s'�&�F.������Vp�s��ΙW
�m���{�A=u�dVq              �q�s�J�m���-���>�m�?4IXB+�_2�\�?L�f��n�A}�˥�O�
               rS��'WL�P�o����I'˄!c��%��m	��3.��@.���舳�kO~O6��"               �=�O�@��
�l ��-G9�^7?�U	C(�S�/��N�-���rŴ�kO~_               �[�b�o=�-�7����L9G����ȮT�d[(�+����J�����/�o<�C�tv9              �Y'��)���-W��VA"_.<�,����l�z�}D�09}�ɵr�5�`��6�yd�              ��q��{�������M�(����ȋ�Qp��s�u\�n�Xn���Qp              �!����I��%��֔ᓻ/o{E�)���'�!�-����i�guOb�R�              ��ϖۓN�+ȑ����~Fn�����#��~��J�I9s�I��               |�O>]�[��ۭ�?C����J6e��~��h+���L:��;              @�,���+�G��?d�L>9���g��~��Ywq*�['�I̮��R              ���ı�J��j�8��Rn�qڄY�Yp�(���)q�r���s���g               �]ǯ�n�2�x��3?����Vp?a�LqW�*�����;��;              � w��$��Xn��}��y��ueeY+�7�h��8�ۭ�fP              `�5h��+-q�r��pr��i�����?ɒccZr�{��:z�TI�����              ���������\n�qܘ�s��n[��G.qC�}�����#��U�^               <3�&qD�}������J���a�K�qB�}oS�N�              `���Ů�*�Ȍ3"Sn���8"k��J�}���'���l�x��O�	Q?1�Y;:�պ;����w����cG�����*�|��:"ٛAs���������i'�����&{E����o�vl�7G�g�҉�{�o{e�pI���ӥ��傴�ou�L�����s���~c���<B���gs�/��9j��_�����k~l�����3�|�zIIӖ%K�8��ma�G�����k\QS�"���ʹ_)�O�?�~�߳O'҇����9���3��y9v�c�3	G�/�����9g��_(��c�w҉#�#��7�;׸�����sV����9�N������>�%�k��$��g��ϙ�d�!r���+�z�����MM�#\ϝlN�f���y{����%��9�|�����#)���W����1��1�j�v��_�{��ҫ<�{e��k}���1�~a��ϻ��1�W�y��$��Lߗ�xW�y����'��z�G����J�ɚ7f��m���gp�c���~�����z�'����m��ǖh�}�Ùh_���c�U�X{��_�9�ń��k�gz�7�~cc��e���=��q     �@���ܾ�����y���kg������ãW�ΤիWSn�#�M��|��JK�Vnk�����of���g>l��x�<�f�!����<QN��z��R�>ٓ}�JHKqY���7��~e}ٹ�/e���&yG�'&�Z��-*�W�����~������ޓRsu#����^iՔ����?n_��{KMŹ"^���f��;Ot�hiNh������}��f�����GYkm��f����os�􉯥K�n6���%���׿yC�O��7̣����,����;���E�jy���'��o������3͋��ߣ��Z.�����'M�~˞���>�h�.9Ü[�h�n%��3�(]Z�	I4�T��}_����U�-{��b��md�wfܧ��{�K*�����^R��YSO�3�o�Ge��S�)�Ŀ�E�}d�7sν�X�X\�����~���yT���s�Z�E�n�S��W��d�6����}�^l�����u��﫞�-��U�����#{{L��W�,+9Y�Z���!����^�_L(�aAE�co�������Q����$ǌ{3��%��3�uڜ�|�|Ұ����}��%K������y��~qku��%U�ym;G)����|��+f����������R�����ue'(_���=     @�,.��J\Pn߷ÇM��6>'���7('+qaWn߲eK���r�5q�8�|_��u���=o<�R�K4>h>}�uY��}GꔨK��a�Ӻ9���ȼ��6�u����?d>}�����ڷ��e�����Z�$���5��Ջ>���d��L�����rWYY�� _a���ߛ�o�/���U�(�R�ھ���|h΢�A������͇�W,-����k�/�[��|����s*�e_T��G��͵�0?�3�\#8(�z�S��*�������|�yu���ܳ��)ǩ6�9oTw��))��_T�.��XP��'��ֺ�O��T��﵂�ړ�WL�wί�?���Դ���J/3�_'8(��/�uG'�_TU�Z��Q���7��f�'͑{�R�z�A�d��ʝs���f�����|���s��������7�￿x��W�l�'�����O���VZn�'�>��A�_����d�)�����7	z�d����Tͯh|%��+�� �MK~�u�3�ko�'���������5A������ue��|�Y��=�^1����$*���#��E����R���}��y]k�g�     ���S�r��M:6w
�cGKPn߿��$�͓N�K�}�����ŕ�쏯7��Ѯ|YKu�|�|[t�쓧�u�d_R�����zE��Ϙ��V����n ���ٻ*�����!�[YcW����|�־;@�Oi�w�\������C�������*����Q��d�ߔp��K*�~�_o����͇k̜s��s�͸,�'�}�w�]\U����zEu/�o3��=fα�
�������PT����zs��^4�m�-���9�d��X�E)uCɢ�_��כ_^��|x��sn4s�
���>���-���.�h����z�U�/��l�)��EV�����)%7/j�i|�=űw�9�]��}�QN|���#���:7����?�ޞ����ʾ.������d��mJ��������z�+�lQ��֚ү�"6��}�E�9Z�S\����z{��yym�ה��D��狿��έ&�����sq�--ե_�J��e�`��9�vW�ۊ5|�?����z{Aԭ͵�_�Z�!�����(y��������d[K]�״/_1�~�      `���ǟO(������g��~��:������fr{u���QJ�����z��,��km^V���*Qc{I����P���5Z��@�W֯\Q[����?5s@|n��Kf�?����~�~AE�=-�JՎ�q�K'{)-�	7����Ζ����M�_h�.~�S��s��Ō�'�$y���`+(��s�Ҳ��1ߑ_8J&�b��SII�e~U�go��W�ז?�k�Wd�`/f�?-I������~"<�����J7���f��,�KZ��\�wIQe�ի��9�h�+{����;�9\����g璹�u�V�>���k�/}�Ow��G�b���ʽxOA�_����KK��v��^M�������d�����{ EU��k�-?��f�5]�3߿�J򒠫���E�o�+;������ڣ{1ٯ�K�K�5���_{aE�m����V�т��}��d¹d��w�jAeÏ��U��8���s�������Z.�S��b���Wԗ���Č{u�`/f�YS���s*��=���?i�Yt����3      ���bs�(�ܸ�)��U�����&���9l�
�x������|^Q�L����KK��\y��￘��`�����%c��ۻ7ז��k�AGe�=L��|�{+�ޙ�}�ۻ߳��ܔ�qOٷG���yXz����@CƲ��o�+;����s(����c�C/����n��>,nx��f�پN?�(E�t�.�{�w�,�i��>V�=u��K�N%��N�0��_=ǽ���.c�ۻִ֖�c��&�)�n&������ej��5+���N��	��|����w����fj��)&�sR��e�1�~U��n&.�a��Z��lOR��p�/i�W�	�9���p{�����J���鿤E?�'Թ%e5����1�k���o)=�����D:}μ���p�Ǟ��3�����XA7{1S��3��nC��a��|����d�7�X{�����F��s�/_��}�F��K�K��o�R����_JJ��9�h���Pj�Ҫ��nʌ{�%      x�Q�r�f���{gԠ��|5�����}�p��7,���co��Q�9䪹���X���-b,�-�R���U(1���g=׽�4���E�溲+���@�����Ġ���,���S��⊚�+<�l��}@�.�P(�������1Z��^�3�Ќ������2Yn�aߐ�3�<l�}n���3߿\��2�bY�
�=漿qMK}����4�g��L�����zKEY]Ƴ�+5/���\ĳُ��3s�+�t��������{�-�_�bi���L������~� ׽䎊̕�{���YV|y��<�����DZ���I�L��{̯�Y״��
�ҏ(%��KVZ��]?E�+X��ٯ�/��K�G�K�9�^��K��g<�9u��|�]	y���͸W�z��/��]���f�Z[~��͸��m;�oL:��6�L���|��.�B��#\�mWn�7xrq&��=�W�׵)_�9g`�	�f�orU���2Wn�aϥ��y��z��d     �Y.��)��ް�쌃�܇�p��r{�ˏ}���W~G�N�#e�+�h�.�����Ę�ug�J^;��&ㅻE��k�)�c>��Ę�>�:�f�p�cޢڿ7W��%�I����z�U�/������֖�1'�ߔ�]ǽn^e�w=��-ե��q��*����]��*���]U����V�����K�kM/��X����֚�[�K�I̳�w�k��٘��]{!eK]٭�`s��>���"�9�f�p��^��ZW6���&yGb���{�V�ϯ�|髇]ٷu��^���^{	I\�����l�Ӯ��R[>[��W1��O:�z{�K��i/�[^]z�(�+3߻S6�<���^��>��|�ՍZ��={W�;m��g��寚�7�����^BT��u�un�SY�&[���[su���1�k5p���oJkGԍ�b�l���W�q��`��     ؇�y���)�����q��?JN�\D���
���<g�ܪ�U������o�Ԕ��<�wK\��rny��_��ᾖ���E�l�+W/.*ox&ۻ-���fKM����&�+��_��t�w;���[�5e_3���Hl�������?j�.�����.1�E�UB�Eu��c��g?Gb�Q�����g{��5����|�=O�J˒yu�e{���b�QR$1�|�DQUã������_�q�l�}�Ĕ���.�j�C��;���׭ե��xS!1���OQe�ﳽ�u�i�.�5ϠRb����+*oz(��]X������j��Ĕ��υ��ym����ҥJ�$�<�KK5>�����n�.��(�!�)_�E����~�*��RSv���?$�ҾԔT6�2��5�)i�)����      ��r�J����egd���troa�����X@0]�r㶱+�ڿRN��m�U��L�N?�i������y�Ŏ�x��ͫ��K{�6n�<�����?��w8�b�}J{ύ���1���~�NqR�)Q�w�]�޸ulMX�O8�S���>v��1���[�-k�:���$�7(�r�vN���{k���χ��N��p�f�&1c�1_�m���ڿ����]7�9g�Č�s^�m�gB�2�7��d�)1c�s����a����/iO�b���3)�_ߩ�C˾ӑ��k�3��H̤����/�TX�w�?�.�y��~�Č�~�;��Dh�O�O�i�͜猗�I��4�k��_���d{^�{�����֛��,��낮OIG�}fΙ(1��N�G�ڿ_��iݑ���9�M     �~�t^�@(���q���{�h���%(�c�<Q^�d����[j�Zͧ�3���P���[[��m�~��LR���{{kk��-�WI�$���ٳ�酵{k���Ҧ8��h���̸O���9u̸���v�P�G�̾�Ζ��5e�q\�._�w�/jJ������M&��}hE��$����K�t���y��m6�W��H��)��af_RҴ����^�Z�2,y���w|�#���l3�ۋz�Gb&�%�����EE][��U}C��$,f��D������no�.��(}�Č+���~WX�/-m��\]�YQ�Tb���S����;�ڿݷyme�j�G������3��?�i�Č#Χ���k�6�֚��1���     �n������q��w���~2>�ʕ\A�������K{kK5ݿ ��'|�:�e�S%1a��d�ð���D��+$V���6n������Z�g/.p$&L�6n�ݰ����5鄲�&{�������H%��dZ}�L9�sRz)�oٰu�}a?�n����}�����6�Cy�z�3���d��u� ̜��J}-��᧺$/��Ul^����}�ֱ_�y�^��wS�)����0��4|ח�~R��$�ɏ��Y������_�yt*��@���*{�۝A�{�~��A-�������|�;���y��~k"�>�;d�ZwNj�yt�h�k�o�}�Ą/���ӡ�	��.�Z)�O���df�wu9N��o���)t��'�w'     ؗ\�Sn?t�b�./�k�e�������W����C[<�j�U)��a�T5��RS���>_b�U*�WU��ZS�;�D.��p��s��E�j��R[�[3
.��0��+�����7�i�.��(y�ą�/��r~�����[k��E_%1�D}1���{̯�Y�RS�3��[%&|G})
�/_o�����m�w�+EE-�����޽��c��<�wHL�s����z{������O�)1��|#���{�U�͸��yF�%.�ܷ8��{�U�͸����&�	��o���x��{KM�w̧0'��s�vw3�|ی��$&|�7
����ZS�-s��Ą�����y�y����^@~�Ą��TT4���<���k��s      v1�(����|%(�����q�(����z��t��%"����Hl
�	ID&{s�c��O�]Id�7��.��H8nt�W�d�bSpO*�{��JIl
�	':�w�9*>�����1����>6����w����ͱ�;�d�U|
�	��cSpwŉ̜�'���]?B�^9�k�cSpϋԜ��M�=�ߖ����*6��R��瘱)���V�����=��;     �����o۶M^x����.|�ea���S��L������TD���o_�e�Z? JI�[�����q��}��#q���y���JD(qВwW9{;�׷���D���|�M��Ӓ>l�a��P��sܸ����yX"���:&�/�����W�xj`��-m�����KD8�����cܛ��A�ID��{ �#�E<8�;E�N"��L����{s:�����H��\7�ދ�����ɾ��H��1�-��32٧�͸�Ǹ�̑�7IG�:�׵�҉�dߕп������~22٧���)����       �#����)���l�ۭ��Б
�nفQn�_�NA���_�dɒ�4k�I�d2�b��D��_�=���9�(H~�#�#٧|�r����Oq}�{��M����0sNd.u�n�ob�B�7�<�2{ɒ.�]�zV���JIη`R�[[��)2']�n�܄�RJT�Rۏ�֯-���y�3t��緬�i�}��.�ו�쒈x�m�Gm��
$�u����w���iuK]�.��`�qf�o�XT�&1���k��K�+��J�K�����~�DD���.�)msD��K��e�%"JK_o�)�b�sFJ�K����;[6JD/_�\S�Y����ֺm���s*�6�Ԕ��3Fr����ŕ��$"��6�c�zs�+9.���%UկID��4m1��u�X;^      bnW�]"����=��q�����ȼ��'���_[�A�i��DHii����J��Cڗ�%B����w6ה�S1xc�W:R�/^������u�2Qr�9)}A"�;���\S���,9�7�R!EE-��������̸�T��"���җE�Q��|��W�c�Kf�#9NG,{{AgKM��]<Nr��s"��R��k��~��8��_��Qʞ��"9Ό��$bQϙ�I��ܸW��?Sr\Z���ؿ1�-9��D�6�^�|�݌��e��cƽ���c��_��qE=�Er��      �c ��)���lu�3^po��.����N�=��r7I�(���{9�Ɛ�T�����s��!W�Ȭr�OZl�9_pW���>��JI�W��s��Z%$*2�����},���I8�J��|�-f���A(-�r�A���D/{3�cq�U����)&����q-�ϩ��(~�1�s"��V��s�������72AG���M�*     � �:V�r{fl��N/<����v�|O\Ǖ�`��Ք�3d[�������R=�*��g�S�s����iN�:��'r٫��{�U�D��>��}FsΑp$z�^$.s�D.{��	J��}��>��?��Q�>&�^3߇&���Q�N)�c��E�4���`^]i����x���)��d     p`�Ђה�3'[:d���k_6�o�q��%�l�}���/��r��~W�1Fvi�����bQ�Q���s�04��Ik�ܸWJ���hO�ȍ{c�Ā/~�O3�8��/ћ�ͤ34��}FN�S��:��gL���q���cp��EG/{3��p����c���7���O�{n"�츏C��
%b̸��uϥ#���	�"zߧ}N��      �~�&(�gV���/�[�wn�|�=�r�ĉe	�뺼Ԁ�z��D�Js�R-�jl�/�i=Q"�f�Z#�bpm���7�k=.v(Q��ޜ6����žM�!QJ������tVS������*��eoD�9e�8��1�}�G�r�J���9�J�{R1H_��e���X��H�h�9�Q��͸�����74���|���ބ��^     �0�E�)�g^�.t�J�}�΍r�D��̳c@k�8�;W���{��LV	$1��s�D��e'��Dn�LPN��_YW6��%����;%��Jƫt<VwD����/=Lyr�Ā��K�ܻ�rDJ��\F��	Ǚ&R[[>Li����K޾�u�J���~���~���Ʉr�J�|�swv�H]T�)	QS$B�����m2���x�{I�s��`W�hL��-Y��Um��1(S�ʙ�웛$�]M��M�J�d��<|� �<"���o������}���nYk^k�~�f�OL�������$�8Pj������ʝ`��#-нHJ����     ��@��r{vdkd�ྦ�5�*����W�����SK:�D[t���z�D@�u��]J�{O10�<���X<���i�D�뺁�������>_�q�w/]tgK$��|_���
�l����K�w�=��c�T�m�p=�� �єs�	�s�S�({1�����yZ�9'�<�*gd�҅��/���WZ��9�0眀�����[k�'ϯ�{E" O���>�԰�e�S���_�H�&{���{:��T��.!jHk]ٴ����%:�;Or�@���~�\��ԗ�XP��D��c�iJ�k��&�8��9�R�+�Kf�4>-�eĆS�(��ۅ;���;��[��'��D�jO�lf�>�m5b?��9�G���M��	�m<�|�7��I#7�d��>�Kt��߮{�}��[�fbM��ɮ�D��Wǜ����v����Ao�w�����n{}�����$&�X7Kk���ۅ9�-�d���W��=7��E"`em��J��}�.��{     �Ly}�z��R��F��M�={^ޖ�JJV
�/o�D��M(�g��[#ѱB?�X Q�T�I]d>��D�R�R���N?�7��1b�O���ͧߕ��\dѽ�0]A�Oڌ�D��ߖТ.�]���sTwa���}��_�U�˦��������U��W����3��c�!@\�}���e� 3�/�]g�%�C���o��/J��.�K��Hb��9AJw��zv��#Q��˂����c/�
���k;�WH�cm�o�+��Q��w��.�������#Qp7�%�|n�і�ƌ�\�}$
��X渷c��;I��k"D'�}$
��;�ڿ��y'O�|M�(_�6w�X��s��q���d�m��(�����.@o����B���>w�f���>m����S��>��s��č      ��}eM�Z9rd�n6L�=��S��=;���_�`��r{v���\�O���O"Pp���ղ�]A��p(oJu��ه^p��w޺V�;�����ƽ��>􂻽�����Y0�3���!��̸�]"Pp���j��Anff�7ս�Z�W�:��������xk�}�7�����5¾0t�=�>���۸�*��f�ˮ�����{wHD
�̛�~��G��g��@K��9'w�w�(����ص{ΉD���k��^�^Y5P�^w�M��f�X�u��d�𧱔t�9�7٨#�Ue�EMA
���v�V"����h�	;{ߗ<7������5;�V]!go�7��O�s�e	6� �xe��͸/�{�=�^"!ظ��XkK�}^��n�{���D���s      2奭�D��N�=�^n{5kYg�ྵ�M6��,���(�ܞ}�m����O���~s$���;CIq߶biըy��e����L��m�ø ����$,��ءӁV�2?���חVVְIB�u�kD�~������c���AN߳Oj��{j��̩�� !�8b�[E��A���7�m�]�dp�����MM�/_/!�4r�UZԤ ������|t���N߳7s�%+��&�-��*�֚�+̜�U��޲s�07������MKN*^�<�[謨/�Di�d۝~������y;3�/h�-�<��.�+|[��]��d۝!k{�?"@�y�s����)��^�-�.�Pi5#ȶ;B�sl�AJwy�{nӲʩ�U�/I��kJ�W��	�m������d��g�XZrԼō�K�̼w���� ����3�p~/�i-��3�5�����ӕ/'�6
�9��c�{Js]�̢��g$D��JOU"'�6
�0��c͸?yym�q+Ꞓ�,+9ټD<5ȶ;#p���>�I����bּE���߽��g�6�q�赕9�?�������M��,-��ٳ�l���e~�#���+�83�d�P�^к��X��� ۆ�=     @�<�e�\:�<����������ܭ�7=/>S�F�=����$wm��^�Lp
����T���2�~TB��� �٢��C´9�!�C����t<�~��]�٨;{/����'9}��U���}���%L��P����9��S´Ɍ��y}?)t̹N������"-*���f�9�q�)�.��Wf�wx�s�HB����e�wa��*a8J�T±c�\�䫻��9�&�i���Rp7�Z'���8["!�N�c�&/�q?"X������]$!r3�N:a���s�[���l������t���<����!�
}ܛc� ً6�����|v�����]*`��һ$Lv܏q�y;{��tڷ�io�9~��~s:��Vc}_ӷ;{ϳٿGB��|P�瘛�v+���t�f��H��]Aߧ����;d���oiV�tg��E�)s΄ K�RJ�Kޡ��(W]��I��|�c�C�;p��q�yN���!g     �)�6� Q���F�=Oo���[Y+�?c���[p��{qr�-�MH{SN)��������lKM���l�	i��%�,�hS����D/6�7��}km���IE�K��L�)�K�6r�����Ma�,k����� �n�]��V�����u�ZԴ��!��e���]g>\d�:��;�h[W��{��̩j����fyM�Ufƾ0ȶv%�г7��Լၶu�*2�/+����+̜si�m�u���a�s�t	��#������V�m�.�܌�˃l�ar����X;=oD�mq殬^�tne�*	AKm�e���A��wG
{eS[~:2�&�;���>֊�v�|s�{U�m�\�S��������ۺ���Z]�4��e����� ����N�6ۂ}��@ۺʹeym��a�,����<ߗ�lk���}k��>ض&��[��|nAU�����3D����=�e[��!{qn\Q[��yu�Il�Z��A��F���O���d�y��#�֚��|��Vj�~D�*��w���9��e�6���IG]�\]zVQe�%�nf����޽XD��;     �M�h[+;�vʐ�`���`���?�<��<�){8d�������9�r{���>�~	2l�!��犓�ru���Zɲ���:��.�(�;%l�L���A/���r��|z�dٽ�*Gt�Tu��ׅ�����`�cm���u��r��Ւe������&�_��¸����sDJu5�O���^:�&����>e~����i7GT�]���ĥ�w ��*V~�C=�syн������9tg�{L��d;����!��Ơ��q/�Tʷ���lg����Y��7�qH�(�S�+�,Yr�yd��83���1�v]$�1�?�}���1��F��Xk�o�o�C�~��{���#�D���Ι=��Y�2��{o/HmS-���9ag�z�вO��J��Y�ξ��<����+ʮ7s���?�9��9"�h;�iY�*�f/��b�z�}��f/ᆿ�ʦ�wL���&�ӳ��}K��mQ[U��V�������P��Ju�^����lgo��I��o5�>`�v�	7�C����&�S��Z�ze��^���A��wl�B^,b�!f��fJ�K�,���e�u      d��}yj�sr�ēC�?���i{M�tl����Vp�Wml���ٻ���{���3��� aWA@�խ�֥�V����m{�׶�%,���mKo��V@	Xm���.X���"��Y	ٓ�d�s��9�P��d���9��w.�I���9gf~�y:dl�h�6��v�FA����7Q���5�gΘq��5�%�f,]�M}��_��h@r�.���j�+�6c΢[$Kt�K��0�8*�c�E{$�jc�}����5U��3�.Z$Yd�oU�LJ���a����U��^7wa�e�T�"EK���ѩ~~],��>���%5ճ�!��FɢDI���)�~����ŋ�g}Ke�ɢ¸�f5��K�4�{��B��wT���,���q��B�y1��*ھ�>��dS�h�!r\��^����g���U��d�.�V�����;���5��M�~�>��dQ��l��I�~�+���~��H������{��1�ɢbK~���SS�|7d����d_ �3'T��T}�=ɢ�����OO���\q��I3{㌉���B}�mɢ���ߨo��T?�5٫��z㿚sN�0�E__~S����i�����\ېf����D�����$��u�/Է|v��_����W󽾹ė��?%�W�[����E*���o��T?����      d��9)�Snϭ5�����Vp��4o�+��0�_�r{��v�ol@��+<�����O#�a,Z2V��/|L����Y�ؔ�pOrÛrz%󰩲����i,T���V�KT��0�c��6���[U�}jܗ�>���U3w\7��G%�̯�������1�ܐ}BeoƤԗƅ�%�_�`��kg/|D�`���?QԟH��.(a��!	�������7K�g�f΂�K,���c�T��9F����xX*��4����+����e?��-�>��1�0������/N�*�_�s�6u���dAMլ�q��t��F��=�����Ӛ���θ~�}�*�o"W�s7\���u����>���ߜ���Ϟ�N�_I�����\Уr��N��$�c�,�������!Y�淙�?#�c��\L���m��SܶC�|������ۮ�����K�f]��}e:�pÜ����u�t��|�U�}[����vɂ���3Ĳf�s7\�������)���Ըߢ��m���|��Ι��1�0�̸��B2�0��}���Ru������,P�k�QsNZ�n7����wm�X����*����7f-��J�����ϭ�VB�cA9�px�����5U�f�]t�d��9N�9�J�u��g     �I��\t�(������.v�Ղ���ײZp�ܞ{���?�!;�v滢�rR񘔏��o��9�1��ɠ��Y?T��w�9F����5����X���N���L˺qU�����)� ��K���1t�S�	�k��hW�KN)��1�e˗T��еs<)����{�+�o:��U�^�	�k:�j�9-���q����T����9�ZR]��M����.\��J��g�%���K��F�2�YZU��k�.zX2hi��o�'3��9�.�4ǃ�;"���a�S��d�j�T���$��VW^���Y:��œ�X�ǽ�眳��^��ճ?vݜH���ò~��1��s�Q�dߥ����,�0E��9'���%�t��+���î�]rv��[�,��iVl��.�R?�Ju]\��1"fBv������61���+1'ļM�����௒A�%_s������n��^]ߏ-M�d���,�Vu��w��E�J�TU~U���nP:���K�wɸ���7�Z�����R�߾l���i{�Y��Gݱ���i����R5�Ԝs�d���K�i�b��}\e_�죝i����K��9�Z:���Z�F�*{�;�i�\�N�}_��S�9wJ��-}�N���RqI�j�I��n�9bԨ1���|���g�������Я�[���      ���ǵ]�e�IY�z��s�/��m۲�5���{ ���_H>\����������!ԖV�]�����g%oPTW�..k�XrM���j�,�#j��^NN7{�(6E�+�eb�;;{ӬR������������mi�5;{�|tI��k3���~�%7�̾��6�?�[��s�i�g_������L��u�yE]m7��f�{���6�f"7ب�O����(4��gMu��s�"��F+�U5��v�d��}:wMgoY�?�̟5����,������Z�#���6���2����4��R��_^3���/X(�7o^���V(i���mV�>!���;�4J�ҟ����}Iլ믝�p�8�?��_�X�L�X��v�֫k�����'j��,��ׯ����0��������N�X�#�.ʾ-����o Vsν5�+�s��E7:����~���4�j��^:�vM���K�{=�W���8��^��,��=嫳d&�=�穯�I3���N����#���2G�_���r�5��&s���Q�?V�����if�����OّiC��Ss�]jΙ��_f"�#*�~�oN;����}HgTZǰ�7�?/V�7w�����ѓ�@�?�����朳-�a�P����{��ޒ;��Y&�?rt������K�`�m�t�7R���s.(��֟H}���O5U3�5u����٫��qk����ߴ�^�ۣ]��      �NwC�Qp���+�J,����j�=a&d՞u2}���:��ݡ1�lߥ��e�XoƤԗ�$n�`�O7WU^i�eάY�ڝ��W�>�ЫYr��{=�&n�W�u,{��T�W�c��3��đ?���_;�4���0�r�x\���H���v�?�������-j��Y_���Չ�f��ӌ�u�e��N�M�6�%�DT��Ei��^�[n�ye��?ө�o��sj��v�!r��[����Ӝs��%7/��y��,����:��-�}�)��V��q��sӜSHw""#��iG1��[tK��+������f'���7�<�
��:�v�x����舆X�t��+��Zps��E3f|}~�ߟ��O�D���x��[qϸ׫:w&�*����cg/R�εW���k�����;{G�غi��������ץ��5f^���k�2{�'��%+��x��s�����t����DH��S_ͺ���o/��ti����Y�ȓ��Us��ܓ�U�"'���cAi�����u?ð,�75�g^v���_���N|5ճ��j2���_���t��-Zb}�e��1�Xe_SU��s����n��k�č6��Lw�xn�:���1���U�?����^SU�e��_�`�4�l[�>�̉�iܷ��^�5� �`�yn�t⨖��t�������N|�XS�>;�˝8���oS�7�9��BG��ɄQ�����v*�[VN1Ͷ5�]����4�����x@&��u��ڹoބ�-��y��kf/��������ڷ�2��;q�.�      ����W�s�~T�R���A��=^hX����Ղ��l݊��)���s���^au]�5�U��
�����>�����fqlɌK�R9�m��99Q���e��J�5m����C��ٷ���W���̂�.���WV�o�L�8K�gOR߳Ěa8�}c��~��-L��pKګ~%���d�L\U3�O�Ŋ���i�wӼN]9:��.Z�҉[��ש���_N��|�5��/����X�������T�s��;�_P�]�J|�p,��]�r����^�ȡ�}��#	�_�����P��_��o��f���1c���um����z��j���Ɏ�/��2b��5U�~Z.]�j�57]�����T�z���Z���q�"�ʾ@|6�إ�\����[4g΂�T��h�̉�q���u�l5�8�lZg�K�n���v�x�\�!�۾t�쟇|�0��Ο;AԸ�K|�a9�����7S���}�^��|�#�S��c��]�9?���Bu}ߝ�qt���������8�}�˲�����ee﷌+bnS��_&
������T�s�-׍�G����Wט��e8@�����55�\Q>Ցc�|�+�~k�ҪY��&�gμ�3���V={\²n0M����7n�F�D_c^Y>͑c����L#���s~�(LT��}͍׎5
�n��u���I�N�]*{}����Q�_�P�>øT]�o]2��}fA�Wo�)�g.�Sh���0�p${}��Έ���5�|���}��q�E�9�����T�����zˈ}S�H�N�=*�Qwe��#
�q�X~�x�@�7��oJ5�[��і?v}"a}K�9e�.��ܓ�|���-5Օ7J4vS�v��M_|n"a~�ˑ�{ͨ�k     �P���*[;v�	c�y��(��GW�Gֵl����z����-���"G���)���i��T�K���J�I�-�(����1B��n2��T���a���ؼꓟ������o��G��,�\�0?jXVa��(�ɋ�Fq�W��U�G8�����2���8����+�����G��|��kj�-�"ŗb}��c�gﾝ V��O�"g���[7��~�������3ꈦW'{#T8]�j����ٻoܯ
6˻Ըw.{c������Ú���0��{:G��7o�!����K��5�|���bI�g����v6�2��f�8�����ͻ�:ǯx�����+�G/Qy6���V�"'�~�ϑE���o����H)�9��^��*��TUީ栻;Ƽ|8�/��O]�}ֲ�P��h�z�g�y��Zj��ˎ�Ù�M����4�d��;���p�/�G.6��Y�[*{�ذ�K����e����jܗ���^�#K-��y�i}_go�uws׸��.��o�RI�{����V�T�;:�rܷ��Ï�aN�{1���?3C�߯�_�ƽ�n�8�ҌK��[��������^�ءo��s,�u��I������L�.�4���e_]=�x�i^dg�>%�����]�'�/�9�B��2Jԟp�/����^Ŀ��s􋟜7/z���٫�/��l�2?���8���
5��^^������!+Ig�~����W��2���u��Y��5u�����R'眗ո7]6�_W��B5���B�PV,����?�-5������F��}��w޼����Uޟ���)}��3�V����w�J��?��7չ�5�����Y9����Ǵ]`����|J��eN^�l�hp�K��i~�ߙq?��T�7,�_�5m��p���x�!�g�5�˜�s^Q�kj��F���*�tw'KR��"���7��T����sX�����'�gT��v<{5����     Ȥ'v=���;�vwy��%I�	ɶ����{��E{k'Qnw�����/�?d_0�ߐ>�t�����o��e��3�7��]\U��O�MbX�b�g�	�\��Ԅ$N��9>����d�K�+��m�#-h��"�.Z;I�8RE8ǧ{&o�?��O6�|��^�K���%b��o(М�^o��=�����q�.��7���"��e��w��uZ�2O���#��g�W��������=��+u�ܫo�Q�R�ϚX�ڧ�C|��l�?{�gM5M�T��!V�w�94d�eM_�������o2��>�9��5TSU�Be�YM���%���d��p�X�s���m�w�jM�䍰��}X��ա�r�C;�$d�5�����^��>���MÚ��7$v��Rd�z��eK$�3*����l��;�{A�}���u*��&V���g�T�n<T�jNh�8~G",�#)-x�QQ+!���ʅÝ�1%)�������.2}�:'�}��8�.ψ��|ߩ��v߸���q���^g�k�V�(�x~�*���h�U��^�w�U�SU�'G{Dg_���#�!��q�o������ˢ_�|�)/����/�o�^E=E����|�e����t��.�>n�*�&�ġ�#��٫k̯vT��ո_�������峷�Hf�桓Deo����3�1��^�w�K��7�Ow8{���Ɛ�b~Eg�=�}�#{1���<����3�H@=\n��[��P��e��^���G��Qm������v�yD2�Ni=Ϸo�pg��+)�]��F�_W����ڑ��5U�W�Vd����T�U�u��M1�տ����'v*{S���ǽ�z�K�����ڵ#i �/��t��}z�[�Iv��WO�o��B�����N��d�>���_,�Cg�>����:{�����ۯ��0{     �Lz�����OHY�sk�Pnw��΅�ܵ'w� �:�CR���L����ѝ�/w˩��8���[��.�]j?��w����^����[�o�to���^���ac3���]��b�.��ӯٗ}�%��w�ʚIzܟV2ֱ6��`�[�5��~���ܜ}��'����E�KTڗ$�����F���^�4|zi�(�\b?T�����h��@��V�Mz�o��S�{_f�H�}����^ddx�?��ӝѫ�䝥�[����2�������qq�+�}�?{�F�,���\��l�
{�Opleٷ(�]�Ҿh���]3�l���sm��d}V&��W�6.T�_������2��������W�5�Y�&8���[�����/�}�k�d�����sܺ�l2�Q��^�{ѫ�5����L���n�~u�Y�VsNE���oT�){k��3��n���F�ֳո]��&�d��P?�e�/��H���X�hu�Ee?1'��W��~��\����V{����a9�J�X]�4{}}����sj��7,     %�DL��{Y>�K9�v�ym�&i4��k����g�_�˦]���(���̫�6����s��r��+O���>�6�-n��6�[�1U�ͦp�+W�Oҫ2�7l�^y�6��e�۳�m��a�[Ը�q�
�I!Ke���p~{�\��m.�a5�u	��#��|�3�e��V�����o�;$��Rc^�;n����F�_�;���f�ޞ��*P'���w��7�|�?�S+u�䛆X@6G�;�u��@����$����Gܷ�xR| �O�c�Q�}���?�)�u��=���ro�����Ը�tŉ�ot��\������Q���ޅr]h��UBLy�g�|n��bd�ή,ӻ�qq�      ��ϭO�U�^"~#��(������k�����d���ŗƠ���N��x\L����Yj�W�>��L�E��/�ݚp�����y�}�Lȓ�]�vk�Z�t5�*,�|a��u�v����(��.�Bg�D�����~�L.ʯq��ƽ.G�qt��:�G{j��6���|?N���|�m��v#*��8��G���B���s�g��iţ$_��{`��i�3Ը?�(���䡞��ݥ&�H�lU��+$_�EΞ]��~k>f/�\���wF��Be�w�x�g�kwgJ�7zn�tȉţ%_��	�t}��FO}��I�c$_��iQs����>�c_㟪�3���au�5]>�     2�%�.+��{'���1(��Sm�nY�wSξ~�
�z��U{��yG����Snw����W�
�У_�_޽M�2�4)2��t#������~�iR�ˏ��r3&n�߰�{�v���Ì��R�ߐ�1�?���ߖW��U�zq;��r;��e�/?�ץ�n/d����{��s��R�'�^�;aq;��r��5�K�??���u�G��_�k��O��JG���k���ϵ�}E�Wٷ'B��w�k�)�^�}����G�sm�/?�}Ӷ^U�T�^��0�_,��逇�W��������{=��=�.˛��m��XP����]j�.��${��]�G�ׯY0\F�H>x.� ���      e�mzH�s�Y)-xM�ݽ�����\���f̲��˹G�1�AM�ݽ�����/�"3tIꡞ�ёǋ׭�k�-���3�괳�)u�xݫ}{�C�B���!�y��W^��췫�O�|�kU�����z�$�P���R����S��O�A�z�Yj��k�����Rً���n�u^�ތ�7|z�I깣x�^��55�x������L>d����z(�>�}�v�L�ɞ�^����u�Bg������*{����"��j�Y�"d���:����~��<�}،�7���g��ξI�"��Ԝ����͵�.Y�#^����~��~E�;�^�䥯￨��t��ε�h����(      C�^���=��%�����^�={�ݫs�=��^��hp��s�s(����`�<���Ц�#
���eG�W�v�S��]y1X*�-;J��Ve�do�x�./�ط[.(�$^U��=�}�<�����������^ӟ}��~�x��}`�x�./<l��ý�}c�׾1�kvF��^����UzeA�J���k�g�y���)�U{����޸ץ��T��{:��}#���볧�5���Sū�J�zp�7����Zy��i�Uz�����%��j�D���NWy8{�j��u�k������ǈW��w��d���9���x�&V/��GT��p�m���m�K���q`�|����^����m��      �{��rޑg�B*���mن�bZfN���ܵ?o���wԙR�{�o�r��ݹ��0�+X/����;����o���{�$$��s��6H��л�wm�����{wK�Q �N�����s�g�^e?���w���ߧ朸��wC��m��P���qߚy:����j�/��<8�u�/�[$��9������w3��m�ޮ���~E_�ʾH�]�q���K��j�^�Re?\]c�ǃ7�v��~���o��{7�v��޻ٯ���{/��DD���n�kt��BO�Īw:��9ӫٷH���`�������^�wxѯ�σ7��٫������/�K<xk���=�\��_j�b)�+GL�	�q��s�<�=     @&����Ws�������mK�{E�\�y����U���	���W���nz@���U4}�y�g�~9�d�x�.�.����7�5;��N)4|rJ�X�
;��͞}#:���Z)��i�^�|��p	 I����֧�N���߈�j	 ��@�}��i�ƉW��q߱���?��b���njꈇ՜�ٳ���z�չ�@��R���}��g��˞�I�ϧ�� ^�/�?���/�z'{]��Ke�|�R�S���e���=�{=��T��j�y��n(�V��9�׌��=o�@���e=*������g�Bp���tS��\�{�g�b���^��I����9z�{�K�=��^�Q�ۗ������P��x�&}�կ�x={     �L�k�r�`�9RZ8���vwӫ�ߺ���|$�w�[��Sϗ���������Ty�K4��K��l�����zt��T����;z[\�-t ��
����*��D�e ��_�d�);��v�MF��.���ҩ�{/�!�'�W��z�T��?�iy��}����|�޾�o�t'X�I�9��sm�d��.�x!{}��z�G���?�e_�{&���v�����{j�qD���D�Ξs.>UsG͜�7Pޝ%ߤ'�vy�����z���e�S�w��6p�vO�M��mP�g\./?���_*{}c����j�Y֕?�뛚�1{%w�g�iپ�      ��;�#���\}�'��)���ӵ/���:qW�C��]���{���G�������pɀ����~C:�������s���m�p����M���To�̨\:�h��Qe�`�N��)�Bg�,\:|�k��n��q���2�e.��"��`���Y��鐚�/q��Ռ�F�U��i��DL�(�"~Ý�o	w�sN���.)�Wz�;\Q>յ�o�t�����2�>����Ӥ���}>gTٿ��Ng߫�s���w眳]e��g��w�:��}���#W�c��F;�]�5��yp���t�z��j�4{ue7�钿��g�z��������]�<�;�[��kR�G�#�qm����{�ּX�`��q��?���w���]��C{%h���.ξ^��������&>     �Lypۓr���c+����)��_O�W�x�o��(�k/�^-+�ʻ�:s��Qnw���Y�q� ��J�i�u�GG/�������Lo���m�Z��$�c=d������\�}�2�x>g�j�q_A�Y��o����#�,[�k���Q��h��������yY]Xy��ϚP���q��_6�����5�}����m�wZ�G�T�z���:^����[��_�ʞh�|���m}���	�cj�_P*n�w2z�ow^g�!�&Mq��}Sz���ܙ���:���������\����������8�u��'q��/$�l�7F7�k�,.n��5�$O��ۻ�     ��tGc����]�����/f@����Yf����5wm��erʸ㥼��r���f��;������ �u��W�>�d\η�+�<ڳKZ!�wv��*��U��s��.}��[�}������?cظ�o��[e��P�^�9Ӈ-�tA���^y�g�ɾ����q�+���5�c���.��q��g�������N���������'�/���&;�]���|�/���rV�Dd�;�}����xH�ؾA�7|��=순g���GԹv�P�>џ���'�9�r�SV����g�9�j���c�\�����s�����ט�C$�?v�q�����g��[��X��=џ��e��Rwd���s�C#��U��${��#�;��u�]G<,�w�쏒w���]�t���4�zf��ND��΍r���V�>�;e���#�Z��v      _m�n�ۖG�'�r�G��_hX%n⪂{G�K��'������nJ�6o�p�s��!��-re�4�������<���VJ�����)��ZU�SebaYֿ���WP^?��ξE�?b�L,�~�}v����7���9G~���~���տt�Ϩ����ո��^�{5�Q��qog�~�����D̄]|Hf��U�����_*���Z�T�Q+!�v����9��<�߃���W�A���{je]_�}�=*�^�����{�vE���?�8�N��E9�*���eM�y�e�D�־������9�Z��nYz�?�ƽ^M_�99�^���{w˫}{��󇊘e���U�m��ڣ�Fd�{��Zzܿ��<䲷����~�T�R42�߃���`��
5�����_cN��9�^�{z�Yi��C-���9G��Ss0����)���qo��)����2�xTֿ���:�`�$Ԍ     ���˦����)��r�	'� ��H���n����6���ҸV��N.�Y������{�����H�^e���;�*䂲��R����}M����~cv�ҫ���c�L+i�|�����ӫ*�f���.��B��
޷ul ��+�޶oΙ��ҩ����^y%�d�!=T�գ�j��tw��>e�d�z����J���ǎ�d�z�?���|?-�d����v�t���;:���{ʎ��+2�5��4�`:Գ�;���A���W��v��F�U�f�S�`0T�����D�9�W��s�f���s�]�e�_S��������fEp�}C�P�wN�k�9��G����k�LRٟ�����/���k�      H]�2eѺ?ˌI��H$����\��r��1�ϩj�m�uߎ���	.�p���Y����(�N(�߾�DbC�M%�Oߔ�-�i?�Dg''��b�߱��WS��Wk#��j;���]���w�����2��N���P���/X�/;�w�+�!��%��s�ij�9�d���]
%��n�-���Ͼ���Ԓqr���[�k�9Ge�F��^��b���o.8]���՜S�s6�ژ:ת�~��q��>�ξ\N����12��q_��}De&����un�o���}����ƺ�k�-*��o�z���45ߟ��wp��;�F{�v��Ͽ�/Sُ�H�uр���0��/����kg_�sn�K�}���:G��C���Jf�w�:}��~��٫��W-'�7ۗ�=�S��Ώ�{��㾝����^�x��������-�5��Md�&�����%��~w<`�B�o��Wgo���k��"ǎ��~��~�     8�!�G����KN����K�r{a�s���;�������F�,�����ۗI�OK$��;7(���*�z��;�$�S�7���Q�V�)i�t����/��<=��]8��]n�c��C�E	�xLe?�ξ?�T���k#ݲK�O�o����RُJ/{=�ձj�g��CK�9�v��Q�eS�G��p蒊~<��׹OKc���Q٥�}��~{Te� �CѻH���F��}���3R�C��:y�ݮƽ�Y���.��xo�=�u�S
Gʄ�Ҵ�ߡƽ��ppz	�x�Ge_L�ٔ���@�L).�i��쟁.�:{}�M^�w�ל8�=��z�r,����u��=��C�;x�Ǔj���g���o'��o��9����ƬSϯ����s�!�<�A�}�3٫���s��D�V��f5���S��}����'��}���^�!�Cӻ�<�u&{+n?����_�t��!��S���g?%y}og?<���\��|=�������iu�=������7��y��w��s�~-S��.�     Ș'v� '�4MFE�2�u(��k����[���5[�Ηdzٹ�s�r��ݷ�!y�q� ��W��Z��1%2�?LF�K�P�s��/%�5U�}Ԍ�o��'��Q.M��>�����~��~�!����t����镦���b)R��f�����񰴙d�����6����C�75:��j�oӸ��u���b_�����+�%��Vyw�Bd����.�m�o���u���"÷/���}�v�j�w���bojt�����-ُ�w��.��1��؛"��O��w�טd�*����D?��-٫y�H�>S��=�ߜ}����������)���T�9��|�k`�)T��9��P?�bÿ_���=�_�!;
�9P��u����}���ϵd�{7�h����e�r�P�(��=�G��٧(���#`F�M�Ogo�Vfg� :{��X���[r��u����>5��J����>�����U���O��#�e�1�}�     d�-o,��8C$��.0���k4ˍ�,��_q+�ܵ�Vɸ�+䔂c?6���{�a�ܽ�d�~�)��.�����ϝ���W=Ev���UO��l#��!��!�ܱ�Xi٥uv���gqج���U�����M�#��>w�czuw�@v��^��     �*n&d��?��~I�h��cSn��h����u�{��.�k�\ƾ�S2��p옔�oc�V�Zu�X˚               ��bA�����I3��J��/�������q;�ܵ�;�}A����>������ �|�f�%�               ���+��}L>1�J1��J��/n���/�"[�w�x��W��v�|넯HQԟ�q(�^c�Y~��|�oE                ��ԳC,|V>Xq�X���1(�^�2�+�Ț���(�k�
�w[o���Z�����)�^CO�����KW�G               �t�n�(~���*.�J��O����K�Ƶ�%�)�kq3!7�q�T�Y/;�ϣ�>x;:�d�s7I���              ����K_",w����+�Sn�H"*�z�Y롕ۓ<Up��J���)_<��2E&�ez��탧�oV�H(               �I��JO�W���Q1��C�����'�+�xa�li�!^乂{ҟv�C>|�t9��$I$<�)�ޓ�^�[��YfB               �L���;�9�~^$r���)�^s�U~�|�4�ū<[p��Z�Nh��7]�}�7�;��7����*l{J               �L��W[�ʜ?/���7�;�탷j�:�^u��A�2Oܵ�{�Im`��>���ۿG�}p��:�+j���               dK,��m�M>2�29��D����)a�r����M�i��u�/�k-}���ʌ�?-�V/'N��ke��?J0�'               @.,�}R�]+�����)��~��q��(�k13.7�)g�?I����6Jpp�N�e����xT,�                �6wl�y��j���c.�0�r�:Y��v	D��O�����e��y|�|�����.d`���zY����Y'               �[D1�Ys�<_�R*���U>Q�f�X�������]���B�yWp�z�A�e����q��8�32q�8�H(�e��C۟�b�v               �Ӧ�mr�?�O��a��_&���=�.�?߰R��ڽ��|��?������}�|�ԏȰ���`~������IW83               �G$�;��M����|�{'�#CՎ�:�mݽ��u�仼.�k	3!l{J^hxU>y���i�;8�6o�?o��=�               �i�m�߾\#���.�?�*���/����W�i�2��wg�[j��%��|������;����Z6�=�)�۶               �u��l�o?�K9����'}X�=U�Us�U���ay��%I�b{R�6����]��'{U���>��;�KyQ��}W���rߖ�ek�N               �ͪ=�ۏ��'<n��稳�g�vt�Ƀ۞���_r���!WpO�
��+�����������.���xs���`�<��y��iu	               ��6�m�cK+���-W�>��h�P<,�կ�g�V���n�ܓ���p��2�(�p�䂣ϕ�e���Ѡ�h\#ϫ���u��z;               0Դ�u�߶<"��xL�9��`�9r�QgJi�0q���5M�兆WeU�:	�#�~C�྿��F����y�?�؊)r������i�ض�1�,k�7������e�$̄                IX��nZo?
��YNw��>s�r������3�-k�6Ț���^�����A�謳������Ic�����ı��1���"aF������I��m������Z��               ��b�ؾ"�6�t��<�r�z�0�X�<�)�e�JmZ�4��;�.���;�,��}���e��쇦Ws?b��:r�L1Q&����ecd��2��\���q��/NO�W�C����&{{ۤQ���F���                ��־vy�^?^�����ˤ�2yđrd�_:��W����./.~�w���z �@�W��=Ң��7�f?t��g����QpO����1�l?��_hl��{����g-a%$�H�LHo4h                �fB�������aRRPd���0M	������X�=C(�g��Ҡ#�%                �I��5��5���;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;                �(�                \��;r+!��L               rϪ��� g(�#�
��b>�-               �=��
IL�	�+�                �@�                �
ܑ[�!>�X                ���++-��.<C               �{��m�^��+�                �@�                �
ܑSQ#&�w�               �^�Ę �D�93���&EEE�H$�               ������5�I ^��b"�
Z-?~��5J,˒��:�F�              ��+--�I�&����H��G�>r��;r�x�)S����v�0{%w
�               �QRR��c�h�4�4Y=>��;r��;rB�ۧv��ܮ��a	�              ���������b��W�I(�#7(�#�t�}Z�89j��������,K               ��x\���e���RXXh��.�-��nJ��:
�Ȫ}�����              �@��u�s����q�DZ��;���;��r;              �;Qr�[PpGVPn              p7J�p
��8��               �@��F�E�              �[(�#�(�#c(�              x%w�
wd�v               o��\���Qn              ��ܑm��(��               ���;���;S��r;              @>:d����1� N��G�����               ��%��z%wJ�pw��r;              ��@��F�i��              0�PrG&QpG�(�              M�ܑ)ܑ��               C%wdw�v               h���4
���               �%w8��;�v               %w8��;�v               
%w8��;��v               J�Hw�v               %w���;�r;               Rq����bH�tSr�AQp�Qn              @:Tr;v�H�Pr�AQpb
�G�����#+Fʔ�S���ΎzI������              ��C��[Z:�@�޴�������MҺ�u�?�(�ةł����PH�����KLYR��;,�>�r;               q��{�1"�`\F��.k[��M]W�)Z(��?$'�r;               �u��{AA�����(��?ttt����4����r;               Җ,��7N���7-�h������,               ��tɽ��I����                p
�                 W��                p
�                 W��                p
�                 W��                p
�                 W��                p
�                 W��                p
��)�eٿ             �C��|b��+ o���X4��H$v�              �.���~)**�� �N���%�P($}}}��             �t7/�����+����III�]~���D"(�             �A����z�`P�n��w���a������               ;tѽ��G�Ѩ�����;����{�m�L<�V�)ɧ �=�������0��cw�ؽً�Fw'�c�:-���v�,D~��G)S�K�P�*ԯ��Ñ���իWQUU          �w{{u]ǳgϢ,� �G�G���Jq{Z        ��I-_j�>��3����pD�&�v         �Cj�R����� �C�Gr}}��"         �|��󸺺���� O�G�4M��         �I��l6��h�a	��^�~]�         ����=}�4���Á�u�_�         �Wj���1�L�v{{         @�R�wyy�����Lo        �� p�����K��         �ߪ��F�����          NG]�w8 �;���         pZR�>�N8�;P�u         �����"         �E��%p           w           � p           w8QEQ�t:��h��         ���i���:��y�6pZ�pb.//��ӧ��ѣ(�2         �_j�6^�~?��C\]]p�p"��������-         �ii��'O����&����ț�N��g��ŋQE          �I�e��ķ�~�}�] ��C���~         ����~���d��/_�'�;d,Mn�        ��|���QUU�z�*���!S��8�?         �~�x�"�����}�4�8�;�&���2(         �~��/uz_�u y���F�A����ɓ'         ܍Ǐ�x<���?������;��E.-�.i         w'uz�=�W�^}r����;h2��b�u��o6�         p���zw8,�qp@)nO]UU���b         w/��������GE���Z�[        �����Lx�K������h�����u         �����ڲ,c:�pXw8�t����y�̺	�         ��>��]\\���������2noo�i����?�_~�e          w'�z2���8<�;�ӧO�/���n�X�|>wi         �#��Kۇ<y�$���Ñ���?~�ѳ�������         ���|���Oq{j�����Gt~~m�����/�.�/��)�         ��������G��l6�x�pd���QE�w]����ӟ�ԟ�Bx         `w��<���럽/u|)n����	�!1�L�~�'�������?�W_}�0         ����m���Y�7��ɓ'}���2���?����~ss��4����w��]<�<�={֟%         �����>^�|�S��z�4�6m�<ȇ�2��%N�Ybik��_L���?���_|џ)         ��׿�5����X,��ib�l6�[��,ȋ�2�����~Kܫ��o�%Q��c�}�]���m<��;{        ��.�M�eSw��������O���Ǐc2����/ߡ����~l1M�p�         ��;;;�7��          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,܁�k�6���ٖ�        ��*���i+���I�ܩ�����        ��Z�)xO�h4�wJ��U:�i�����-         �k��,mUU�4�]���;��UԾ
�        ���m�V��x<�{!p��PR�^׵�        �K=Y
�Ӗ���bw�m܁���=�         ������bѿ�B��d ����3�R؞6         Xg՜	݁M܁OZ��M���        �&���&��G��}u�         ��j�j��G�Q |�����m������5���m�>W����_         ܙiE���Ho���F���KS���eه���]w�gR؞Β۷��muS/P���ٻ          #)z�)|Ũ��{Y�/FOX��y���~+
#Q�7�@/,���=��~�6]N���I���O�        `��o�RM�Fl�|��~�z
�ǣ�>z�G����~�4w`E�D�4���}��iB{�T�m         �)DO/�KS��帏�ǣ�r��4���i���� <pij{
�w�um,�y�mݿ        �=�uo��VQe�˳��w������c:<p���@�����2��m���ET�"b���         ��4�jnc��&��8�L�,�����Ե��������������51��Ѵu         ��nQ-�q9��d��D�U�"�]&��I��.q{:+nQ��S�        �CR�޴U\ϫ����}�i�WK��t:��#p�$]�e��.N��:��M)         "MtO��l2��x��ǧ��$wxX��@�uUUm�q)h�]�D��q���y]�]�        ��+R(vǟ����:��$f�󍦹�&���}4p�	��H�۷�ۛ��*�z�����(�����;V;��        ��ū?%c�/w�VJĚ����&f���7KXW���?�;�s)nO�h�D:�mQϣZn{Q��R̞��U�>�<         �ܪ�z/�J�{�o�����q[]Ť����l�4��k[,b6�m48=w��V�&�ny𰸎�mv���)l_qX        pZ�����_}�^D���W�mߩͦ����<�ө��1�;�Sm�n�/n��u���x5��         �U���/��b��MW��m�ˍ&����~��=���ۡ��ϯ���u[XE�         �X1ꢟ���V�YM\߾���E�F�a�u� �������	�C�q�b˸��v        �mՏ�3Y��?����z>���F.�r����p�4M�/�C�M�}ܾ��xs��rˉ�         �+}S��Զ觬o4s��6�ܫ�Z~�b���i��=��HK�]���mu��'Jq{
ۋ         ��+�(�/]�E侸���e�e9�CR��-
A�w�G�B=TץK�\��&�pE�<vܐ�7go���������M�        ؏7]�f�y��u\�_��S��N�� ��;�u]�܇H��⪏�Kg��S�O+ O�Ĵm����C������         �e�"�k��������A��S;���X���d�R���n����fq{Qv'�~���ti��Mi��         �������������p�N�{���7a� �jMS��"N"n�x���/I        �q��m�T�$E��"����oj�&�I �M�'.���4͠}�f��׷��<Dd��QS���         d.��D���<F�Q�����>���<	�ᄥE>��6t�yu����<��>l�S�nZ;        ���4@�������A����t����	K����{��w];�W��3#l        xx���y�f����m�oe�3�S%p��.�2h�����o�ۋ�gv���Yn�h�G         ��TU��$F�Ѡ}Mq��%p������onq{:�U�/���        ������������M�'*�a6Ģ�G�*�!��+n��~        �4v5�}S��t	���u=hz{�gQ���b���+����V��         �H�[Q����������	�)��r	〡�p�Ң;D��>T�ɕX�&Mn/��        ��aHܞ�>Mg?;;[���N��NL:�,m��x�v�e�~�����~        ��Y,1�L�F�)p:ȇ�N����}���֗w�C�^�5"         ��M����rY8%�c����|�~E���#�],��V�        �0�Lq��i�'�m��̳u�z���������j���         ���!�z���V�e �A�'���a�5ՠ��>��E'n        `UU�ΞBx�;��;���Ȯ�vm4��>�m/������v         ���ƦI�Ś.MpN��N��v���G��)n?��x         r6$\O�����O�������Nľ�8�:���$         �qCc�4�}]���o4�?�;���i���u�r^�_��r���к���G        ���ں!���p:�p"�Lp��z؝#n_@tq;         ��"��x�v��d@��p���o�0��8������        ��	��!�&��'p�04poځ��[~Y݀�         6UUUL�ӵ��o42�r'p���[�O�okzz{��2         `SC����>���O�'`��f����L���r9         ��.Z_i�&��Og����8.�;��!g��]��������o6         �CC�u��4�!s�K��3�̲�-�]z1�        ���n�$��uv��	�!sC��n�{��\��        �ݬ�ۓ���'A���g6���        ��!܇Ngr_�q	�!sC�~��jM~3L�          ��&+p��	܁�3�        �C��� p�{aؙg��5˃��         ���p}�w�x!�i;t�=Dwވ�        ؟�q�	�p?��!I�]������         ��2P�wȟ��L&��M          �����4.�         ����^tm�C�         ����~�          ;��і          ��{љ�         �������          ��ؙ�         �}���          �]	܁�u          ;��3�         �=�;��w          �B����v          �D��X��         �>܁�t�v          �D��/܋          �]	܁��         ��܁���;          � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p8q��(&�I@Ҷm,�����Lz�@R�u��3�N�(��$��I?s>%=^��V��yt]��}ʲ�����$=^��f��x�o�4MUU��/��I?s I����Yg6��9&vl��noo����>���>���>���>���>6��>���>�1��> ��h�ĥ_Z��{V���+=f���d�_x��:�J��!1�5�w�5j�/�<nxא_x9&�}C~�3~��J:�Y����Yû�����}�1��ر��|��|��|�c�7��>�6���}lc����c'�2��> ��h          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�          Ȃ�          �,�����:���&�o�h�qܴ��(�2          ��ڮ�y����]�g��=/o�QM�F��M����Yn�G��7���g�f1�j���}D�          ܙ����U������On�+��3.�;�v��ݳ�g�?����4q�u          �o��Z��?�ў���V��B;���o�X������DQ          쬝D\�KՋ2�C�|T�����v������4w          ��\D\�۸�����I�e?��(��F�         �Vڋ"^��(�i�'	�Y+� ��_�x�ߛ(�          ���I���3���A�$��.���l          ����Q4�����2��8���         ������E0����\�cg^��q         ��2��ˀM��Hw^���2��W�         �q���hg����;������          >j�����9�;k��<��          ���q�o�)�;[�>/b��          x_�������J�Y�&          �}�3�;�����2          ����lK��V�i          �uS�َ���tc?t          ��n��;�ѷ          {&p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p           w           � p     �?{w�"�u�a���O�-am��I���&��%[aG�q ��5��U��	e2]U��u]�0�Z�N�u�     � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "��r�ݮ�i*h殅�fS}�4�8κ����ƜuӮ�n�7�9eݰF��}���7w-�=q�u�0�i�1�(�͹�X7�iΞؼ�}�}�1go�xF��ކ5�<��=ɺa)�>�-y�i�Ǎ�{b r	��r�˜/�,վ��B�R��`��rúa){ְ�a������a){ְnXÞ�5�mXʼ�5�mX�ކ5�� ��E�          @�;           �           D�          A�          @�;           �           D�������c�s�m���v�kk��h�a��rrrR]�4�^��9wi륭���nk��;���a_[/m�rttt��f��ƞ�}s�6���i��9��ކ7m6���X7�3�c�>�0�c�9�>s�����yk̝��˄�-׾�y�΍�/�� �P�m�8g(tvvVp��o��<�Q�kϨ9��uþ9/�ڞ�vn�{͜�M��x�žC�i�y<��7�^c��9�y���Xü�5����mx�yk�����y_���������\w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�         x'L�T@6�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D�          A�          @�;           �           D���T           ?*�;�t;�;          �놪I��
��tW          �ꮦ���`)�;��,          �UkM��	�Y��c         �m��M���	�,'pg���O          �9֚����Ŏ����m          ����t��;ŝe�,v��_�          p��'c���Q�w�/�u��j,          ���WS]~4�x�w���Ƚ�C��         �Cƪ��N��S�;�	ܙ�����          s�<��Q��Q_0���Y�S]|1          ,�ޟ���~W�{Nr�0�;��S���Xݮ          `�n[�-����5��ܹ���;�����=          �ѿ����z�Y�$w�$p�:�f��/'�         �k���χz�I_�G}�m����r�{��k��         ���U��i�͇S������i��'�;��������������         ��D;���ۡv�:��_^�/k,�3#p'uWSuߏ�}��ý����?�����׏k#n         �'֍UO�������r��骞�xZ�Ϫ~qR�}M�Nx���1'����ɫ��o\�����w��m�ق� �:���;�N:��{�﹀��ۘڻR������X�xF2ǉE������(�N ������/�z          pW���Gq�?�"�>뿖i��?Nc�O��C�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @� n�\�|>H]��o�XD۶)G��Xû�<��>~oxאu���zn3t-�az����UU�!�#��d��]C�)�7�o����x���؆���Ɛ��6�Ϲ��|������}�x8|w��'�N�ٔ'��t:�D>Q���M������Me̓lb6�l�Ŧ�۰������k��|�pN�6<��6<� ���          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"ܡp]׭ߩ�,�         x��JD��C�v���ʺ��        ����~�C�,��]NpwB         @��v"x(���.          �O���m��        �͘����
7x�ͭ��/����Z        ����!p��]t몎�[�;Z\M\ߡj��        ��u=h?!<�O���7�ƚ���}�~5=�V         �u�ږ�i�A��C��P�\Ls�����g���J�]�Ϸ0         Ґ(}�>C��wK�`P�^���ƬWy\W�        p7�Lp7���@^5ֶ��4�,���z�λ^;=         nǐ��&��a����*u�u��!|ty��Nr����l        `�2\������� �j���X.�ػ~��V         ��u]7(Jo�f��Lp�� p�0tQ5�X.���t����j��t�,         vb����h}��2���DF�m{�t�Q=�鐃u�Hw�K�ww         �l�w���p��@��.p���r��֔��n��^�?۰�y        ��t]7h�z�uC�����Á����q����Ի�j����'��q        `F�a)�)�@�p �����k��u��k��v��p         p�!S��x<t�����H^A�\^?����h�Q,�����?9m}��{sy�E�         ܪ��>$\7���H.����4㵁{�)�Y���´�򭫻��+�         �]C���l���/H]���f]w����h��ED�~�z���G��.:�;         �([�!��W�p8�p`rA^,�Og���b6�X�_�UQe��)���?����         p&�ɠp}H�E�fh�>O�Oq��~߷���Q1�         v-��܇����ÁɗKɭm��^]���I�3r_���	        P�M��j��_�}���F1����7�|9[?�=�b�j��5�lMq        `������x<tL���0	�� ��*�ք��˰��b6�X��Cu��E�y�nyy���o         \o����>d����p��p��
��S��y��r�A�7��w4x�w�N�         �\��1Id�P��5t�{����b~�����ݛm]z�i#�;*�        x�����W�u��I�,�0�����kF1Z�c�\?��j�{u��wQ� r��m�5�        �����;���p����Ex�\F۶k����b�.�����Oz_��!�q�L�        ��r{�C��e�Á��1�N��WWuON����*`�[FT;X�/�:�Q��/         ]�uQUÇ��?�:�	�����6�I��4u��Q����]���FT7�^����n��	        �=�M�>t"�h4�:�	���+Ά�)�e���>��˓����a��˟q�'7=         �h��=����󸦷�� p�{`�0��â���q\t�h�v�t]t�W]T7���?1�\k&p        ��rj{No*cx�~���D.�9�}H�^Wu�L���,�"������i�[��q����         �w]�m4�=��'''�oW׵���p�L&�����o�G�q>=��ׇj����D�[b�����8s��        �m�������������;�#��z6�ڿ��~���٫~:�`]ݛ��W��檦�̋�I�         ��6S��jr{Ndj<ou_@��p�4Mӿ��b������Q\��7���f�nyyR��[�ԣ<L��        �^�iܞ�P�o�?p�p�ݶm�1jFqR]E���ۼ�]E��o�W�(Tu��]A        p�Va��q����F��s��?��រL&1�N���!r����Q������{�t���I�         ���I�ۄ�)C���7�}p?	������(...6�M'��o"��vw�&t����ݫ|����nV��c�        ثm��w5M'''��������2	��[]�6��Or�_���qL���n���۩���3]t�U����d�F,���        p�ޟ־ٶe��)q;�w���
�4��6����8�j��<;��qy��!��yE����{;��r~0n��w�:         ؏�C�����X9�}նmr��x,n�@�@���n�F�f���q1{�v�����}���&x���/ߏr�{o��        �c�F���㻎�G�Qou܌�7���$p�b������d������Q,���.^G׶��Cv����&ku��y�yk�;        ���c"z�G���os�l��ZC�����k�NrO9ͽi�l~������Uy^R��-���-         7�q���эn/n��E�LF�y%�t:�h�{�.ߎ�'1Mb6��b�y(U�^u���        �d��۷�or;<\wx�VNrﶘ�^WMON.o{��t���s�;        @��M�m۰=e�~�c �K�T� ��q��<���VǨ����>]��v]��>�>t���s"        p2Dω��G�Q,������䞁{��ݖS�W�������"�<�[��?^�*t�"��Ƚ��        �[�!znM���xٳ��X����	ANt�N�[G�k�o�8�c�e��2ڮ��n�<����7�{����M�n�;        �Meg�ֳ9���<n���@��r����Q?�='���x�o�f�o)�������{w��������[��Jw���t�0�        `�l�V�S�}n��]�G�����x+O�%^2F��f;����f�Nt~��d�|����O�/?����w�F�U��v�e�;        �pd����6��|�����4��䞡�m�OS5        ���K���� F�|P�@����|>��b         ��U�~����&p�ʓ��2r��         ��F}�0��,O2r�        p��Ҟ���������V��r�|�        @]�o�v�m܁��	��$$��g�޶m         �pdԾ��LknJ���j�{�uoC���s         �WQ{���$pv*OT2t_y7xϏW         �a����p[���z?xO����	���"x        �ە}Wn�k�>^}}�����ػ�I���          x��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�          (��          �"�ဴm]���      `�� �CTU�s8 w(T����<f�Y�-�          6���h4�������I��ɰ����q~~nR;         ��j�ln��5M'''���;P�;d:�Ư��*l        �[�\.�իW�0�'O����Q e�C�ʰ\(�0         `?r �˗/�I�?6�
 p�;�q��/��=         �/�f���GE]���;ܡ��+���b         ��ɖ/���?��$w�Cw�C���         
�M�˗/�I�����9??��l         @9�������4����X.�qvv         @y��;::��i�/�;܁W�^E�u         �'�l��={�~	�a��EL��          ʕ��r�4��L�{vqq         @���{��Q �#p�=3�         ���O�{�/U�         P�U��4M �!p�=���         �l��?w�#��        �h�`��G]�         p8��_w�#�         ���          �"�          (��          �"��@UU��$��q4M�         Y�u�\.c�X�t:�?�����i|��G��ѣ>l         ��m�x��U�|�2���8w8�����g���;         p�����ӧ�v~~ϟ?���� �&p�����UU         ��.���3�����駟(��
�׿���         �����>������?P&�;죏>�        �e��X,�ŋ�G���F�駟         �[9����,����}s�;�?wأM��ۛ�	         `���;���.���a�rA��ӧO         �O�<��.��k�3��K�{4���E�K�         ���N/{�/^\����K�{4��w||         ��:::Z������;�Q^�5�Lb6�]���I�         ����[��l���Q���^�w�!         ܾu����q �%p�=�����,ڶ��>��"         ��5��?���i����~	�a��j����x�����n�         v�^���d�w`��p2p������_�5>���          nO�zf4��;�w�#O�<����O�7��b:�zi         �%����������S����ᎌ��>r���_ϟ?����*         ������������w�n��;�/_Ҷm�����{����s�         v�իW���l�����;w�c�=��������}����wX��         ��M���������O��ۡ w(@�����/�\.�~=����7��_��        ��^�~�~�m��4MϞ=�;>���K�B�����O�����V��3x�����>��?�8��
         `�l�~���������y�㝞���6�!p�����ѣ~Z{^%vqq�v������ŋ����R         X�_~��1��i�yNj?::�[���(��
�f��e�>����������O?�kn����Y         ��Ξ��b��̞���_o�&�<y�ɤ�(��
�i��f�         �7��ٳg�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;           E�          P�;PUU|���1��~����          ��z��i|��'q~~ϟ?x���?8==�Ǐ�������"          ��gϞ��������d/^�����%p���i�mu]�������         �ڻq{���X,�i��w	��'M�'���~��ˋ_�~:�8b1_ƿ����ꫯ�F�_~�e����          �~ܞa�7�|�����w-봞��u����"p`��g��?�����������[�V��E�          �gq{b�忖q�sz{?�۲�W������Y_>X��         ���q����9�;$r         `�v�%p�Z"w          6!n�&�%r         `q;7%pg�;          ���w[E���|_~���         ����]������Y��         ���[w6&r          =}�T��N	�ي�         �a˸��������������         �����r)ng'�܈�         �a�s��ܘ�         �a�P���?�vvB��N��         �7q;� pgg2r���E���#�/��������         ��#ng_������c=���E�UU���.r         8,�v�I�����W?��         �Љ��7�;�B�     ��o����*����m��%!��}a�����!�x	ۉ}�'�=�N&��so<���8��x��1ccC �`��KX$��RkCKkW/����c�Iݒ��T���s��U:oש���{~   7q;� p��tE[ra��         �8��)�;�*���P��         �(��)$�;�N�         P�������         ����4��7"w         �t��w�J�         �.�v�D�N�)r߼ys477          �oРA�vRE�NA�v�^WW�ܓ#�H�         �C���������I"���"�7ǘ1c���2<          �ǁ������[�l�}������j���ͱ~�����l6          ȏ�{��"�����쌶�ʀB�SP��1xpM          Px���P(w
�_g��<yr          Px�:WE���P�           ���          �T�SP---�x��          ����y���"p��:::b��}         @�e�C
I�          @*�          H�;�Y�	          
/;�2���Tgu&:&؆          ��          ���          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�          H��q1`X�0"F����cp߁1�Or�DUeU����{������f�@[c�?t0�6Ʈ�=��iWlol���ۑ�          �w������o��'��뀓&�oU�w�����ƶ�8��[�@���ݼ/��hl���I̱�wS&��1GŬSc�Ic��1qh]�?�iO��l{l޿-6����n�����=s?          �M��1%��49&��IC�ň'��u���{7����c�����aM�m�t����{��9qƨ�1g���g`��YUQ����	���Y[�=V�^�m[�-�u{7Fggg           �oe��;rF�9zn�6jV�8:7����7$��g^�˶Ɲ����`ےx}��hnk	ޝ��mN82�7?.�;+��AuEU�1-w|b�swu����xv�˱b���vf          �]��~q֘��q�s�y�����=�6��|Qtd;bю����W�-�`kc��x�
�u��h��q��b�I�"풻:��zI��ռ7���\<������          PN���� �+'_�=3�TVG�UVT�������xy�xt�ӹ	�_�y�>v����i��E��ݭQ���7��@\?��XtxS����b������          P��U��K'��zi�.FUUqnݙ�cG���'㑵OGc[S����g�������)Q���R�<��G���o�V=Onx!:��         @	�wPn��US����D�Y3<n9���q�����+�]�{�ܔU�>aH]|d�����Q���n��⣳�����y<��Y�;          E�u��f�%q�̫c@u�(U��n��q������Ǐ��K�i��,���㓧���͋L&�"����y7�5S/��-�'^߱<          ��TVT����ξ6����������&_�N��Mto�h�RWҁ{���a�5�W�.W�����}_�ݺ0�XxOlol          H�3FωϜ��;ht��~U}���|0��tA�����7���d�9���y7��f~��ǜ����,{0~����          H�dR�ͧ�^n�9o�0<�ù���(�񵻢�iw���ܓ;>}�G��IF&�	�*�d���~nݼ��Kߍ-�          �Źugƭg~"�����O��_5=�XxO<���(5%�O6!�x�gc̠Q��%�����Sܷ����G��4w          
(�|˩�ǵS/��U����O���ķ�0���RQ2��u�.�O�zCTVTG��fc���1�sRL?������Es{K          @��<&���[c��A�444D�=1�⟷<KVE)(�����*n�ws\:�{��}ժU��ؘ��r_g�������ڽ          ���1�ǟ��1���=Iܾq����쌦���%C��=k�bWԁ��~��K|>&t����.�����c~/�\<���          �ޔ�d��7n�����t�Ν;sq�okmm���s?������F�*��}T͈��}!�t�{��]��ĥΊ�)���          ������y���~'�dr��M���ϒV���o���[�k+���e�>i����Yn�;�s����7-3.�x���W�          p"���y���)#gݗ�����G}\gcG��S?�XwW�l�Ŧ��9�����\��tOw��.���Q�:$�l����ߙ�          �W� ������S��K���7v���-m�I7�w7���E1)��}�ɧƟ��ǹ�$�{z���A-���>_[�}�;          �%��������2lB�}ݝ��v����o�o��$�4m�bQ4���#gƟ�wkTWͯ\p��w�i�:��$w          8UU�X��3=���vm����?��-��E-�|�_��9q{������C���������{          z�"S_8���Q���;���o����N�X���ES{K�]���k�/ο-�U���D��]F��7N�:�]��          �����?�����x'��]gk6�8���_�'�;;"�R��S_���1���{z#nOtvvƜ�ɱe������          ���s>�N�,�5���2-���Y��ۗ}/�,��{E&����ƘA���魸�KGGG\;�}QpKl9�=          �\8�����k��;ѓ�߮�P�������FZ�6p�����s����KsSs�6���E߈C�          o7qH]���[����;;;{m��ܳ�'�i#f���#�R��[wf|p�A��+n�Ҳ�)>7����;          ~[��~�������ݓ���K[[[�0��X�ch�O��܇��ͻ%2�Lpt��ۻn���?/���|          @�?:�8y�Ƞ{�����>�k�6�?�������3/Q}O�*p��T�����ԧ&8�B�퉓O>9>3�c�d���Ѹ+          �ܱg��~'螮���6`���>yz\s�xx��&�
ܯ�rI�:rfpt���Ǎ#G�yW͟�����nOݝ          ���~������������ӧGeee|��b��e����H�����Ms?]Z�����q�������          ��g|<��	�.q{���:7��/~��"ۙ�4HM�~�OD��~���)n��So�W�X{[�          ���1���u�KK��e���q��㑵OE�"p?{��q�����1nO$w�$�����         ��RUQ�:�#�ѥ-n�r����^����߮��{nC�zCpdi�ۻ\6���]k��          ��w�_c��,�q{b`������~�V������ĘA������=Q���O�zC��S�          �ap�Aq�k�#Ks������/�<[l�B*h�ޯ�o\?���{+����)#gƩ��E;V          �/i��W��[1��ʊ��؜����)
������.�!}ﮘ��.7��p,z��          J۰~C��S.�[���]ί�?��ذwsJ��dz��_��b��3�O��G͎�ۗ          ���f�?�V�	�]��퉊LE�8�����R������Ǡ>5�;k���Cӯ�         ���U���I���.玝�kjc[��(���I��˂w*��=q��91i�X�wS          Pz��zI.r睊9nOTd2q������P��}��s���R��R�ۻ$oZ�|�         @iI諧\�S���].�x^���Es{K�[A�+&]�U)��Ɲ�[���lj          z���ƈ'oU*q{"������uOG��=p�h�?���7
��?>jkkO�y�M}�����u�          ���IoUȸ}ڴi'4n�r���#p�x¹��%�M��w�d�yw         �2����?��7
�WU�N>u؄�0dl���������qgo*�=1s���0<v6�
          �߹��Ee�"xS���]�7����5�1i踠���D&�������          ���u�7�zܞ����ђ"����7ΆN�C��圱��         J��>51�vfPq{b̠Q1~�ظk�K^�y�O�rWNq{b��7����          �8����L��r�ۻ�9zni�������S���[ܞH��N93���j          P�捞����ę'���z4o����R;#*+*�\�c��%�[G�         Pܒ&���cܞ�=bj����֎�����g9s��(W��'f��          �Q5#��C�\�kܞ������&Ʋ���Y/�d�)Q��=nO����ā��_          �߬�;캜��.�k��V�^���U��F���L&ӇO�W�X          ��'M�r$nӌ<��yy�u�O�>��QN��o5aH��         �HM:.ʍ��7�����Y'qs9)d�>nܸ��퉉C�          �'����!c�����jĀ�b`��8���}t�����92�h��;         @1�X�T�r!nw���e�{}��<�Q5�(����m��=�ܽ����         8>c��r!no�֖R�><J�����U���}žC�         ��1�Z�����FՌ��:y�
������3j��;         @��P�-pB�~t%�Wf*r��K������          ����v*n�|���~5��L&J���g�          �Rn@��ݗ�}���{��(E���ܷt��          J�����=���ׯʀ��Qj��Ǧ��         @��g@�q{���i�������R"n?v��         @q��(��H��Ǧ*���ׯNUeq� �F�~|J�f         �rPJ����%7:d2�^�v��gJcj����UW���;          堲�4z`q��I���Le�w���:�~�::;�؉�O��l��         �r�-�X�~bd;���F�����I�~�e{�n          N��"r,n?1�a�%��eۢX��O�֎��          媽����O��<u�~Ś�Z���O���C         @qi.�x׮]��(_��ׯځփQl��c�         �r��Ё(6I�^__/n?����������fq{���R|on          ��@k����!n��H�ޞm�ƶ���i'n�]�	�         ��ޖ�Q,��g_����fh�wq{��Ѵ+          (.;������;�N^�⎦��8�.�J���:���yO          P\�aȱ����h��>�˕�v0?��������ol�<�a          p��l�4��G�nt���ܸk���=6��          �7n��l{TW�/�����}��N^�h}��LO2n?~|���F9��         ���llڷ5&i"nϟ����yo^��S�%��7NE&i nϿ4��          @���ߒ��]ܞ_�8�:/W���-8O:.
M�^�v�          �Ӫ]��	�F���oŮ�y[+oWwyÚ�����hhڝ;          (N�w��4���Rܯ�zI���p��         ��ٸok4�5ǀ����텑\����m��]��;W�\&��|�֢�+         �����ҝ��1�d}q{�������zy��{[�����b��O���[�}i          P�^۶� �����^ݶ8����j'�s>wq{�mط9�v          �-	��M�^x�~��z�_ܲ ��yu^�����[_          ���Ɔ���C�򲞸���6Ɗ]k�f^�����c[��]ӻ�==���r          P���j^�B��5551}������|�;�y]3�<��^��.nO�-�E��-         @ix�����9��5����\�]�=pz�K��������/          �c[��X�{}L;iR��_ܞ���ƒ�+�n��d���]�b���'����t�����          J˯�?�+���=]_�ld��Z$��']��	�������bw��          ��<�����i��U�N�9��钼�v]����Û������<�s�����k�          JOs{K�z�q��KN�������ű�qgA�.H�~��5~����Ȭk��<��tڰos��}Y          P�X�h���Q���y���t��G�vA��ë�~U���>��/nO��W>��7          �g{cC��eA�[w�1�CܞNk��ǒ�+�~��}��ǯ�?�zi����=�v4�g7�          ���V�<~g��9�)�����w��]�`�{��?��']}+�t������D{�=          (mɤ.�E�=!nO��״�
��i��\�d|p���z��=ݶ�Om>�X�  xIDAT|1          (?^�/q��Ӣ"ӽh\ܞn?Z�@�_��+h���w��㒉���>��8q{�ݹ��xC         �?�m�'6<�O�ਏ��ۢ���7��(|�~��1�^�@�љ7��c���hǊ�׭�          �凋��͋����1���ӦM�E2��{iP��=�躧��S��Խ�����ב��.�;          (?�폟,{(>uڍ���������_��A*���l|�;�]��Q���������+~�o          �Ӄ��ǟS�Mx����鷧e_�h�����wo���<�M�<����8l=�=�]�p          P����_��q�e�)*+*s?��|�hlk��HM���k��1o�)1��V�^���l�7��l{          P�6��?]���Ȭk��E��/�K[D��*poi?���Oq뤏�=n�d21a>|x�=?Y�P,oX          ����c��IѾ�%�k'q�ԩS����д;����H�T{����U11F�u�q�Ɖ�{`�uqﲇ          �d;����_�rK�4�/r7��g:�N�������%���^}���?����|$A2�}ĈA��;�?���?�66          ������P��qՠs������3���~�觱�au�Q*�������ߏ�8����ګk��{&{����KwDCӞ          �w�¶���a3bdǐ^]�+n�����-�տ��Je��hlm���>qud{�΍L&�Ǐ������/          8�﮸'�jέ���;S���=�a�������H�V��+�������<��_Dq{�=���xh��          G�љ������M��hoi;��������_��z4��D��:pO<����礘[=儜���c�|���          �][��ό�>���O�9��=���_~���iw�]����6�*M��	���\���[�cy��߉l�?�          �t�t���Ѷ���#wq{ϵv��y��~�(E�'~����m��cxǐc��&�����W��f�eO�3          ������Ϫ��4:�;�����k�h��<��X�sU��	��Z}w��bLg�#uq{�-kX_~����P          ��X�kytd;���+z���{���%��ߎ�ۖF1)��=q���⦉��䊱�z�����mK�>���G          ���xϪhjo���\m݋���=��e|����{��]���kÃq�؋���#�������u���W~���          �i큍����I���ܫ��{n{cC��O-�8�#�QQoy2v���(�Z�9e�������{�?�,{0�5          �-��k�/��tDӻ���܆}��o����ݼ7�U�v��Z�3o���Co��q�Ɖ�{���9��ʝ���W          z[c[s|eٷ�Of"���D6���]��s�l���֫?�涖(fE�'�l�//�V|~�'�Sun�x2����6螵{��o_�N�~          ũ#����θj�Eq��3�P�!q{�e����W?����DkG[|u�w��)&\�#�����'���7t��k          ���Ƨc������c�xq{wm9�-��ߎ�}��T�D���k/�X_<�31e؄�5�5�7^�3���j          @���[_z�����ک�F&�	�ۓ�/Ʒ_�+��[���T��H�B��%��zI�4��ѯ�o�V/o}=���G�д;           -ڲ�q����_����u�N�jO˾��w������xp�������y7ǩ#g���XxO���          ��Zְ:�����Gf_�qUTW�d��#���xd�S����;�ښ�T��+����n��FΊϜ��7�<��h�h�W?�-�y�}          �)��~ג��uO�'�~8�7���d2Q��Xw�~Olػ9J]I�]^߱<��ؗ�I������G9��v�c��{�?���          �&�`��_�G�=7��P̩��bݞ�q���孋�\�E��h�h���<�Z�L\=�����+cX�!Q�ڳ��T�Kqc���          �nY����'�����}]I��k���\��uatvvF9)���ˡ�ָգ���_�E�ώߝvEL26J����ܝ)�y"v7�          (5�v��S�M�͸*έ����(vIȾ`�Ҹ壇���(We�wI&�?����1���r�E���D���Ql�;4�����/EK��          �R�fO}��߉���eϏ+&_�kj���i�Olx>[�l�qpG����[���Ww.�/�{F\P7?N5;*+*#�6���mz%�����         @��۲?~��񳕏ĬS㼺yq~��\��V[��-�ͯƢ�ˢ�3�I��[�ښ��������i�fǼ�O�3F�)�o˶ǒ+�mK��m�c��          �)ۙ��;W�;�8f�g��g>&����~�o�ۖ�ko,����=�����=hm�MGO�L&u�F���5bZL6!����7yC��X�wS�ص6V4��ջ��"w          �Ȳ����aM�k�����3GL��çƌ�c���zKs[K����v�{��ص&7i���wC���i����u��~VUQ㇌��A'Ǩ�1�fx��?,��rx���}F���w=_����s/����bG��r`[����          ��K�_��uQ��2���?�.F�Z��&xh���8�����;Ε���s=pr����Z��M;c㾭��iW�q����%	�n���q$Օ�ѷ�O��lG4��          PX���掣��[;ZmA�����Û��F         ����/�;           � p           �           ���          �T�          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�          H�;           � p           �           ���          �T�          �
w           RA�          @*�9���Nw#�    IEND�B`�PK
     �9s[�Ƚׇ  �  /   images/ce527fa2-4558-4370-a5e7-21077342728a.png�PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK
     �9s["1^FHo Ho /   images/e2a053a3-24a6-43e1-ac97-395cbc045e87.png�PNG

   IHDR  �  �   �r��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ��IDATx���1mA  ���+w!`0�t ^z )�-(R^$E�}i��_]���s� ����\k�       ����|��5 ����cp{��朏��s p'         �%�          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     ���<F��~��k�fq�\��PVeqU������T��T��aIl���6�4���%��5�j)mm<j�j����J�"" �s>�V��@X�3�x$��?;3���_�y}     � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	w           � p           	���7�o�=���������r�l��ʲ����1(5���z��7       �Z�vm�1�@����}����c�3?�7�۲7�S���?p��͹.x�%K�
���q�GF]]]6={��#�8"�u����o����///�~>�y�>/         ��k��o��F�ڵ+���Ν;���cǎؾ}{6���Jl۶-{=I�~s
^E UEEE444dӫW�l���ߺ���UUU         t���ټ�bڏbϞ=Y�e˖x�嗳s�l޼9���g�>�;�\.�썍�q��G�QG}����޽{g�         ţ�����z�󝝝�u��,tߴi�[�q���}���������������c�9歨�v         `��r�^�ze3x��w<�w��x���^Ȃ��lذ!����ަ��>�?��8�㲨=���#          TEEE{�ټݫ���ׯ�b��������6x(UwJVuuu������          ]�{����ܜ�~�v��>�~��l�}��رcG@��S2�8�,b�O���������          HEMMM455e3al���/�O>�d<��Sٹm۶�b%p�h����'?��2dH�766F.�         �B�o�d~�<���M�6e��ڵkc͚5��+��;E#�����YО�UG>j///         �bҧO�lƌ���y��,t_�jUv�ٳ'�P	�)huuu1t��lN<���          ����!��ڲ��������}��ձe˖�B"p�����/ZZZ���'>��z         ����ʷ��mذ!���X�n]tvv�L�NAhll��O?=N;��         �ֿ�l&M��ms��b�ʕ��3ψ�I���d����)���E�MMM         ���իW�;6��_~9�ꞏݟ~��T�IJ�޽���5���\.          8�����7o�U�V�_��X�~}��$p��ѣG�1"�          �NCC�[����?+V��Gy$��]M��a���>dȐhkk�SN9%���         �ë_�~�L�:5֮]˖-��<�����t�#�<2F�g�qF�m          ғ_f��ܜ���۳����}�ƍ����C����[[[���,          (=z�c�f�nݺ,t�Gb������C�gϞ1r��8��3���>          (l�|6ӧO��+WƟ���x���;�	'��ƍ�aÆe��         (.�����֖�ڵk��{�������q�9(�!�СC��sύ���          �42$�M�6e�z�سgO����TWWǈ#���}��          JS�>}b�̙1q��x���O�S������RWW���q�YgE���          ���)S����_��{^z)�����Y�����ڢ��2          �TWWg��?��X�zu�}�������;Jccc�{�1r����r          F�=mii��g����+�zꩀ�"p�}����ĉc̘1QVV          p�����_�B�Y�&�׭[�vw�S�޽cҤI�v          ����2dH�^�:~���Ɔ��C�^�b���q�gDE��          �F.�����:th��o�%K��K/��63����7n\�;6*++          �B>t?����SO�B����7�iӦ�4	�K\MMML�81۫��          �����a�b���t��رcGPZ�%*�`�ȑ1cƌ�ѣG          @
***���=F������{��A�^�\pA80           E���1}��3fL��W��U�V�O�^Bz��ӦM�6��7�         @����W_}u�Y�&n���ظqcP��%���2Ǝ�'O����          �B����_}<����t��عsgP|�E���%f͚���          ����<[�<r�����<�@�۷/(�"�����͋N8!          ��t��=fΜ�G������nݺ�8܋L�[)�sNL�:5**��          �����c���q�w�믿6t���^x��	          � ��E[[[477��ŋ�'�
���TUUŔ)SbܸqQVV          Pj��k���+W�/~�رcGPx�N��s�F}}}          @�;��bРA��_�:~�ᠰ�TmmmL�>=��          �_=z�/�8N?��X�xqlٲ%(�4|�������.          ��6t����W�w�yg,[�,:;;��	�HMMM̞=;F�          ��֭[̝;7Z[[cѢE�m۶ ]�1p��X�`Au�Q          |4'�xb|�+_�[o�5V�Z�I�������<yrL�4)�          L]]]\u�U�|�����c���AZ�	�������hjj
          ����r���'�pB��'?�6��'jԨQ1{�쨩�	          ��jll�뮻.�.]��sOtvv���=1ݺu�9s�Ĉ#          8t*++c�������-��[����=!������իW           ]#�_���ӟ�4�x����'���-f͚�          �juuuq�5��=��w�uWtvv]OM}��ok0gΜ�ԧ>          ����b	�����rK�ܹ3�Z�èw��q�W���          @ZZZb�q��7�ƍ��#p?LN>��������           �ҧO�����zk�X�"��.��m����cڴi�5          �������KcȐ!��_�2�x����w�����袋���5          �����G}t���?��۷��������/����V          @a4hP,\�0~��ĺu�CC��������/�nݺ          P�z��_��cѢE�bŊ���bcƌ��s�Fyyy           ����2.��hll��K������r1eʔl          �Ɀ����;�#����C���".���1bD           �i�رQ__?��c�����'p?Ⱥw�W^ye4(          ��6lذ���?7�tSl߾=�x�QCCC\s�5ѷo�           JÀ�뮋�}�{��/N�~�80��ꪨ��          ���e�K_��o�9�|���������������           JSmmm\{�hѢx��G��N��1><,Xeee          �����lyvuuu,_�<�h�C[[[̝;7r�\           ����y��EMMM�w�}��'p?@���1k�,q;          �.�������"����w��#p? &L��ӧ          ��9�󢪪*�����	�?��lʔ)          �a�lWWW�m�������&p����"���          �����=���c���"��!p����b޼y1f̘           8mmmQSS��rK�����	�?@>n����O?=           >��ÇGEEE��G?�������r��vq;          p�����%�\�E�����K��?���ٳgǘ1c          �`:��Sc�����,:;;��#p��M�g�yf           
�G��]�v�m�����{�:ujL�0!           ���:+^{�X�dI p���>;&O�           ]aҤI�{����	�ߦ��=fΜ           ]鳟�l�ݻ7���(e��o���1k֬           8f̘�v�e˖E������5�ϟ�\.           �|�<w��,r��G��|�����^zi���          �ᔏ�/���رcG�Y�&JMI�q�e�Eyyy           � �7_q��o|#�{�(%%�y���}.jkk           %555Y����=�l���$�����ꪫ���>           RԳgϬ{��7����z��������K.�          @ʎ;��⦛n�}��E�+��}�̙1lذ           ('�|r̞=;/^Ů������Yg�           ��3Έ_|1���(f%����Ĵi�          �������'{�(V%�80.��(++          �B���b���o}+���E1*���G�q��Geee           ���������o��[�F�)�����<��޳g�           (�%��N����v�ݻ7�IQ�3gΌA�          @1ijj�iӦ�w�Ťh��#GF{{{           �s�9'6l�?�p��܏=�ؘ7o^           �9s�����c�ƍQ�.p����+��2���          ��UWWg��׾��عsg��
�s�\tttDCCC           ��>}���_�������3
YQ���g��O          �R���'N�?��QȊ&p6lX�{�          P��N��ׯ�����Q��"p����V��r�           (E��z��q�7�֭[�|��.���֭[           ���ݻg}�w�����BS����ɓc���          @Dsss�}��q�}�E�)��}��1iҤ           ࿦M����?cÆQH
6p�������(//           ����"�o���سgO���gϞ}��	           ޭ��1f̘��v[���O=��=zt           𿵷��O<�V��BPp�{�^�b޼y          ����r1����b��푺�
��܋.�(�w�           |��������w�������
�'L�C�	           >��N:)������L�޷oߘ2eJ           ��M�>=V�^�7o�TD����b���QYY     ��ػ�(��;��)00�.��4�R#�A��c�&z�9ɉ���$'�����I�;!ш�b7�=XŀH�D�I�����DQʔ;3��9Ϲ�/1̝�e���     _ݺu��+��o�1�����Z�i~׮]          �#WRR���_=rQ��M�6���??           8z�]vY̙3'6o��&��+��"�ׯ           ��%�\����"��t��F����7           (?C����z+f͚�$g��+��K/           ���_|�A���F����=��5
           �_������Ϗ|0rEN�%%%��{           *�i��3f̈�F.ȹ����(������           *N궿�������سgOU�qr/p?묳�E�          @�;��c��SO��S�V�%��f͚�g�           T�s�=7�x�زeK��9r*p��⋣nݺ          @�)..�"��￿J�9�w��%           T�#F�K/�+W���?CN�yyyq�e�e�           T�������K㷿�m��r"p6lXt��1           �:%%%ѷo�x��w����<p�W�^�w�y          @ջ�Kb��ٱ{��J��*�ǌM�4	           �^�V���N�g�}���J�}��          �i�����cӦM�z�U������U>D          �O�W�^�w�yq��V��VY]ޥK��۷o           �{��?�|�^��������??           �M���1f̘7n\��g��%%%q�	'           �k������OǊ+*���$p?�s          �ܖ�����w�qG��_��{��nݺ           ��_�~ѩS�X�dI��W����}           ��ԁ�3&n��
��J����           T}��Ν;ǢE�*�~*-p7�          ��:��s㦛n������}���Ѿ}�           ��9���{��1o޼
��J	����Mo          ���?������+��WJ�>x��8�c          ��k׮q�	'�|P!_�R�Q�F           ���ѣ�o�޳g�h߾}           P����+k�W�XQ�_��w��          j��O?=&L�P�_�B�T嗔�           5�����G��?��\�n��G�����           ��(,,��#Gf�{�~ݨ M�6�           5ϩ��O=�T�����׬�����OϪ|           j����6lXL�:�ܾf����ՋSN9%           ���8�x�����\�^��#F�����           5W�-���1cƌr�z���ȑ#          ��o��ѹ����y��          @�שS��ܹs,Z�訿V�rJ           P{��<���-[�	'�           ����z(�m�vT_�\�#FD^^^           P{ԩS'/���Q}�r����c�С          @�3|���	����M�4	           j��;F�bٲeG�5�-p?�S          ��+Mq�ӟ�tğ_.�{��ͣ��$           ���&M����#��r	�������           ���_�~0 ^{�#����S�~��'           >���޽{GӦM           �t��ڵ�U�V��u�>lذ           �}N>��x����*p/..��={           �3p���4iR�ݻ��>��~��Ea�Q�          �i֬Yt��9.\xX�wTuz��          ���޼���FIII           �?K��C=eee��9G����?


           �Y�ƍ�k׮1o޼C��#�SM           3`����5jݻw           8��?��QVVvHD�{�����           ���7\}�ܹ���G�80           �������&M�D׮]           �H�������={�|��v�>`�����           �"6�����={�~�a����           8T�{�.���~��ѵk�           �C���'~��V�ޫW�(((           8T-[��֭[ǚ5k>��+pO�<           ��={�_�����Mp���m۶^߾}{�ݻ�S�N)**��z�YV�^�          *_�ѧM���sȁ{�Ν�A� Gc׮]�iӦ���c��ͱe˖غuk��p}�J����Ǝ;b��ݱs����={����N�:�J�{��������ׯ���o�{�q��ѨQ������u 
         �w��{�%<�C.�N<�� �ϓ��6dk�����/jO�zUK?���I��*E�M�4ɂ�f͚E��ͳ۴Z�h�ݦ8         �?u�֍nݺŜ9s�1w K��?����裏b͚5ܦi���)�W�>��4l�0Z�j�[�>���c��y         ��z��u�{
�:v� �7n��U�Vp{�S�k�-[�dk��şz_��޶m�l�k�n�m�         j��={~��)p/))���� �fJ1��e�b�ҥ��%KbӦMA�HS�Ӛ;w�oO�{�P֡C���{Zyyy       �^�v������ۣ��4{yϞ=��;w�ݻwǎ;����y��ԩ��}�ի�@�����������կ_?�ur= G�c���-[�ڵk?�������# �RX�����hѢ,hO7T���ͬY���O�F��S�Nq����_�       �����6d���͛��~��[�f�z��sɾ�=ui5l�0�6m��6n�8{9�k޼yR�@-�����⋟�>�;@VVV+V�����g1{Z�ׯ��t���{�e+I�����w��%�u�mڴ	        ���}͚5��裏�f#��7fa{��^]�&�ɻ����f͚e�{�-�պu�hժU�� ��Q��J�!@�KA����c���p�;wn����c�޽�z��l���k��҅`��޵k�())�:d!<       P�R�����=[+W��?�0��S�^ZZ�#�Ok�ҥ�z_�Ҕ��(��]�vѶm�l�	� �\�wK?R�Ͼ0p�޽{ ��V�Z��~̙3'�����I��f��V���J�{:���O�vA       G'M+_�lY6|0�i������5�[�.[i��'g�{��۷o��;��c���( ��4h�=Ƨb�L�P�lٲ%fϞ�E�i�c���6o�o��f��6m�d�{Z)|�[�n        �-E�i��%K��im۶-�<����O~~~�Aw�q�J'�w��Q�PMu��M�P]�ݾ��n���{1o޼سgO��Jǟ�5mڴ�S�Nv�K�޽����1_       P��ر#V�X���,�ŋg���=iZ��ի���odo����=MyO]D���� r[
�_x�O��s�F�E�֭�ʕ����}�̙YԞ�a��k׮���|����}�{��      ��n�ƍ1���+��ij;��'���ӧgo+..�B�N������[� ��!�n����b�����E�bƌ��[oŦM�*Zځ��SO=�Ms�ׯ_0 �t��9        5Bj0� �>� �׬Y�l۶m�Y�fe+)**�Z��D���C��#7n�Z������܏?�� ���޽;fϞ�E��	���������c�ԩ�jڴi�4H�      @��N7_�`A�ϝ;7�-[fB{-WZZs���֣�>��;w�b�����T��x|X�{� �W�`Z�pa���曱y��\��c{��լY��߿6�=�       �&�qi��{ｗ��i� L
������-[F�^��O�>ѽ{��S�N P9�@��ӧ��ѡC� �|�Z�*��׿fQ������u�d�c�=6C���w       �
eee�|���Q�ҥK��ڵk�Lq{ ػw�l`ӦM���Y���o�>�֭ ��۷�[o����ij;Tw+W��?�����#�dGt:4N:�$�       �p�v�9s��̙3��wߍm۶����l�t��z(�,�N�O}D��@�J�zQQQv��>�Ӄ2 �o�޽���^{-�y��I/�4������dS�O>���رc       @y�Ϙ1#�0v��PYR�hѢlM�4)ڶm�Mu8p`�2 G/???:t���������5�Óv�I�S�N͎-��"���wLWz�p�)�d�{�U       ����,>����>}z6���]�*�^�:��l�݇�Z�
 �\�N�-pO%< _l�ҥ���/gU��Sۥ~��4hP�92�=��       �ϓ&e/\�0����o��͛r�'c�4pȐ!Y+Ѹq� ��w�q����{aa��3 >G
�S�>mڴX�re JG¥�iu��=N;��۷ov�       �f͚��_���6TG�N�4)z��'�|r���'


�/�σ�?3po߾�V�ϰiӦx���^�-[����͛���-[ƈ#b���ѠA�       �vJ�g͚�M�;wn6�j�={�d��*..�ĩ������ �M�6Q�n�عsg��g�L�dɒ��_�o��v�D8|k׮�ɓ'ǓO>��TNS�[�j       ���H�g̘���5ٶm۲Miu��18dȐ(**
 ����{l,^�8{�3��P[-X� �y�lW%P>v��S�N�iӦE�޽c̘1ѩS�       ���7���矏��FK�.�֤I�bРA��|������{*�j�t��{�O<�D�s��{m߱\]�t���:+���       T�W�Φ�O�>=�o��?���Z��0 
��k߾���?�Q�m۶P��޽;^{�lb�ڵk�<i��m�ݖMr��W�}������       ��H���Ν��Ꝇ�ׁϖZ��z�8����N��M�@m��~�S�{z�,..��"��o��VL�2E�U,��0v��h׮]�y�1d��;      @�+--�7�x#���lr;p�6oޜ�L�?i �Q������&5c�~�;j������'�x"6l�@�X�jU�?>��K�����#???       ��q���˱m۶ �\j�f̘���ݻg�DϞ=j��F�F���?w��ٳgO���Yؾq�� r׾���瞋��;/۩      @�Z�v���}׮]��y��e��c��ѣG��c���>��m�6 j��{���o��<�H�Y�&��cŊq��gGp]p�QRR       T����4��7ވ��� *�ʕ+����=�X�~��q�)�Dݺu��J�g�mڴ	�����ߏI�&������/^���o�G�q�Fǎ      ���hѢxꩧ�����kݺu���f߇��zj�5*�ի 5�1���
܁-Ű?�p,X� ��#mZ�;wn0 �[�l       ��}a��Y��z�7o��<^x���,tj�V�Ze��EEEѨQ� ��6l�O<�D���+vC����z뭘9sf�;��sύ���       ��,\�0�L��rϖ-[����_�"������kݺuv[��o����ꪴ�4�}��x�gb׮]�|{�쉩S��믿g�yf�~��QXX       �U�Ve��3�}i���ɓ�^j���q�i�E�:u��jٲe������PݤI�/��r<��c�7��ٺukv��ꫯƥ�^�z�
       �غu�⩧��~�ZVV@��&��f�^���>;��� �Mz�j޼��'�T7K�.��'ƢE���?�[n�%����]vY��      �O۸qc<��Y؞N������ǽ��S�N�.� ��� �M���`@u��5�c��M��Mp��Y�fŜ9sbĈ�E[QQQ       �s�ά�x��'cǎ�,�V���o�=:w�_|qt��% ��Գ���� �.��.��L�۷o��ٽ{w�+��wމK/�4���       �U ���oǤI�bݺu�l�-�믿>N:餸袋A��Գ܁je����1:K�,	�C����;�O�>�}-Z�h       ��ܹs㡇�+VP{��-3f̈Y�f�g�g�uVԫW/ rէ�f͚@.JGc=�����s�e��D�XK�h3z��8�쳣��        j�6�#�<ӧO��ڵkW<��S��k�e�܇yyy�kRϾ?p/..�+�I��NL�81��8Z�6̼���o|#:u�       5��ݻ��_�G}4JKK ���c���1mڴ����u@�9`�{ӦM �l޼9~�a;��
�|����/Ç�K.�$���      �&H�[?���v�� �,K�,ɺ�4���/�F�@.HM���=�s�3f̈��?��*�޽{��_��s��UW]ݻw      ��j�ƍ1q�Ę9sf |��M��iS�E]�	�����TXX��{�&M��mڴ)��~�� �,}�Q�����i�      @�TVVӦM�G}4JKK�pl۶-���x�����_�z�m�6 ������@UKS���غuk T�}��?�����ꫣs��      ��-[���K�.��1����Og�qF�{�Q�N� �
��ƍ@UرcG<���YX
P�֬Y�_}�5*�?��(((      �\�&�����^x!�P����<�L���;q�UWE׮]��	܁*�dɒ��{�� W�����ڼy��k��֭[      @�HS����?�-�
���o~�>|x\r�%QTT �E�T��>��s�裏f�� r��ŋ��?�y\|��q�)�      @UڱcG�ZL�6��v�¥Ǚ�_~9�̙�Ms/))	�ʰ?poذa T�u�������� �.�ѽ����~|�߈���       �l�g��~w�~�� �L�������iH�i�@E��7h�  *ڌ3���m۶@u���D�k��&�u�       �a׮]1eʔx��gMm�Lz�y饗��6��ַ�K�.PQ�)M@����c���P]�I7�pC�92��կFaaa       T�իWǸq�bŊ��4����7q��gǘ1c"??? �[Ve�׭[7 *¢E��������K;��N��=�}�;߉-Z      @yJ��|�W����;w@.)++��<�̙�\sM�j�* �S�7k֬(/// ���/�'N�ݻw@M�dɒ�����ճg�       (�7o�	&�{� �,���~�_~y:4 �K�7mڴ^ ��]�v�������j �T[�n�[n�%F�^xa�0      �ٳg����شiS T;v����ǬY����F�����@9ٰaC�q��tc��.��3���ի�ꫯv�      �4Hp���1mڴ�w� �͌3b���q�5�D�n��hd�{qqq� (��͋��+;.�6I;�����;����h׮]       ��+W�=�ܓ�Tg�ׯ�n�!F�_��W���0 �D��QTT$p�J�=����#�<eeeP�Y�&~��_�UW]      �����/�ĉc���P��l�ԩ�lٲ��w�M�4	��%p�ڎ;b	���o@mWZZw�}w̝;7.���(((      �OڵkW����+P-X� ~�ӟƷ���8��p�ܝ�?�0Ǝ�W�j����hذa�۲iӦ�z��W�ݘP��I��߳�ȍ7      �dÆq�wĒ%K�&ۼys�x�q�ęg� �*��֭k�;p�f͚�ƍ˦S}իW/5j4H�X���!�ԩ��~�����y��׏���O}Ϳ��o�q�ƀ�n����_�"��_�5�;�       j�y���]wݕE� �AYYYL�<9V�XW^ye�|�;pD�d�?��O�rS~~�����mڴ��m�F˖-�U�VѢE�,lO�zyK�!p�H�������k�_�~      �>��g�}6y��P+����jժ��w���K �'��������<[��w��%N<���ڵk���ѡC��رc6q����}���C:�"18f̘8��s      �=v��&L���~; j�4��g?�Y\}�Ն�k_�� _`׮]����>�z� w����N�=zD�n�8�gԨQU�gJ�;p�}��D�+��"
      ��>���;vl�^�:�Q�F�Ջ�?�8��J�~Ґ�ѣGǅ^yy�U�Ӳ�����#�6o���v[,^�8�z��q�}���^�zEQQQ��;\:Yaݺuّ[���      �fJ�� �t�35Gf��֫Wo�˩�(((�n�`�t[\\4�VӦM�y����������?P��!��<�L���k��O ���yyy�pk֬�[n�%��j�m�v�ްa��Uw�|s�΍_���q�u�E�f�      �Y���x衇����!��-Z��V��4i���"���p=M`?�
�?�f͊_���o��oѦM� �'�����	��gZ�pa�~��e˖�j���={������:Hxig�����l�V��_����}/ڷo      @�WVV'N�_|1�=�e8��G�1��شiSt��)[�s�Q��"�yyy6?�������W���~��ѽ{� HLpꭷ�ʎ�ڵkWP�:v�'�tR�x��qV�M�q�|�� n�ƍq�7ĵ�^�"      ����Ҹ�����rG�WRR�E�)d/((�ޞB����4>�����[��M7�W^ye:4 ���IO=�T<��v�V�t�U��~��'W�cw�ph�m�7�|s|�[ߊ���      P�lذ!n���X�bEP�RD������7�t�?j�i����{��l�~�w��j�� �'S�L��<�<͚5�dۋ���&H�;ph�Iw�uW\u�U�/})      ��c�ʕq�-�d�;U'???�v��{��&���=W��b�(c}��'cݺuYC������~`��ᡇ��>��۷�aÆeV5mס�OYYYL�0!v��#G�       �͙3'�����|T�&M�dQ��A����M|��_=>�����w��������V�{��ꫯ+���|:4;��r1�/m4z���c�F�      @�z�W���˚*W��|�	'Ā���lѢE �o�ܹ��_�:���h֬Y ����?5x���A�IGa��ib{�֭��KO,

bϞ=��?��ñy��袋      �-�wz�'O�g�}6�\�5ʢ���GqqqTW�¡Y�jU\��Y�~�1�P{ܡ�KS�Ǎ3g�*F�%|�'�i��V�vঠ�y����Gp��y����/�v�      ��JC���?�k��T�v��Ő!C����G��7nEEEQZZ��[�n]��W�����N�:P;ܡ۹sg�;6�̙��4��W�^1bĈ��GK��w8r)r߾}{\q�"w      �bi���~���1cFP�Rw���/}�KѦM��iRK��S_l۶mq�7������ҥK 5��j�����o��s��+E��k�ȑѬY���Z�j��~ G^�����oֈI      P�����w�y'�Xi�y������I�&QS���w8ti@�M7��^{m���#��M��P��v�-�ĢE���չs�5jT�m�6�Z;���믿;v��|�;QX��      T�4�j�ر�U���СCc���Q�^���R���x|뭷Ʒ����ׯ_ 5�B
j�H��Z�.]������g��:u
�O����w�}7ƍ�E�&�     @�H�����A�ٴ�!C�D�:u��04�L:Q㮻�o}�[1`�� j&�;�";w��v����O�ƍ���O�>}�D^^^p�t1����ݻ7��7s�̘0aB|����      l۶mq�M7Œ%K��W[��}Lp�#�gϞlH`�:lذ j�;�i��w�����^��JX#F���u�����(5j�6m
�|L�>=


��+��     @I����c�ʕA�*..�SN9%���7_KC���eee�����?�1��ӀR�f����I;���Θ={vptRLڻw�8�3���|���X����W_�z��ť�^      @�Z�~}�����5k��'<xp><�}gm���&M�Ć82{��|0�o��sN 5��j��Sm���1k֬�褝�g�}vt��%8t)p_�hQ �����&�@     ��v�ڸ��ȝ�N�0`@�1"6l���T���M�2%��P@�!p�,�P�����7��\�:ubذa���|4֑Jc@�Hh�1��3�      ��lܸ1��.n/?�;w���:+Z�n|Zj*�ϟ��KEj��cP�)5�{���W^	�\III|�+_Ɏ���ܡb���Ύ�;��S      82�7o�o�1����K�@�խ[���Z�h@�IE���8� �7�;�P�'O����/��iРA�=:����;T�tZ���ߟ]���&      �óm۶���c����ѩ_�~�92������T@�KCaӠ��ÇP}	ܡz����g�	�LϞ=����"w�^�F����(JKK�)r���{���E      ��ٱcG�t�M�lٲ�����E�>}�a�z�C'p�����/k(@�$p��W^�)S���q��q�9�D��݃�.b��ʕ+�8eee���.6l%%%      |�]�v�m��K�,	�\�6mb̘1ѡC�����I�i�P~RC1~��,rO�o��G�5��ٳ��g�4�=]l�O��cϞ=q�wď~��h׮]       �m�������͛��u��ȑ#cȐ!�����T�X�"���;�3��_�%kÀ�E�5ĪU�����v�q��.�Q�Fŀ��ӢE� *���۳)?�񏳓)      ��;�o�[pd:v��w�����w��63]w�uѭ[� ��;� 7n��o�9�9t�;w�.�@ Z	�nc��]�6n�����~��      ��޽{c���1cƌ���$x�I'E^^^p�4P�v�ܙ5������9@� p�jnǎ��6�&�5bĈ8��S]lUcP��.]�ƍ�k���q�      ���w�}��o����$ƌ�5
ʏ�*^j�� ����Ѷm� r����td�=��˗/M�&M��/��;.�<�8�ئ��@�5kVL�<9{�     ����'���_~98<���ѣGǀ��'p�ʱe˖��[�'?�I4n�8��&p�j���EM�=��΋������� �5k�֭�r=��s�&��#G      �Vo��V<��c��I/���h޼yP1�[C�r�v��[o����� w	ܡ�z���^�X���:�4hPPuҎc�;T�|0�G��}�      �6��Ϗ����޽{�CSXX_��cذa���T�Ե4m�4֯_@�[�ti�7.����ls	���P͘1#y�����d.��lG1U+�|�A �/��Ogir�N�      j��>�(���ؽ{wphZ�j_|q�i�&����C�5kVL�4)�ʀ�$p�jf���v��;fOB6lT�t1T��;w�رc�?��?���      P�mݺ5n���ؼysphҩ�cƌ��u��'5�������/ɾ�F�@��C5�.�Ү�]�v���:�����Ow�L�C�۸qc�v�m��(�ԩ      PS��"�nl͚5�KA�9�}��	*���ƃ>͛7�6� �E��DYYY�u�]�aÆ��
��s���#�#̀��lٲ���{�ꫯ      �������b��kӦM\z�ѢE��jܡj�&oܸq���?�?�� r����I�&9��4j�(.��h߾}�{�ի6�-[�P��O��:ur�      5��ɓ�7��X�޽�A�i�;U���:;wc�Ə�cߋ�C�P̜93������9昸��ˣI�&A�J;���1[�ڵ�N8!      ��x饗��g�>_~~~�v�i1|���5h� ���c۶mT��?�8n����я~�����	�!ǭZ�*Ə���g�ѣG\t�EQ�N� ���}ɒ%T�t���w���_�͚5      ��.\'N>_�F��K.�:�#M��C�I��]w������M@@��C۱cG�C���4�lC��3�<3������-�7o�;�3~��Fa���      T_i�n��מ={��k۶m|�k_�&M��%\�|y UgΜ9��c��\@�R2A�J������ի�OKA�駟j�U�V�ŋ��ɓ��K/      ��RԞ�ȝ��ٳgm֩S'�=�Bnx�駣}��1p�� ���r�SO=3g�>-MN\�z�
�����=�?�|t��%      P�L�81,X|�4Dpذa� ��2�IS�a�`�֭[G��w�A��~L�2%��z���W\��C5��8K;�w��@n�0aB�k�.;�      ���^{-^z�೥��_t�EѣG� �	�!w����;������P��c6n�w�}w���JO����8�c��)�OGj��� ����Ƹq��'?��#	     �V�X���ي���k_��!��D�f͢�� ���@�[�vm��]w�u���@��CIǛ�?>�n�(M��ꪫ�8��-�8�CnJ� 8iҤ��       ���b�ر�s���Ӛ7o_���u�H��S䞢Z 7�������O��g�@��Cy��b�ܹ��R�&��ȝ�ϑZ�ۦM�%%%ѯ_�      �\��s�=B��h߾}\~��ѠA��zIM��א[{��ԩS�x�T�;��˗ǣ�>�M�6��v]5��r߄	�c
�T      �5���={��c�>��:�Ï_��Җ����e�K�jX�l��j�؊�=��˼�8�E�v��$��E�U�UHt$$!�*zG4�����h�([���g�_$v{�9�>�뺃ˍ3&����:����򣩀ғ��~��_����0`@ �C�%���1~��_GSSS�aÆeq{�޽��p��w����p����,*++      J����c�����&L��=�XTUU婶�6��s�ԩ�������Gt�;����~:���|j������XܞC)pO/z---��>� ���C=      P
N�8��F���r�3fd��UTT���@(][�n�^x!}�� :���؆��^>5bĈ,n�իW�?ݺu��������(m�`���}-F�      ЕR���_�:Μ9\쮻�o~�A��Ci�7o^|��_�q��б�Ѕ��%&�/6l�0q{���J_�i!����?�yTWW      t����\�[��V�y�A>�^���� ������W��_��ѯ_� :���H��Kq�ɓ'��?��O����>� ��w���x����'�      �
�w��>�TEEE���1{�� _RS!p�ҕz�������}�w1�1��E/^��np^mmm���w��A��R�˒%K���.Ə      ЙΝ;���MMM�y)�|��b֬YA���f׮]��6d��}��@��Cؿ̝;78o��Y�ާO���P^ҭ#����㗿��A$      :��O?��:�y)n��c�̙A>i*�<<��s1f̘���hw�d)���~���AD߾}�?�i�ScP~�?�<�L��'?	      �iC�e˂�R�������Ӄ��T@yH7����g���kTWWо���,X۶m"z��?�яb���A����d[�Ϟ=@�X�bEL�6-���      :ҩS��7��M�H����o�����6��o߾x������}	ܡ<x0^x� �����1lذ��ҁL����C��̆�      �#��=��'O�λ����;��/-��֭[�(}/��r�(�_�j �G��$�~���Fccc]eee<���/})(�t���ݻ(/G���s�fCJ      �/^��npޜ9s����!u5)r?|�p ��m(����e�Ў��I��k�֭A��?�ƍ�m�����W_}5�M�f�     �vw���l��͚5+��ޠX��@�;��#G�ĳ�>?�яhw�Ǐ�?���A�]wݕE�P[[@yJ�ǿ��������      �������o���A������'�@yY�lYL�:��Wh'w�O=�T444D�}�k_���/ q��6g������|'      �=���+�u�� bԨQ��c�EEEEP<�B�ICZ��������ߢG���;t���z+֯_E7bĈx���������[�n���@y�7o^L�>=�      p#�9�?�|p����~�}�N1Y���ѣ��?�9����pc�A����?��Qt���GQ]]Ц��2�
�<��?�����       �-m���o~Qt�{��Xt��=(.�;��ŋǔ)S��n��	ܡ����ǏG��W�*���	�T:�	ܡ�mٲ%֬Y�g�      �˖-˾w*�^�z��C�ѳg��ӧO�>}:�򒆶~����/~�7q��:Ⱦ}�bɒ%Qdi�>C��ǐ�<�LL�81z��      p-N�<s�΍���������G��gA�����1����w����CHSXO=�T���D�}��_�������`�p�ԩx���_�     ���ӟ�gϞ�"Ky�5jT@��T�ܹ3��4o޼�>}z6,�k'p��v���_�5v��,p��#p��H���q�q��7      \��7�믿E7gΜ�4iR��4Pޚ����C��g?���k#p�vV__�=�\Ymmm<���>��B�0�~Nҭ@yK����K������      |��������7n\�s�=�J�P�Ғ�5k���ٳ�6whg/��R�8q"��{����OF�=�H�y�۷o�<y2��u��X�n]v�      |��W>|8�lذa�lp�|x�gb	QSS���C;:x�`,^�8����!C�\����!G��l�ĉ�       \ɡC�b�Qd�{���^��2`���֭[455P�N�:�?�|��?��	ܡ=�쳅~��1cFL�4)�Z���m۶�Ǐ�~��      �J���?�������}�{1p���ϒ6����f7����k��]w���rK WG��d˖-�~��(�#F����p�\�����/g����      \(�6l�"�ַ��F�
�"���C�kii���z*����9^����Akkk<��3QT麬'�x"�	�U�6򥡡!�^��?�q      @�����}ERWW�g���
ȏm۶�ڵkc֬Y|15*�����k׮(��~�n���ȧ+V�׿�����[      �ġC���R���#�\-M�˳�>�&M��={���p�������dq�Ѕ�կ_�쥭��>��H��<��s���      'N�����GQu��=�|���ѣG���C�|��G�g�c�=����Z�dI;v,�hРA&�iiJ}�޽��{ｗ=�ƍ      ����s444DQ}�;߉!C�\��STTTdƀ|X�hQ�}��ٟo�	��|��ǅ�.����'�x�d1�"M�!��Νcǎ�~�     @1�ٳ'V�^E5y��8qb��J]N߾}��ɓ�Cccc6�����|6�;܀ę3g�����7��\���k׮x��cʔ)     @1=��3���E4hРx���W��,p�|Y�vm�{�1r�� �L���ԩS�x��(��Çǜ9sڋ��-mq�4iRv�      �����{�ETUUO<�D���Wj*v��@~���������������rw�N/��R���G�t��-{���E��v������;�#      (�����瞋���7�7�|s���T@>m߾=֯_�'O�rw�ǎ�e˖E}�߈�C���t%[�hnn �^|�Ř9sf6(     @1�%H���"���g��Qwȯ46q�Ĩ���b
#���͋���(��n�)n���������Ƒ#Gȧ�G�ƪU����      �/u/��RQϞ=�G�����U[[@><x0֬Y�Ƀ+��5:~�x�\�2�&ȏ>��i1:L�8�C���/�e��     ��k��V��z��߿@{H?K������@����1c�-\�F���/���9s�Đ!C:�+� ��;�]Cy�]w      ������͋";vlL�81���� ���?G��e˖�7�� >%p�k��GŊ+�h�*F�ùR�!mq�={��c     �{�W��ɓQ4}��Gy$�����wȯ�R�q�ѣG� �S�5H$E��2;|UUUt����i�x͚5q�w      �������~���ݻw@{K�;�_i(l�ҥq���p���R�)����ӧ�M7���Ơ8�ϟ��~{6D     @����gϞ����׾�ƍ�����ۂ�{������ҢE�
��=]�u��t��={f?s�O� �:o��f6D     @~�����ŋ�hz��=�P@G�4�/5S���j|���@�W%��-[E��<I�1t�t �C1̛7/�M�     @>���gΜ��y����n�Q����jkkk ����/�׿�u[�!�pU�dTѮ��җ��Ǐ�L)p߹sg ��gϞx���]�     �iy`
܋�+_�JL�4)�#u��=���}�Q ������k�o}+�������
w}VUUU|��ߵU�N�J-(�����     rbɒ%���ޭ[�x��:Cj*�,ȶ���(2�;|�U�Vŉ'�HfΜ)4�K���bI�ӭ#G�      �Wccc�&w�}w���t��Tl۶-�|;y�d�\�2�瞀"���hmm-��Y555�t�;ϢE������     ��|��,�+���y���0�cΜ9QYYPTw��6m����G��{�ѳgπ�п��z�s��P�֭�����_80      (?---�[�<��ѭ���ci Ǒ#G�7ވ�3g��,�E;�6,�L��U***����@��_x�����c�      ����_�ÇG�����m��Й�P,/��r̘1#멠���<�mp/���ߵ&t�t �C������=z      �e�Q$UUUq�}�t��}�fߩ644�{�쉍7�����H��!moomm����W��F�
�j&��xΞ=k֬�9s�      �#�w�w�"����cРA�-mq����}��Pi���������n���Q���{�(w(�ŋ��w��j-     �2��IMMM�u�]]E�Ųe˖صkW|�K_
(�;\��U�
u�ϤI�bذa�@�Ŵ������E      (}�M�6E��s�=ѳgπ�����Y�ti���?(�;\���ˣ(�u����7JE�6������� ���W_�     ��E�EkkkE
��N�Е�P<k׮��<���P$w���͛u��̙3����"]0 �;@����[q�ĉ��       J�ٳgc͚5Q$�������*�+	ܡx���������w�D��HE�B��o�=�Ԥ-�w(����X�jU<���     @�Z�lY444DQ�9�MĔ��STVVFKKK ő��x ����B�8y�d����Q3f̈�}������|@���kq���g��     �����H�+**���P
�2�~��e7c�q�ԩX�n]̞=;�(�p�+Vd�c���vJY�8�)�ްiӦ?~|      Pz6l�G����4iR�1"�T��_���
(-�S$w�?����r��(�iӦe�P��a(�4p&p     (ME�ޞ��{��$5[�n�X�m��w�[n�%���ҋߡC�����;�(Uw(�w�y'�^�o߾     @�h���(,�i*���-[?���@���H�ۧL�� FI����޽{�ٳg(����x���m�      (1i{{KKK�偔���� �i�����ODϞ=�N�����!�|��(���*0�B�8���(��˗�     JHZRdy t=ܡ�R�v�ژ3gN@�	�����Q__E�`(uw(��{���ݻ�[n	      �������ɓQ�R����mo.J�\,-�Sw�_�V��"p ���8��'�|2      �zE��>y�d�)i�����0�xv��{�쉛o�9 ������c�֭Q'N����;�����������      �Ή'bӦMQiy�]w�P�RS!p��J}SOy&p��֮]���Q�g�(w�ԩS�y��7n\      �uV�^---Q�R�w��R����G�n`��O7���"=zt:4�\����KXSSS ŕ>��      ]+�tE�n���r`i ۙ3g��wߍ)S����Bۿ�ٳ'�`֬Y�$�� M<x0��z��7�?�aTWW      �o۶mq���(����flʁ�X�r���\�Shk֬�"H��o��r�dw(����l�x�ԩ     @�[�zu��픓A�e?�---ӆ�ԩSѷo߀<�Sh���zA�ޞ^j�ܘ8��y-p     �|���ٍ�E0v�X�QS6�u�-�<v�X Ŕ\֭[��sO@	�)�]�vő#G"�w��*ʖ�߀$M744D�=     �γq��8}�t���PN�@���--��Ww
뭷ފ"�<yr���3����s��e�<��     �s�]�6�ছn�[n�%����b˖-׶m���ѣ���Kw
��{EEE̘1#�\��X�9nmm���՗w     �Γn�}�w��㎀r#hRS���?��y#p����������(Wݻw�~���G}@����������     @�{���=��ƍ(7ii �����SHil̚5+�ܥ��������{/&N�      t�7�x#�`�̙QYYPn�@�gϞؿ>< O�R�2λt�J�����QUUP�ҁl۶m��[o	�     :A���K�O�<9����D�^���?��RO!p'o����ǳ���kii�g�y&���ƦM�(7&��6��n���FEEE      �q�y�hll������޽{���T�޽;�b{��7㡇
��;��~��,�+�ӧO����cŊ1jԨ,t7n��(w�ͩS�bǎ1z��      ��M�E0cƌ�rV[[+p��>���;����Q���oߞ=}���I�&e�����2�;p��9.p     �8is��"�7�tS@9�T m�pڷ��퀼�S(�Ν�-[�Dѥ���S.�@FϞ=���> R��裏      c�ƍ���y�������M>E��m�|�M�;���By���ȝ�.��>hР�:ujL�2%jjjJI:��ٳ' ҵZG�ͮ�     ������Q)ܴiS�����ٳc�������@��;wƉ'b��y p�P��W��رc�hѢX�dI�;6�Ꞷ�WTTt5�;p��5dΜ9     @�J���w1E�n_�n]��F"������
(i�e�ymnn���g��⮻�
��;��6����o:��'Eœ'O�6����;���8.�6i�     �ߎ;��ɓQ4)
ܾ}{����7&M�ӧO�������s�n�H������8t�P9r$�z�?���}�ҥ1f̘lRy�����Up��6o�---QYY      ���ݩS�b���bŊO���7�wS����R�$ipcccTWW�;�;����r}���>��B�4�<eʔ�޽{@gH�1�6gϞ��;w�     hg��Npޅ[�S�N�Z�����R����$���!�l�uuu�N�Na��$n��Çc޼y�x��?~|̘1#�Б�]���� I�\�     ���Ǐ�޽{��;v,-ZK�.�1c�d[�}WE�����6�6�;y p�ZZZ��$�O��Z�n]��1";�M�8��&t�����ȑ#�����      �ǆ���|����ظqc���ٓ'O�z�^�zt����&��7P���Ν;��ٳA�طo_�,\�0���5kV2$�=���h��������={      7nӦM��K�_���˖-����ǌ3bذa�m����&}>����N�N!l޼9�x)4�p�{
��!.m߆��Pssslݺ5��     �ƴ��h+�SCC�E�D��>q�Ĩ�����޽{[�	|"�͙3'��	�)�>� �\i��ܹs���mWr80�z	܁K��w�;     ������̙3��I�DzR+QWW�-2dH@GKME�s����{wʞ���KS�۶m���ӧc���bŊ5jT��7.*++�����6     ���6��~���?��~뭷f��رc���*�#܁����Y7�ѣ�	�ɽ��t����ؾ}{����7&M�3f̈���\�����v�ܙ]�أG�      ���M�t�ԭ��O�>1y��>}z0 �=���@��g�fM��ѣʕ���۲eKPZN�:�mu_�re�9�Vw�J
X�pD��H���cǎٶ      �Ϲs�eut�ӧOg�Ċ+bԨQZ	�U��p���]�N9��{|�AP��5(m[�S�N�)S�DMMM������P���     \���}SSS�9Z[[��;�;p�����
(Wwr-
�m���cǎŢE�bɒ%Y��&���rEEE@�t Kۚ�lݺ5      �~v��e���ѭ[7�*�'� UsssTUU�#�;�v���8s�LP>҇�ƍ�'�̓'OΦ�{��`���Ν;�A\�     p}҆W�֕Z�����+�j��KS�Z)����!>���lp
ʑ��\KSH��#G�d��K�.�1c�d��ѣG�%p.U__��n�)      �6i۳[�K˅�D]]]̞=;��ERS!p.����+�;����@�6�<bĈ,t�0aBt��=(�;p%i�M�     p�RW������J�_�>{�Z��'Fuuu�������>�������ʑ��\��Ͼ}��g��1~���1cF6,(�~��e��Ν�6�����      ��֭[����J,\�0��>k֬2dH��,.�>�[[[���"���ɭ4a�w�� �bݺu�cR�8��V�8޿ �1�     p}�m������OZ�[o�5�ǎUUUw�R�q�Y��ʍ���ڽ{wv]�gR�XҁL�\(���~�׳g�      ���ܹ3(O~�a����'&O�ӧO��%p�$-�S���֮]��b�pR9}(��}���&�sƁ�T�NkϞ=�|%      �:��S�N����ӱ|��X�bE�5*�M��ƍ���ʠX�B�4�~& ڤ���;�(7wr+mp���F��s�f[�Ӥr:�80(w�J���     ��m߾=ȏ�*�w��~���ԩScƌQSSGmm�����{ʕ���J�0�I���Wb�     �ڤ����ɓ'c�ҥ�lٲ;vl�J�f���"ȷ�T�ڵ+ ڤE�����-PN��RSSS�߿?�ͅ��}���I�&e������K�6N
---��`     ��ٹsg�o��ͱq���I���ɓ�ؽW�^A>Y\*us�3?<A9��K)nO�;\ɩS����+W���#G��ٳ��n3�\&�u��cǎ@�����w      �/��{��	��ȑ#�hѢl�{]]]�J><��;p%�f�;�FD.�޽;����m[�S�N�)S�DMMMP�ҁL�\����[n�%      �|�{���Ơx��j�ׯϞ#Fd�'L�ݻw�_mmm \JOI9��K{���)�n�T3fLv�5j���%*�[�l	��۷O�     p>��À��Zz.\�mu�5kV2$(_�n�N� m|�S���R�4��^�7nܘ=)��<yr����+(�����?     �ձɕ���Ǻu�'muO����㣪�*(/i��A��СC�&�����=z�(wr)M�:r��e[�G�t=�;p%>�     ����ϒ�s�;wn��=-�>}z0 (���jmm�={�ė���r!p'wҤщ'�˅[�Ӥr
�'L�ݻw�����     �X���|�ӧO����cŊ1jԨ��7n\TVV�MS\I���SN��N�$M�1���+=,Ȯ�1cF6,�\�{�Ξ�g�@�ÇGcccTWW      W�n3������پ}{����/�N���555Ai����K��PN���t�tS��u벧m��ĉE��h����k׮ h�~�v�����[     �+KK��z�<y2�.]˖-��c�f�D��^QQ�܁+�URn��N
۠3�mu_�pa���ŬY�bȐ!A�J2�;p)�;     ���q����c�ƍٓ���<yr����+�z鿓4t���1�F���;�
�
�
�����zk���媪����R��Ç      �M�N{:r�H,Z�(��>f̘�={��T]�G�ѧO�8u�T �9{�l|��Gѿ��r p'w�m��?�0{���S�L�&��ܸt�َ;b�޽�?\�{      �������>��>bĈ���0aBt��=�|i����TzаQ.��J�ZG�F)I���^{-�/_��v[v�K������;v,�y�x�������y��     ��RW�{W:ھ}��g�QWW�f͊!C��'��J7�;6��ɕt�FCCC@�iii�͛7gπb�ԩٓ���r�*�?�U�VŮ]��j	�     >�ѣGut����X�n]����)t?~|TUU���6 .�ʉ��\���rp�ĉX�xq����D\��>j�([��|ؾiӦX�dI9r$ ��ɓ'�_����3      �����B�<w��l���ɓc���ق@:F��p)K)'wrE�N9inn��7fO��M�{:����;�(f_z�ػwo ܈4 s��7      �U��N�>˗/��+W�m�ݖ��_��W,l'�q��yǎp)���;�r�ر�r���[�`A�ٽ��.��o���(�������իWGKKK ܨ�w��     �r�6JE�6oޜ=�:�)S�DMMMpm�����~l۶-8���p%��lll����R'p'W{�_�>{��M*O�81z��y��,?����0@{9~�x      p�C�����ޢE�bɒ%1nܸ��9rd��Μ9o��F֗襀��`R�5|���R'p'Wm����㥗^��_~9ƌ�f���V�49���OG}}} �'��     �2�)e��ͱaÆ�<xp�O�4)z�����G�k�����i�"��J�wʁ��\��G�@�q���馛���������u��e�~�r��	�     .׶��A
0�͛���J�H�VbĈQT�t��x��ׅ��1�F���+w�n�޽�3��� 7s��:th����z+^|���' ��      �������ƀrr�ܹx��7�'/K��{���_�ԩSp���;�q��٨��(�4�����'M(O�6-&N�X���?����v�C��     p9ߡP���Z�����~����^,�\�ɍ4iE�o߾�I��)S�d���A��Լ����v�S�w��wMEEE      p����h[
����92��>v�ب����H���ٴ�;���;�!p���-+V���+WƨQ��нTp{��^xA�t������Ě��      �<[ɛ� �ر#{�����R�D9���������<ڛ�ʅ���8u�T �p۷oϞt��<yr6��U�3g�ğ���,8�,'O��     \@�F��>}:�-[˗/�d)�q㢲�2�I���z�8w�\ t��Y��c�w�P���F
ـ��\:����]q�K��s�=��'��ҁl���     �yǎȻ��E���H��ӂ�R�u��ls{SSS t�4�6t�ЀR&p'7lp���U�%K�Ķm����     �؉'�$�̿��+�t��;vl�J��Qj����ӟ��@��S�䆐�N�.���v[̚5�Cp��6�t�      �ST��ͱq��쩭��N�:5z���������SOŹs��3|��G�N�Nn��צ��%6oޜ=�}�K��͛����     �������ѣ�hѢl���1c���G��?��x����:���r p'7Μ9��i�����cǎ�U�      |��ٳ����yMMM�lu1bD�IL�0!�w�ީ�>R��k׮ �L'O�(uwr#ƀs�n�С1}���8qb�����5���c�Е�      |ʦV�l���˞�:L�4)k%���w7o��V�
��潀r p'7�lо</��R����QWW�gώ�Ç�?o͚56']��?      γ��XZ藚���muOK������VCCC������ ��{�@�Nnܡc����ׯϞ/��+]i�v�� �j�      >eS+\����K�,�ɓ'g������_�ҥ�\]��?��;������ �`��?~|̜93������7ް�(	w     �O�>}:�k���,_�<V�X�F��B�q��Eee�u�k>|��@�K	�)wrA��+]��nݺ�i��^WW�W��R��      �S���imm��۷gO߾}cҤI1cƌ�߿�5�k��/���� �*�
ʁ��\����k�mu�?�������      ����O�|����Z�*ƎӧO��#GFEE��s�n�;v�����������m����¹s��Z�v��455e[��H      ygS+����}�ƍ�S[[S�L��S�F�޽?�bŊ �j��H�o555�J�N.����X��޽{      ��б�=�-��K�Ƙ1cbڴi1z���w���g{;P2����R&p'� ������      �̙3t�t�t�V��Ç����c	���+W��R�vJ���\� ��~      p�������/��B,\�0���bӦMP*�P��䂀 �Tccc      ���@ר���u��@)�n@���w �R�      ��	 p!��:�;����  ��     �< p!��:�;����  jmm      Dl �żP��䂀 �Tsss      ��[ �bwJ���\�� ���     ����&ߛ  �S��䂃 p)�      6 �rnw��	�� p)�      �3 .���P���� p)�      �3 .���P���BEEE  \��     �� ���:�;�PYY  �~      `C+ p9p�:�;� ` .��      ��V �rwJ���\� ����
     ��� ��~@���w �R       ��Z[[J���\� ���     @S \���N�N.� �K9�     �� ����R'p'�u� \�{��     Pt6 �R�(u�`rA� \��     �� ���J���\� ����     ��� ��~@���w �R�      l �媪�J���\� ��~      ѭ�< ����R��\� J�H�      "��� �B�KJ���\�ѣG  ��ٳg      p~1P�����  ���R'p'z��  m�      |*Elw ����R'p'��4q���  w     �O����ٳ ��)uwr���"z��gΜ	  �;     ��Dl �����J����H!�� H��      �	��y7��	���Z�6�      >e9 p!]�N�Nn8� m�      |J� \HWA���}�� ��_�~     �y"6 �B��(uwrC� �1�     �) p!��:�;�!d �|     ��� hӭ[��޽{@)��B6 ���7     �O���+  ���;�!d �|     �TMMM  $nv���! ЦO�>     �y�
 �M���J�����. ��I����      ༾}� @⽀r p'7R�^YY--- נA�     �O�� ��^@9��)nO����� (.�;     ��Ҧ֊��hmm ��lp��ɕ�
����      ����޽{Ǚ3g (6�)wr%m۷o ����      K1�� ���r p'Wm ��     ��0 ��� @��*(wr�_� ��     ��� ����y��u�����0�0�30ð�"��b�7�D��W�TJ��m;��{�U7�][��ʹ�̫�l�i'��Ina*����2��,2���t��PYf�.��9�3�R�����|>���xO@>�SP (n���     �_�իW  ŭ[�nQSS���A ����l{M      ��i� @z?PRR����������  �O�{      ��� ���B�NAi�ںq��  ���\      vM� x?@��Sp���#p�"%p     �5[ ��w
N
����? P|�      �VYY555�y��  ����|!p��� (NMMM     ����B� �K_I��Sp��� @q�>      �ͥ���V�
 �8	��w
�� �SUUU���      ��w �8UTTDMMM@>�Spz�oݺ5 ��a�     �[3� �WZ�VRR����ܷo�xꩧ (���      ޜ� ���\�'w
R��*p��b�;     �[K������  ����|"p� ��
 �ǅ     �[�������ظqc  �EWA>�S���� (.��      o/�@�18�|"p� 4( ��&����      o-Mo}�� (�������/�����,tkii	 ��80      x{)p �KCCC�����;+Mq�@q�     ��; ������;+�n<�@  �O�     �{R�VRR��� �;�F�N��@�H;�      ��z����/ P����;k��� �����ݻw      �{R�&p��ap �F�N��իW���EKKK  �k�С�6�      ���w�} ���J��;w
Z
�V�X @�J�{      v�)� P<�y��@����&p��'p     �3w (�7w
�� 
[Za�|     �gjjj���.ZZZ (lw����6dȐ(--��;w Px���UUU     ��IM��~��  
����#�;�{��1`��X�fM  ��E     ��I�Y� P��������|#p���9R� *��     �sÆ ���m%%%�F�N�K��w� @�5jT      ������s��  
S
�!	�)x)pO+�Z[[ (������      칊���߿�]�6 ��d�����WSS}���u�� P8Lo     �7i��� 
S<dȐ�|$p�(�)�w (,��     ��1bD�� ��������H�NQH^�_ P8�      ��� (\���|%p�(�3&�n���5 ��WWW��4     `����;;^|��  
��l�3�;Ea�������X�fM  �o�ر     ��K�� 
���|&p�h�)�w (w     �����˗ P8���uuu�J�N�H!��� @~+))�ѣG      ��tW (<���;�;EcĈQ^^۷o  577GMMM      ���	�--- ����? �	�))nO��ʕ+ �_iW      �Ϙ1c�W��U  ����$F��������� ϥ�9      �G� �c��ѳgπ|&p��p�q�7 ��z��Ç      �O�A7M{mmm  ���k�������hjj��> ��������      ��&���v��  ���B p��L�81~� �&L�      ��4�]� ����<F������	� ����f�     h)p���� �_#F���ݻ�;�;E'�N����-[� �?����     @�5jT���#^}��  �S �@�N�i����_�: ��1q��      �c���Ř1c���  ?	�)w���,p�<���      t��	� ?���/���P��q��EEEElݺ5 ��7hРhhh      :N
�KJJ���5 ��bz;�D�NQ�޽{�[u ���v     ��WSSC��'�x" ��"p���)Z)��@~8蠃     ��7q�D�; 䙪��>|x@��S��Yyyyl߾= ��5`���۷o      �����[n�% ��q�DYYY@��S�***bܸq���. �ܕn�     �9����_�~�nݺ  򃶂B#p��r�!w �qS�L	      :O��~�� ��*++c̘1�D�NQK�r���#^}��  r�СC�O�>     @��@��0aB����;E-����}��� 䞴�
      ����9B�~��  r[Z��F�Nћ2e�� rPIIIL�4)      �|tP�v�m ��ݻǸq�
����7f̘����M�6 �;F�uuu     @�K;�
� �p�QQQPh�������?�i  �c�ԩ     @�8p`���?�}��  rӔ)S
����a�&p��V|��     @�I���� �{���b�ر�H��k��1hРx�� �z�'O��     @KSao���hmm  ����[70��o6���ӧ� G��U      �Z1t��x�' �-i�(Tw�?i����Ŏ; �:MMM1lذ      �륞B� ����>F�P������������ t���JIII      ����3m�4mM�o0c��; t�����"     �ܐN�81��  r���B'p�7=zt455���? @�;�����.      �i^�; 䆑#GF߾}
��� m�q���M7� @�{�;�      �q��E}}}lܸ1 ����A����8����[o��۷ �yc���      rKiiiL�2%n��  �NEEE|���N����:&M�˗/ ����i7      rOx��Gkkk  ]c���QYYP��)��@�)//��     @kjj�Q�F����  ��GP�Æ�!C���ի �xiK˴�
      �+Euw ����Y��@�o��|g|��_ ���.      ������hii	 �s͜93�X��ML�<9n��fe ��ƌ��2      ���������G?�Q  ����29䐀b!p�7�.���Z��zk  ��v     ���Z���Ǳs��  :ǴiӲ�����B�(�����ؾ}{  �O�>1a       ?���g�w���  :Gj����-���Ĕ)S⮻�
 �����%%%     @�H�x� �9ƌ(&wx�gώ��;Z[[ h?���1}��       ��=:���c�ڵ t�#�<2����m455Ł+V� �������       ��)��^{m  �O�>1~���b#p�����w hG)l�9sf      ���N���rKlڴ) ��������;�!C�ĨQ���G `�͘1#���     ��ԭ[�����  �_UUUz��H��)Mq���+++�V     ��Ҏ���~{l߾= ����UTT#�;즱c����c͚5 콴]e�^�     ��V[[�M���/~ @�I;�H1��n*))��s��W���  �Niii�+
      �a���q�w�Ν; hӧO��={+�;�<0���c�ڵ �iӦESSS      P����{�7 �}��}���L�{ Mq�7o�)� �Lo     (L�z׻ⷿ�m��� �o�±>}�3�;�!S�`�L�2��v     ��:�ѣG�ʕ+ �7�sL@���JS��ΝW\qE  �'Mo�3gN      P��=�X�; �������������A�5k� ���M�fz;     @>|x�5*}��  ����'w�i������K_�R  o�[�n��'      �4��s��\  {nܸqق1@�{-mb�1 ��#�8"     �:
- ����/���K.�$ �]����w��]     @qH;�
�`ό;6F����a��@&L�>�`  ��#�����      �8�=:F��=�X  �g޼y����Q����CEkkk  Q]]�sL      P\�?����K x{'N̆�!p�}����zh�}�� �EZ]ܣG�      ���Ho	��� ��JJJ���~w M���㎋�����u��  "�#�      �S����CEkkk  �v�!�����kwhuuuq��G�~��  "N<�����[M     �b5`���<yr��7�	 ��ű���SA;�={v�u�]�q�� �b6jԨ8��     ��6��X�bE�ر# ��v�a�E�>}�{wh'ݻw�VS]{� Ū��$.\      ����~x���? �/***b�ܹ���ѡ��]�=��� �(�      �̛7/��x��W ��c�9&����5�;�����X�hQ\r�%��� PL*++�m&     �MMMM��]o�9 ������>:�7'p�v6lذ�:uj,_�< �����={      �ёG���/�^ (vix`EEE oN�`��q����^��ѯ_��9sf      ���֭[w�qq�UW ��ƴi�xkw� ���1gΜ�馛 ��I'�eee      �2y����OO>�d @�:�����$��&p���׺��cݺu �,݌;vl      ��I1ߢE��3��L��� �I�&�������CISl/^����\�P�*++���      �vӧO���+ �����ǂ�=w�@#G�ta@A;��㣮�.      `w��K+V��-[� �9s�D�޽�=w�`i��<�7o ($C��#�8"      `w���ļy����n @1hhh���>:��'p�V]].����: �P���Ʃ���}     �=1k֬���c�ڵ ���O���� v��:�ԩS�W��U<��# �ਣ���      �4DiѢEq饗Fkkk @�?~|L�81�=#p�NPRR��vZ�˿�Klݺ5  ����Ҷ�      ��F��vX�y� ��{��ق.`�	ܡ����;�ϟ7�pC @�J���8㌨��      �'�pB����y�� �Bs�q�eC�='p�N4k֬����� �G3gΌ�#G      ����X�pa\}�� ����9���#p�N���.Y�$>��O���� �I�n$      �^�M�˗/��+W ��	.^�8����;w�dMMM��w�;n�� �|�v�UYY      О���d��m� �����aÆ�����:�x���� �3f̈q��      ��>}��q�7�xc @>�ݻw̟??�}#p�.PZZg�}v���klٲ%  �544Ă      :ʑG+V���<  ���Ē%K���"�}#p�.R__��̮�� �\ն(���2      ���(��N�O~�}�� �|3cƌ3fL �N�]�����S��=�� ���̙Æ      �hMMM1o޼����� �|RWW�| �C�]lѢE�jժذaC @.4hP�     @g9�cbŊ�z�� �|�v!Y�dITUU�>���z��g�uV\z饱s�� �\PQQK�.����      ��RZZ�=������k�� ��f̘�Ǐ���!><�����   �r�)��      ��c��o}+  �544Ăh_w�s�΍������O t�I�&����      �J����#�Ľ�� ��Ү#g�}vTVVо�#�Nv���'m�@�I+��,Y      ��/^�V���7 �9s�İa�hw�!)*<���k�	 �lm��z��      �ժ�����O�/|���� �+��@��C��>}z���=�� Й�?�x+�     �)cƌ���:*~� 䂊��l�`YYY C�9hɒ%�nݺx�� :�ĉ�裏      �5���φ�Y�& ����=�� :��rPyyy��}�O}�S��+� t�޽{�g�%%%      ��[�n٤�O�ӱm۶ ��2y��6mZ K�9*ņ�sN|�_��;w t��EU���      ��_�~�`������ �cɒ%t<�;�1c�Ĝ9s�?�A @G8�SbРA      ���xG<����� t���HX[YY@��C��7o^<��S��� ���;,?��      �|PRRg�yf|�ӟ�^x! ���x�1x�� :��r\�8;묳�3��L�_�> �=6,���      䓪��x������gc۶m m���1s�� :����/ζn� �/jkk��s�Ͷ�     �|�����zj|��_ �HMMM�dɒ :��	�Ā��UW] ����ʲ����>       _M�:5�x���� �***������t.�;�C9$�8��; �ƢE�b�ȑ      ���O�5k�ĪU� ���ŋ���t>�;䙅Ƴ�>�<�H ���5kV̘1#      �t��-����O}*ZZZ ��QG��t�;䙲��8��ⳟ�l���7n\�t�I      ����6�=�������رcG ��=zt,X� ��#p�<TYY\pA�ۿ�[l޼9 ����/�9�(--      (4Ç�N8!���� �޽{�ҥK5���m�.��2+�xS��_�(�G�      ���#��5k�į~�� ��Q^^�}�{���&��%p�<6bĈX�xq\s�5 +]x-[�,      
ݢE���}�ڵ {���$N?��<xp ]O�yn�����K/����� �6��묳Ί�C�      ����x������g���% `w͛7/9� r��
@:�n޼9~�� $'�tR|��      Ť��.�?�����Kc۶m ogҤI1w�� r��
��'�7n���? (n�gώw��      �h���q�gƕW^��� ofȐ!q�gDIII �C����4�.]�]vY<��@qJ�e��      �,�v|��ƭ�� �+�{��.� �w�@n�CI'ڴ�ֿ������? �1c�XU      �gΜ9�~��X�|y �UUUŲeˢ��6��#p�SSS����K/�6 �aذaq�y�E�n��     @�C�v�i�y��x�� ��V���������PP����㢋.�"���� ��80����GEEE       QVV�{n|�s����~: (nm��F�@��C�jll�}�CY�iӦ �0555�>��l�,      ��UVVf��.��X�~} P�.\S�N �	ܡ�����/�V!oٲ% (,}��/�8jkk      xs555ٮ�)r߼ys P|fΜGuT �O����9�@���?[�n 
C}}}\t�Eѳg�       �^ �lٲ�����^ �G��~�)���P��~\~��}��  ���)n�ݻw       �oȐ!�| ���/P$<��8�3���$�� p�"1z��,r��;v� �SUUU\x�ѷo�       ���������j( 
ۘ1c�sΉ��� ����رcc�ҥq�W�Ν;��RYY�Mn8p`       {�-x��+4 �mAS�nRY�7��B�9蠃���O�k���@Iq{�*q���      �<0�8㌸�ꫣ��5 (C��:���� ���дiӲUi_������_ r[UUU����aÆ      �~�N����^{���@477g�E&�'�;�ɓ'g'�~���}��  7����E]�]|      �o�����k��7� �>}�ą^����/�;����g۰|��_�.� �-={�������      �q���wƖ-[����~ ��z��u����7�;�Q�F�?��������J �z�>766   �-�رc��}�{���  @~�7o^l߾=~�� ����..��⬷ ���!C�d+׾��/��/� t��}�f�����  @�Ν;�)z)"O1y�ұu���{���j�1}���g?���?���f?�>�}�~����+�L:v���RRR��<�����]}��������O����ʲ�����\^^���+**������ا寧m�Zڞ9}���
   �����]��v�m@~HQ{�,(w 3hР�������?---@�8p`\x�QSS   �b۶m�y��?��)VOQz:R�����������):o;
͞��)�o���t�ħ�-�O1|����6��G�QYY�}La|:z�����  ���p�	����o�9 �m)j��?(n���3�g������q�e�ņ�Εv���>��,  �Ui�?��Y���+�d��H�-To��S��>���s���.$H�wW����I��c[���t��b����/�ӑ�  ��fϞ�����|ǵ-@�J�[��^WW@a�%�d��⋳�}���@�5jT\p���  �Ζ"��7f��7mڔ}�"�4a�m��`�]i�}H��ۤߛ��65>M�O�H���t�§k����,�����~  �+̜93[�{�u׹�1��/�0���;�wz��Mr����㩧�
 :�Ag�}v�0  �=�����HS�����i�)H��UڦƧ�����V�b�tݜ�����)�Oӹ��� ��2cƌ��ꫯ���F�˖-�& �I��Rz8�&����g���@ǘ5kV�|����  `w�M]O�_z�l�z�����q�6�7���w<���J���"�4>�'555ّ�u655Euuu   �C9$�ָ��+�]� �:�F��.���(pw�M������}q�-��m�� ���ϝ;7�=��   �[)�}��c���Y̛&��p�m�q���ߋt��'iǂ�������S߽{���g������eccc���  ���8qb�w�y�|E��E&L��}�{�!@a�o)m�{�	'dx����lR ��[�nq��ǔ)S  (^)T߰aC��	�i{[��A9�����?�n�����#�<��_�L������uuuY ��ܜ��  @q7n\\x�q��g�� t�ɓ'�Yg��ݿ
���-3f�Ȧ]u�U�m۶ `龜�iw��e  P�^~��l
{���D��y
kS��	���o����Y����{���o߾��  ��0r�ȸ袋�K_�R�� ����ŋg�Z�� pv���G���i� {&톱lٲ��7  P8R��nݺ,do�طnݚM��C�x��==\M�{eee���D}}}455e���  Px���ǲ���� :��ٳ��㏏��� ����#i+ޏ~���E�ڵk��3|��8���  @~j�ƞ\��5}�B���-�Ȑ��#-tI�N|���{m����o�l�{�>}b���Y  �4�*	��W��=�X о�@�E��G@��{,=����?W^ye<����[�>}z�UV�n�z @>x�����"���]
ٷmۖ� {ꍓ�7l��?�x�}���C�4ݽ��*jkk��}����W   ?TWW�E]���7�7��M �>***b�ҥ1q�� ���
�+i�������w◿�e ��҃�M�1�  @nI�z�ľnݺ,dO�_}��,d��u(E��H�C�W�ξ��'���)|�ٳg444D������>  �ܓ�\�}���{��o�= �7i�\C�	�x	܁��.�N=��l;���ر# ��4�!�&;vl   ]+E�)f_�vm����iӦؾ}{���@�I�{Zp�����O<��雷��!occc6�}РAv� �PRR,��}��u�]�����K���-[�{�����	�3fdo.��կf��]�q�v�hjj
  �s������3�ĳ�>�MD~�W���bv��;6lȎ�+Wf_K�{Zh��E�E�555  t��;,z���i�& v_ x��F�=@����Ç�'>��"��'��b5q��l����   :N�p�~��x����---ٴ��u�b�v������W��_���QZZ�ݛ�������)~O_  :֘1c������/����Ҁ�E�EYYY $w�ݤ�%_|q|��ߎ��+ �Iz@<��8�c�- ���&�=��ӱnݺظqc6�=M1`��b�-[�dG��"I�+***���6��{���!z ����k�E�k׮ v-ݗ8餓b֬Y�Fw�]����i���F��믿>�n� �.m�����i  ��IQ�3�<�=�}�bӦM�}��hmm �^zM�ґv�X�re��{�)zoll�"��  �������h|�[ߊ�˗ ���:�9���Kw�CL�6-W\qE6]�P�92���ٳg   {��_�5k����?---ٴa1;@�H��iG�6dG�������l�Φ��>|x��  �siA�g�����[n�%[�@Dsss�w�y��� �"p:L�~�������7��{��B�&��-�.\eee  �������g��B�W^yŃ]��^���u:����+�{��_6�2�9C���ݻ  ���s�ٳgg1�UW]���(f�'O��N;-***��܁�&����&L�뮻.����Բ�O?={m  v-��<�L�]�6�ξiӦx���Mg�C�����cv�^�:����֭[���fS��i�;  �k�ƍˆ~�+_�u��@�I��ϟ�sL���܁N1mڴ<xp|�k_�n�ѣGǙg��m�  �EKKK�Z�*���H��
ێ;⥗^ʎ�+Wf�{��My4hP6̔w  �i��'>�����w�uW �4H�Ί�c������_�~�},n����; ����s�̉y��YI  ���_�'�x"�8����۷{�P��[�lɎ��i���Q^^�MyO������a6  ��>���N�Q�Fŷ����
@!9rd,]�� A`�܁N�.�N>��1bDv��v ����8��c�С  ��瞋'�|2��&����� o%�:iAT:~��(++�"�4�r����=  (VӦM�����W\6l�B��̚5+.\�� �w�KL�4)[�w�5��C= �*�XZ�hQTVV  ��;w��ի㩧��^x!^~��l2/ �tٱcGlܸ1;y��Awuuu���7���=i=  (������o|#x�� (UUUq�g� {C�t��5�e���;�o�1�n� �"M[�d��-  ��k�����O?�t6e7�&h���sMZD���gG
�{���{�����l�{�ne P�Ң���??k'n��l'$�|6t��X�ti444��rW�R�Ō3bĈq��Wg��ڸq����O��={  �m۶ţ�>�]����K�� ��R�Y�c͚5�|��lW����6lX6�҄w  
Q[;�y~�k_�g�}6 �Mz-�5kV,\�0���`_܁�Я_���G>?�я��?�q�U-@gK[d�x�1}��  �B�s��X�zu�Z�*^x�x��W r]
��9+�0����<M��۷o�92���  
I������x�|��q�w@�������>;�^hw g��{�{lL�4)�����;@g?~|�z��E  ��{.{�X�n]����Y$ �,���9���ώ4�}����>}�Ę1c�w��  ����<N>��l����_���J ��z-^�8[��^�@�I+��4����gq�-��&�Pij�	'��m�  ����%�׮]��9Mm�B��u�6mʎ��gϞ1`��;vlv�  ���ɓcԨQq��ƃ> ����2.\�� :���I�AđG�=���7��m����M�SN9%jjj  ��k����|O=�T��⋱}�� �b����7f�C=�M�L��<8�"�{��  ����6.������;��o��[�@.H�L�y���� A��~��Ň?���{�������v����-����  �;vd�W�^��h�[K��֯_���{o6ѽO�>1bĈl�;  䃒��l:rZ�y��Wg�� �JZL>��lpiz}�(w �7CӦM˦��t�M�|�� �iw��3gf[  ����%��Ӕ�M�6Ekkk  {.�C� �'�|2;��ʲi�)tOCҶ�  �������G�g?�Y|�{�3� �tÆ��N;-X
���@�H��6ӧO�뮻.��� �]��SO=5ے  r�Ν;�)\�V�ʮ{�m�&j�����ƍ�㡇���7���  �4�+MM�8qb\{��裏@GKSۏ=��8�裳�!�� p���������w�qG���?�*xK���1w�ܘ5k�-  r�k��+W�����	����q:�#�C����&Ӎ92�w�  �KҢ�}�Cq�wƍ7ި� :̈#���MMMЙ�@^J+gϞS�L�[n�%�/_ o�Dv�a1���o��  r�s�=�E��֭�W_}5 �ܑvTy�����{�=zD���c�رѫW�  �\PRR3f̈ѣG���_������TUUł��"�� t6�;����3�<3=�и���g��Q���;}������Ir��@¾( ⾡�(�-ڷ��u{z��{k��<�5U��>������wf����]^���Kk7����l�����dO���"\�n[� Y^/�S�sN�]b��������]���/bٲe  S���H�2��ѣq� `�K;���Ç�TTT��ʕ+�;�c   7]js������O���������C<��C���Q__ 7��;0#������x�w�W^�7��g������<_l �ͦ� f����hooϓ������˗�]wݕ��  �f���{c͚5���/��o��k|)s�w�w��fpf�Ԝ�e˖x����^�m۶��̗n��_�U���?����  ����ɓq���8w�\ 0s��Pooo�۷/O�X�%K��}�ݗw �-�7M;]�_�>������� �&�,�y�x��d.�)C��q�[jp~����׿�u�޽��d���Л6m������5  7���D?~<:�C�Z��522��Z[[s!KKKKn�[�ti  ���z���?���Ď;b�֭��� �w���?��X�hQ L%����`���������/⥗^�#G�03���Ń>���.  ��R�=]k<x0:::,� �&������ӧ�{SSS�~��  7B���aÆ��{����w�ɟk$)W������{�7 �"w`ƻ��������y���q�ĉ ���z����+W�  �QR#�}������^�v ���^��������X�vm��:�P  �S]]]����a�_��q��� f����x��b˖-yA6�T�;0k�P���_�+v��������`����[�g?�Y�[�.  �FH[7��q������ �*5fvvv�����>����X�jU�y�Q,  ��T �?����O>�$����3!0{�]}�������FCCC Lu����N�z衸�����W_}�ELq��rK������y  p�uww��Z[[��ŋ p��a��0�q�ݻ77k.[�,o_[[  p=��ʹ���wߍ������ f�T
���ݿ�ל Ӆ�;0+�����?7n�?�0^y���0Ť��-փ>��  ��r�,;u�T��� �����i�����s�=5�����  L����x���G�!���{/����Y�,Y���w�uW L7������6l�[��޽;~��Ĺs��y�/_?��O� �������>�� L9)��O>���<W��iS� ��T__���>�l�������>&&&�ޚ��r��M��P(�t$�P�B�=�PԦ�������8�W�������7�  �zHA�O>�D� �V�¼49�~��w��M  ����������ǹ�=�����2gΜ�`%��\YY әO� �"�S�6��Ç㷿�m? �G�o.m��V�z�  �mdd$���G����^7� �i-��|��Ǳw��ܶy���wܡ� �I�dɒ������Yگ��8t�P S_]]]<��39�^UU 3��;�7X�fM��G��믿�oB��H+�7nܘ/�,X  0�FGGs�i����  3M��:��?����裏���1֮]��v��;  ?X�}��������lꩧ�駟���� �I��E����������.�{ｼ%,�ݥ-�7oޜ/���X  0Y&&&�/�����7���"�uvv����cǎ9�~��w�1 ��J1`*�x���a�lfw�k4������=�\n�y��7��ٳ|��˗Ǐ~��ذaCno ����P{
u��  �ٕ������������sO,^�8  ��J�������Y�?��?������R�`
�?��Q]] 3��;�w�N�x�x��������o�>��GR�������  L����ػwo���� |����8}�t��Y݊+���"  ��m������?�{�7b�Ν>�� �r���?�y�b� ���;��TVV��w_����x��r+N___�l�Z����{,���  &C�ٳ'Z[[cxx8  �v���q�ȑ<i��U�V����n ��-[�,���/���ױm۶��H���J��=��3��#�D�P��ħV �`޼y���?�i\���C�iug�H7��b��Zxݺuy  �P��)mw|������u� 0	��>�;��϶��޸��[  ���*��_�"g%R!�R@��R�⮻�-[��w� ���;�$J!߇~8OWWWގ�w��]ttt�D�/��7jk `R�<y2>��hoo��1 �u��ϱS����}��ʡw  �.���ڵ+�x�hkk�ڥ������'?�I,Y�$ f;w�뤱�1�t>��q�������w�-�^]]]��jӦM�|��  ����ߟw�jmm����  ��ˋ�TWWǚ5kr�{�X  �V)��aÆ<iWƷ�z+>��S%�455œO>�?�x�c p��;�u��Z�n]�����sn!����������Aeee��*}q�}��&  ����F_|񅭋 ���������yZjsO�m�~��  �ŕ�Dwww�ر#�~���/Y�'�x"x��(
��I��@)$��xM��}�Q�ܹ3�=�����$������֞ښ���  &CjM�ϝ;�Z `�J�i)��}�����c��9x���  p�Ңɟ��'��3�䅔��=���\�٨��!6n��7o���� �L��&����[�I7	҅\
x���Y���S������O `2����ȷ��-��� ��#���>}:OMMM�^�:�X,  �Ej�N�i�����C^L�>7��,�ݿ����������o'�0466�m��������w
�sݥ�P�b���{�'���  &Kڱj�޽q�  `��E-����m�i��e˖  \��;��~���������������H�L�p��x��cӦM��� |7� SLڎ(mE�fxx8��S�{
���;L����JS{
�WUU  L����سgO�kk ��.]��w'}��7���2V�\�<�Vw  �YYYY�q�y����s��������|��9s������Q��
��O�`
K��+[t����]9r$>���܎s�ԩ�k������[sC{�J  \�� f����8|�p�[�;  �G]]]<��Sy�B��螚�O�80���)׳aÆ\4XQ!�	0|7�&R@���n����<����СC�����{�����?����ijkk  &��v  ��� �dhll���~:O[[[�ڵ+>��hoo�
�5�]wݕ��w�}�y �w�i���>�(�I7R���r�=5�\�x1�]�E�ڵk�"��*���9  �z�� �_�ǭ�>�`,_�<  �H;����~�O��A���}kkk����r��ӹ������: �~�f�����u[�l�x��/��{{{��%5�_	��cz  ד�v  ��+��۶m�� ��dɒ<���Ν�ݻw�'�|ǎ��0��{��-�h0]� pc��@_�?��S�����8q�D��I�S��CUUU���n��I�v�  �(�� �_muoii�͇.  ���y�O��<i����}
����/^��{o�իW� 7��;�,���M�N��t#!��Ӷ]'O�̏Ϝ9����͕��R�=mכ��[oͫ��B  �����w�ؑ�\'  0�R�f{{{���Q]]�=x��� �����œi�g�i��������?����_2gΜX�n]nh�뮻r���O�`�J�&���i��ӧO��4)�����/��mjjʫ�.]���)؞V��� �͒�v��n�  p�ŧ�~�}�Y��tÆ���  �}����r����/����{
�wuu�[EEE�Y�&��<+V���0	�pU:�O'�i�*m�B.W�Y������٩����i��4�-ʓ��͚���  ��mbb"��I��t�  7ZZ\�>~��s�}����Y5  |W�������I����ȑ#9�~��ᜃ`f+��p�J�=S���M��o���J[Ħ���I!�+��4.\������3+�
�EUccc477�c
�/X� �׬� `*Ja��;w������=  LiWѷ�z��N��<�]/ ����C=�'I��ʡ��G�ƩS�|V:ͥ���zk�Z�*�\V�\��^|��{K7�4��9ccc9�~%����J�nN\y�&�j�T>���������;�ܹscΜ9W�ijj�Gv  ��Ԍ�k׮���ٰ( ��itt48�;bnذ!�U  `���G}4O2<<���q�رxO� )��Ԕ�멝=گ���ϟ L� \7�B"5���9�~�&�䇆�b||���tA��U��k�&կ���ɍ�W�UUUy;������+�^ ��$�?�ݻ7o��έ `�H�2�"�_|1�ׯ_+V�  �l)+�v��<W�C:M��'N��ٳg���`)ױt���Ⱦdɒ���[n��0C����q%\~��x  �ۥ�v�ܙ��l� �t�v}뭷���2V�^�<�Hޑ  ���cX�fM�+R1ߙ3gr���Ǵý�����-�b�r�%�]�   f�tCe׮]����
  3���h8p <��.6l���  p#������R�=���?>O{{�������ei���������㦦�(++ f7w   �"5��޽;}ҍ  ���bδ���_�y��Ń>+V�  �R�}�ʕy�XZ��
I�����4�q
��݊Ҏ��]
�ϙ3'�9z:���tL��t�;wn �_"�   0ͥ#��=�W���  �F)��[oE�X�;�3���(
  SA
~�݇�|���n___�������ϡ����̏�1=ʏ��I�'###1666)������\���:�s��~z�����D]]]>���_�\O� ~(w   �i*x>����X��+ �����?�8>��X�fM�_�>**� `�+//ϭ�i�/_����|O�}&�%�_��W� {�g ���'9    ��ٳgc�Νy;[�v  ��R{��СC�hѢشiSn� ��L�: 3��;   �4q�ر�裏�ִ  ��I�iף�[�Fssslܸ1�ϟ    LM�    SX
��ݻ7>���  �����W^y%����G�e˖    S��;   �422���:ccc  L�K�.Eooo���Q]]�֭���?    ��   �����رcG?~<��  ����P|��Ǳo߾X�zunu/
   ��#�   0\�p!v���O�΍�  ��3::�;(�X�"6lؐ��   ���   n����������'  ��+�vSJ��/��7F}}}    p��   �ǎ������   ����R�]��_����x�Ǣ��9    ���   n��ƞ={��ŋ  Lm)����/��r466ƦM�b���   ��#�   p� ��������J����ƍc���   ��p   ��R�}׮]144  ����{{{㷿�m444�   \�    �lbb"����}�Y���  0��믿uuu�aÆX�lY    ��	�   L�+��O?�4FGG  ��R�{l۶-jjjb����jժ    ��p   ��R����>�������X   �K
���~��عsg<��ñz��    �p   ��R���?��;  ���P���{9�~�}�ŝw�    \;w   ��hdd$7�<x�jc{YYY   \��҂ؽ{��{
�   ���   �Q
�l߾=�9��  �&�:��?�����<�֭    ���;   ��Ha��ؾo߾���   �E
��ر#7��_�>V�^    �)w   �o���)|�F�  �CCC����Ǯ]���G�[n�%    ��    �g�}�w��-�   �-��}�ݼ[�ƍcɒ%   ��;   ��8p 7)��	  �����o��f�����?.   ��L�   ��/���;w���`   �H�.]�A��^{-cӦM���    ���;   0��8q"�o�}}}  p�uuu�+��MMM��}޼y   0��   �R[[[|����ӓ�  ��t�������ob���y�樫�   ��@�   �U�������}�   Lu��^�E��F����    ���  �Y���#��Qc;  0��k�3g�į~��X�ti<��Q,   `&p   f����x��w���-   ��tO�6���/cժU��c�E�P   ��D�   �������C|��� �%]�9r$Z[[��;�3    f
w   `�ٳgO�ݻ7��  f�t���Ƨ�~7n�+V   �t'�   ���}ǎ144   �E�z�w���.6o�---   0]	�   ���ӧ��ދ���   ��.]�����ꫯ�{
���;   �t#�   L[������o����  ��A����x�b�ҥ��OD�X   ��B�   �v���rc��'rx  ��K�Jmmm�����w�>�`
�    ���  �icbb"v����y~  �_���������z(n���    ���  �i��>�]�v���X   �݌���|�|�I<���x��    ���  �)�ȑ#�}��
   ~����x��ף��16o����   ��D�   ��.\�۶m����   `ruuu�o~�X�|ynt/�   0�   S���H����q���   ��:y�d��?�c�}��q���   ��&�   L{�쉏?�8���  �#]��ݻ7<�6m�e˖   ��"�   �t�O��w�y'  ��chh(�m������SOE]]]    �h�   �M��ߟ���Ν�K�.   7_ggg����bŊؼys
�    �Q�  �nbb"v�����l  ��ҵZkkk�򗿌����ڵk   �Fp   n��?�<v�����  �Ԗ�ݶo��~�insoii	   ��I�   �!.\�o��Vtww   �K��꫱hѢx��'�X,   �� �   \W###���Ɖ'��   LO��̙3�����w��ׯ   ��&�   \7{�쉏?�8���  ��abb"���G���{,�/_    �E�   �tmmm���.  ��ihh(�z�hll���z*���   ��p   &M
7���q���   `v��ꊗ^z)V�Z���B    |_�   ��سgO��U=   �˥K��ȑ#yG��<�-[    ߇�;   ������%���@   0�Ƕmۢ��9�l����   �]�   ����X�������   �U����u�ָ����{�   �k%�   |g��y�ر#��  �ϙ���={������'�����    �6�   �5����[�www ���(�]��,.Ey���𤋮����ңKQ(���2��~OMMM��}��先�?�ߚ�T�.]��|hh0.��/���h��\�M�cc1<2W�9���c� �����x��WcѢE9�^,   ���   �*�������-� 7B
�� z��cDMU1j�����*��������X�������ʊ�����b1��K�����beeT/?���,���4�QV������(��,��f�ti"�FF�>�A��O��������q������X����p������|�q�}�C�������qpp(.�fpx$�t�zKגgΜ��[���?k׮   �?G�   ���;��^��� |_��2�����p9�^S,Ɯ9�QW[uu�cMm���Du���zu�Kϋ��L�Sz^(��l������W|��dI�F��r ~xx$7��c鵡��.�P����?0�}��S������o |ccc�}��طo_lٲ%���   ��  �?��ŋ��o���� ��Ԭ^,/��,*J�k�����>�룮�&���Ŝ�ڨ)=����buMT��U�c��:7�s�
��.�{J�]������P^,�;���`i��b�_����x1zK_��틾�{�@���/��R�Z�*{���    q�    �{��ɓ]�}�eQ����XQ�ڪb4��ż��Q?gN�ח�nN���Eu����%-R�-��H3����?>1C�����w9��ן���7:�����?�zz�b�= �|i�ӑ#G��ɓ��OĲe�   @�   ���ٳ��[o��U f�BYD��<������be4ϛ��^���������S��)�\QY��򨫛�g�_x���H���F�Ł��닞��|����=�q��+�GF��a��}۶m���[�l����    f/w    ���r��ĉ��V^V��<5�Q_SM�Rp}^�K����������!���(+�����X��������DoOO���EWww\(M�����s��14< L/����[�n�x ���    f'w   ��Z[[�wމ�Q-� �EE�J��<���PW-�͹����1�4̍چ����vf����<-��_����N�����t���������	 ������裏�������F}}}    ���;   �Ri������ L-eeeQU��W����ǂbol����b�ܹ1�a^�WVU�uUUձpѢ<lhh0߻.tEǅ�����;�t��� n����x饗��;����   0{�  �,���o�ccc�͓zի*ʣ����幕}������%�����)7��k�U5�L���X�(͟���GggG�?��:���s��8���.]
 n��}w߾}q�رx�駣��)   ��O�   f����x��7�ܹsZ 7P��,��s������X�2?̟s���~^c4�+�P(��)VU��%K�|U
�w]茎��8{�|�>{.N�k����w^p]��/��W���{�t�T   `�p  �Y�O>��>�(����룼P��QWY5��+VDKsS,X� �5��ܦ�h(M]}}��	f�t���/�s�W^����=5����S9�~.�/��;��:r�H���ŏ~��X�xq    3��;   �p�����oDggg 0y*R���<�)VDS}],Y�(���4�DCSS���f�bUu,]�2��J�.��F���ўB���ƉSg�����{�!����5�ҥK㩧���   3�;+   0��ٳ'���D ��e9�>�X���X��%ZZ�������9j��@RV�5�an�[V������pt�?gϵ��3g�ę�q��#F���%�w�k��g�&��>�x�X�lY    3��;   �@]]]���G___ p�
eeQ]Q�f�,����X���Fc˂<��GyEe |W�UU�xي<|����htu���z?{6�N��ֳ�h4ƅ������ضm[,X� �~��(�   L�   0�|����'�h�)�^[Y����^U��2�9���7�,��M�R��~����EK��u�����;ݝq�T[�:s6ZO��g����� �����غuklذ!V�^   ��&�   3D����o���@ 𧊅�h���2�^����/\��_ifof��B��ۤ���˯ƅ�sq�̙hm;�J�����@���X��������3�<UUU   LO�   0ͥ��w�y'�;���K�B�I��U�cE4��Ăŋ�y�hZ�8�,��� �.����+n��ࣗ_����Ϟ��S��h�8q�\����D �V���������o�=   ��G�   ����������P �V兲��,�9iR;{�����/�����ļ��(+��I�����u�x����h�\舳�ڢ�d[n=�}�d<&,�f��������������Fuuu    Ӈ�;   LS۷o�}���l�����1��27�ϫM��K�)��/X�[�+�U0�TTV��.�s׃ǥү����8w&�N���'�TGg���؄�;0�uuu�/�7n�U�V   0=�  �4�nп��kq��� ����hHa�bE��sr�}��%_��/�B� |]ڹbn��<��'~Tzmhp :Μ�S�Nű�q�ԙ���q�w`f���{/��?���Q,   ���  `����O>�K�������<7�7�c^Ue�k��2̞Z��ļ���໫���e�n���Ãq��\�=}*�;G�NG��h���L���[�n�'�x"V�X   ��%�   �@������ 3͜b��v��U����e�}i�,^����QUS�Wޚ灍���{Ǚ�q�T[o='Ξ�����8:a�%0�6���~;�-[O=��]�   `�p  �).5��ڵ+&&&`&�/Vļ���[]����0wn,X�<O��e�]��#ޗ�Z�g�C�q�T[�i;G�����=2���������矏'�|2/^   ��"�   S���@�������� �Ϊ+�s�=Oue���F��e�p��XP�����Ԕ-_�6�#OF\�뉎3g�ܙSq���8}�;��Fcx�bL`z�7�x#V�X�7o��   S��;   LA��۷������BYngO���h����%KsC{
��76EY� �OZ��f��u���~=���v2N�8_k���C�72��`��t�R���Ư~��زeK455   p�	�  ���^��8w�\��0�ʢ�x��}^Ue4��y��h_�tY4-Xee1f��Xi^sK���=O��EǙ�q���8z�X����ޑ���q��688/��r�~��aÆ    n.w   �">����v`�+��E}UE��2Ԟϩo��V����ce�* �]��+�π4�=�9����q��X9v4��^������(�v�ԩx��g���>   ��C�   n����ضm[�8qBk;0eUʢ15�����TUV��ũ�}EnjolY �U�5��r�</MDwGG��:'����'�kh4���bd|" �����x饗��{���?   �O�   n��'O�[o����0����E]e!������U�Q����E�WFEe1 �Z���b�4���P���q��h=z,:�rؽw�nF�͗��ݻ7�;?��O���6   �G�   n��������_|���2*
e����4M���*��e+r�=Mm}C �d���������x��j�3�����cq��B\����p��<�����/ģ�>k׮   ��p  ����;^}�ոx�b �l����\S��U1��2�kkr�}��[��pC
�WS=���q��'���9��#�32�#�p���۷o��Ǐǖ-[J߳
   \_�   p�۷/v�ؑo���ee�PU�[���������@����b^KK��~��RW?7��}�G����8}�H?v,.E��Xt��rw�F:s�L��?�c�ϟ??   ��G�   n�h����ԩSq�$pcU�rK{
����ʊʘ�xq�/�uM���	 ����kb��uy����q��X�;g�z�sh4���b�96p�+��w�yg<���   \�   p��;w.��Ӎp�%5�7�TFSM1�UWFuuM��Y�lETTV L'��W�=�ēq���8}�h����sp4:��bd�nI�����hkk��{.���   �\�   pm߾=�������幩���"�VUFM]],�eu,�uu�,Yee� �� �L[�ty��6m�������#q*��ϵ�f����v .�  ��IDAT������կ~�6m�[n�%   ��#�   ����@޶���' �������,�P��Ҥ�{��h_��X�d�P; 3^Y�Wc˂<w=�1.��ę�c�v�p�8y2������`2���Ż�Ǐ�͛7G���   &��;   L�Ç�{����p=4TU�@{K]UeQW�KnY�V�M� �Vu�sc�����j����S�98]C��3<�X&Kkkklݺ5�}��hll   ��p  �I211۶m�7�&S�,����5��T��B!�6��M��V����� &���H\����xi"�FF�����t���/�����<^��x��cc��mtx�k�/�~��|��+�7)��GEŵ}��vq��,���ߓ~oR����g����/�^Q,�]"���+K�w**��+K���ǅ���π��a����h;�Ei�����04�����d��_~9x����{   ���  `ttt�k���ohL��Ծ��*Zj�Q^(����X�zmin�9s��R}���xdd8FGFJ3c�#9t�B�iF���|<r��ޛ�c�D��+/��BEy�U��9_���)9_����=�yeUuا���b�ZX�"��\���y�{{.�ݏ|���5<v��]���.]��w���S�{�X   �p  �h׮]�w��|#��Hm����_S�uUQY(�a�h_�f��vf��A���H��xh����/�P���3.ޫ.�߿r����TU�DUMm�X���t,��ǜ������yz�.��#����Cq��+�h�������[�n���z*�,Y   �w#�   ����H���q��� �!j+�cAm1Ω�b�,j���@{jkolY0SLL����`ib(����p�8<4�/�K����.)$�f���OZ�B�Ś�|��������{u
�פ�5QS[�)�?���)�Z�!υ��rн�ȡ���C�����266o��F�\�2�|��    ���;   |i���~;߰�>R����X����(���Ukr��y��(+���bbb"�.�������+K�����_̡�^O�0��"��/L\��򊨙3'�k뢦�.k��DUm�׎�����Բ0Ͻ��3���������1�;Gcpl" �U����^�����Q[�9   |;w   ���o�����*|gU�XPW�QSQ����޺:��,Yee���&��^�X��+=���)Ȟ����S㺟�L��c��ӝ�/�,�nW��W��7D]CC>
��li�Y��yx�Gq��8q�`�>v4���s����h��߮�t���/��͛cŊ   �e�   p�FFF��_���� �V�BY����9Ŋ(
�p��X�v],^ykn��)~SX�b_OiJ��t�-��{��f���y��ȅ�����I;o��{m}×���W�5u���=3C�P�f���#_D�r�{ϗ����؄�>�7�;��\�2�|��    ���g   pN�>o��F�����)��ESMe,����ұ��ZCSs��m]������itx8�sp�4����@�qOOne׾�]Z������?���Kǜz��C��q�c}Cng���,�-��ʓv�8u�p;�?�:�G��x��ą���m�&�����K/�s�=U��   ��p  �o�}��ؿ�����cAmUnl�,�EMݜ�Ծ�u���p�\�4�ep�;������+�z�s� ;�iaI���<,�ޑC�s�E��ƨO��ω�yM9���~ί���<Ο����Ç���@t�������?�[:oۺuk��G?��˗   �u�   �R[�?��?������T�r�}aij*
��u٪5��ۣe�2�L����ׯ��{R��+�'&&���Ǣ��B�?VUS�E͙�)�^z\?o���)��ea�{7>gO��C�Ǚұh$�ӌ��>�����x뭷bݺu�裏   �/�  ��hoo��^{-FFF���ʢ��2�V�cY�����s[��[WGyEe��511�C�}]]��}��0{O��t���h 3���`�<�O��������˶�yM�ϻ<�kL�B!�ܲ*���@�8|(��=:�{x,�/�f����8�O�����U��    �  �O�޽;�����N��H!��bynjo�-Fy�yjӽ��;Jsg�Ω�.R�=��s�sg>� djc�3�c�����|��J?�jJ?�����mj�y�[r|�P�<U5�q�=���:�������Pt|���;< ����u��زeK,\�0   `����݇wTס����M�����@�M��N��o��%\�Yy�ɻlc�m c�cS%��*H��4}Fq�QT�|?���b��،�>���&�    �7
��z{{599) x��4����v�Ô�phs[��־iK���S��/��>�^���� ��� &_�����[�wk�UM4�H}�"u��QB������^��{�ɑ{Jds�N<
�g��^�\N��v�ڥ_��W    ��p    �hffF~���� �4E}.m
x���jcuڶc��tu���
�!�Ĳ�g5,/���!����� ֝���_����з�{|>��?�jc����ُC�m����sniﲇ�(a��n]�B[B-d�Jd�0�?5��d}v߸q�^x�ꫯ��v    �jD�    P���ǟ�9�C v[��Ծ)��4�r��ұ][�w*��$ౕ��K�Z��f�5��Ѱ� P��ɤ��F�����DU��-�Vۻ�6������h��~c7�[����=2�+z��hr9�4��@U����;Ｃ?��Ojhh     Ն�;    �j
?~\���ہ*��m�Vȯ��Y�v�Rs{�N�U�\6���3���������̞�� ��:^,~�YC��~�
�[A�hCc�Ѿg��g��[��ܦ��G�nZ݁*�-�~��G��/~��{�
    �j��9    @U���Woo��� T'�ӴC�߶�{<�ڽK��(T�S>������4�`�ne_Z�g!��d�J11<d�ǂ5��44*Z�h߇c�r�\³ki�ԍ������Vw��YǠW�\����x���)     �w    @չy�>��s��@u��v��L۾s�Z;�	�U�������v�}~fھ�`J�|^ ����`��;��s+��D����ZM�ֽi:�'
GT�=j�����mvvV�����^{M�pX     T:�    ��r�����@u��v�é��Nu����<��_���ķavk��9 ���.l��1��~�j�#�56�n�f;��Ddo�aV��͟�?F�;P��鴎=����C     T2�    ����d��sssPC���`{�����hL���m�9]n�r��	�NNhvjB���P{.� `�Y;%=�ݺn���x�oP�q�bMM�54�s�hi���K��k�mu/��TN��i���Zt �2Y���}������;     ���;    ����̨�����|VC���nۭ�v����vm۵[ͭ��V�������v#���};��{H� JH6���ب=,Vy(��彾i���U��⟅5�?���ud�:��4���T"�\���@���u���kr�Y�    �<�    ����:{�,!G�
]5��j�e�|��:��Ӷ�����ʑͤ5;5���1;eڧ�˲�	 ʉu|��-�P��6ہ�ئ&; _M����O���߼Sm5^���$3�XJ+�+@�v�{��w�{$     ���;    �b�9sF���P�b>���E�.�y]S�:��S��)���f����� *�r|������n���?�Ge�U������?fR��m��LN��&�PY���;��������     ���;    ��Xx�=j���L.�Ц���{��Z;��s�
���R�Y���531nߧ�	 �O&����=,�áh}�wB�V�R�F�
G�_�yL��i�TMAS�M%2�X(T�B�`�\7==�    �J@�    PQfff���k��T��ˡ��W~�LÐ��W���صW��c�������F5U&ƔN& �+�󚙼o�>]�_�j�вE�-�jl�"�ǣr��ީ[W.����:L��x�Z<�z��hb)�D�  �a``�>'��k���v    �rF�    P1nݺ�s��ie�6B����)�Q��_��7�s�~���4M�|�������};�>=>j7� �,���u�F�!\W���V5���-��./夥�k��c�F�����&�3�Mf��Y;ٽ��v�=�    �rU^g�     �gΜQ� T�i�)�-��S�á֎.;�n�Q�@���=Ӄ�q�L�W.�. ��g-t�{0m�����p{lS��7����EцFFi/����)X������_��i�T���匦��
,ʙ���ѣGu��uvv
    �rD�    P�_��Z� T��a�ڭa��.���إ�/�(_ (�������Fih l�|>g��ƍ�*S�kܤ��-�k�\�����N���Һ���ijk�W[j��Jdt)�t��;P��?gϞ����t    ��p    ��������!w �/�v�9�S��m?��jԱk��w���JW:���٧�P���E Pjr��7?�F���"�Xc�xohnU��^F��Z:��=���Y��o
���x<�0���RZKټ �������k��&��-     �w    @Y�u�Ν;g��(_�a(�u�9�Q��e��kP����ҵ�$[U!�sY�LM�-�V+���>� e'��|'����T�Ԣ��m�\.��,����kia^�x����e��LN��2v�@��v�{��w�{$     倀;    ��9sF���P�L�P�߭-5^��;�n�ɶ���Ꚛ�Ҳ�R�܃i; 8=>�٩I� *K:�����=�Ex����ukq��{�{��]��RP�v�&�T"W��g��(/��wG�Ձ���)     Jw    @��f�:r���7����q���n����.>6�vt�{��T�
�#�J���1;�>1<�TbY  Tkg���	{ܸx^�O��[��ҪM[�������w�L��1��TWا-!�&�3�Jd�+uʅ��v��Y����7���     (e�    e!����T*% ���0���WNӐ��U��Աk�<>���V����)M�kr����n�`  ���_�������ݭ�{��������g5�B5Z�/��X�um5^���Y��S�t�F__�r�7d����    �j!�    (y���:~����� ���۩�W�~���s�ϯ��{յw�\n���2锦�Gii �)X���`ָu墜.��m۪���[s{�����Re���p����l*��xZ�s6�������ӡC���0/    ��    ��v��5}���e&�q��Ƨ��e?�#�~�EmپC��6-�  ��\6k/���6Vg��7�mS�q�3���tt�t��1�0T�s�����tN�񴖲݁R����w�yG�������    @)!�    (YgΜQ� ���ץ�Z�B�G���u����K;�e��XoV�njlD��jr�ҩ�  ��Y���G�����|jڲ��7�l��ޟT��A�P��E��0+Zc1���bZ�{ �+����?��~�;utt    �RA�    Pr
��>�����@y���j��~l�۴��oj�J�}��	M���M�VS�r  �/�L�^�M{8N�55�a��m���?���1T�|���MM�pw����_��a�c�TY;:}��g�9��_~Y     ��    ���H$������ J�������֧��a���Ҫ]���b�M��Z�/؁���w4;5aU  @���s���ճgT��i�Vm�ڮh�\���Y��Ǭ�{Mԩx&��4Aw��ݾ}[�ӟ�$�4    �F"�    (����裏�-��.+���V��尟�tti��_�6V'�����f&����A{,�  ����Y{�]�,�F�۶�i�6�7�|.���V�{ryI�,�vhGԯD���xJ�I��@)�����Çu��!��n    �Q�    JB__�Ξ=�B�  ��0�z�G[j��9�[;�k�/)�k/��jr��h�V&�  (����\��.�[�Z۴yk�}o��_��J�w�����F��� ����%���;z�7�    �F �    �p�}��p_YY��c��������B���Z6������hjtD�<�\  Pɲ��F���jr�C�4Vн+�Skȣ�xZӉ���#����ѣz�W�u�V    ���    6���~��q���	@�q���n����v�v��y[�v����k,�N�j��؈
��  @���LK��T��1fGا�G�iM.tJ�����'�h~~^���     뉀;    `C$�I9r���@i��훃^;h�"ؾn2�&��j  U��4���W<�hl�Fw��@I�ꫯ4;;�?��    `�p    ����رc�d2P:L�P�߭�Z��K:�����P��ݒ  P�<V�{�X��
�ǿ	��F�v�{����׿�UN'    ��c�	    XW������O�BP2C��{�V��3M�Ԗ�;���_+�VWryIc�w4^�S|  �;��w��L2�1����;���7�T(     k��;    `�\�r� J���󹴵�/��ߍ�{^����aa�d�i����'G��  x�1jWا�G��f�Y�8���jr�ӟ����&    �V�    �ũS�488( �!�s��֧��a?oli�����±zau��9M��j�������   O��4��+�i|)��)���F)
:y����G۶m     k��;    `MY>�?���1�x����S��贐l�����o�_�������>>tW�,�+  ��*��:���i4��B:' ��:�s����q�۷O     �6�    �5��dt��-,,�ƪ�����Zϣ�A�MM����75�g�x{85����ӧt2)   ���S�cNͧs^Li9�N9�F���/�s>���     XM�    kbiiI���R�� l��rK�OQ��~mh��~���-�󙝚���~��P*�   �W��T�>���tO*�+������/�i�    `5p    �������(��
���j���ﶟ�D��������)�xóI./id�OC�ohia^   �x�SaOPS9��SJt�����>�������I    ���]    V��ȈN�<�B�@�<S[j}j��e��5����ߪ���`�3�e3�;�{��5;y_+++  @i��}c>��^�������䙗�eaaA���:$��/     �w    ���q�>��s�p��ZB^5�|*>���U��_�k�~��Cx:+��éI�뻥�;}ʱ#  @Y0����b�:�K�����i噣�"�J����z����F    ��"�    X�Νӭ[����Q�ǣ��>��N�:������\n��t�jlp��'�  @yr������\v��T"# k/�˩��G�����,     �w    �s�׿����AX_u~�l�92C[������ˤS����ۚ��/   T��TGا�A�F�i�&ٙXk�BA���?���/���[     <-�    �gf]�<r�fgg`��x��V��-�������[�?)��krdHC�ojjt�~  ��e-
�����ix1��l^ ֎�������E��׿     O��;    ���R)���{J$�>�.��j|vs�%ڰI{�;�7����ZZ��ȝ>ݺ���   P]j=N��M���R9:k�֭[������      �w    �S�.L>|X�tZ�a��r9L����\�߸P8�ݿ����;���;�s���&��4t뺦���&A   T��ϥ�ש�DV#�)�9F���ؘzzz����4M    �s�    ����z{{�ϳ�;�����A�Zk�r|��$�Ш���d�~��̴�nߴ۳�   ��d���n��\_J�~qs����]�p��!��n    �S�    ��ݻwu��i
l��%+ʾ)�Q[�_.���v�!�������h��u�=�   �s��c��n��}&��շ�����{O����+��/     ~w    ��u�Ξ=��m�T�ǩ�H@��{���r���K�>+�n��G��)�%�  ���u���ks �������\��L&���_o���jkk    �!�    �YW�\��˗`�x����j���V�-�]r�����l:�{}7�`{|~N   �j��[�L*�{Ie,�VS.�ӱc��ꫯ���^     �7�    ��t��y]�~] ֆ�0�R�UK�'���_�u�.��v   �=�x�^�s)�uj,���rFv4VM>��G}�����jmm     ���;    �G�>}Zw����������?'�(��I�*��ibxH׮jvrB   �z����x��wih!��tN V��ʊ}�������     �p    ���ǏkxxX V_��T{دZϓ���ڽK�U���yݾ��[7�I�   l�ӡ]��p����\^ ��r?{����v�b�2    �#�    �Q(t��1MMM	��r�������>��F�뺺U-VV
�֝�W5=>f   �R�8��>��DF#���U��p��%�R)���    ��;    �[V�������ܜ ��w�1���Z�\󩿾�m�|��*]*����ۺ{�k%��   J�Q<�o
�U�sid1��d�E��*�~��������V    ��F�    `�f�z�w���$ �'�q�=�W��x�ﱵ���i�{0m����  @�p��:�>m
�5��T<���300`7�<xP    ��E�    �d2�w�}׾�:|N���^�w?�����ڴe�*M����{���K�NM
   (W�bֽuA=Hf5��R&_�g7::�?�P����     Չ�;    T�x<�Ç�[@x~�!��������ںw�4MU�T2��[vc{ryY   @�����85Oib9# ����:z���|�͊�    �w    �b������Q.���W�q�3���X��ٶ}�*��̴�޼��������  @er���������|RKټ <���99rD���I�    �	�@    �Rccc���U(�u:��S푀��U���MM��DU�V����{v[��ب   �j�w��[ЃdVË)e+���<��[o��^�97    �tp   �*t��]�>}�p;��Ц�G�a��Ըڶu�R9�f����Tb).   �Z��\
{���� ����L&��_��W    *w    �2�n��ٳg��B{�<Bn�:#�<ksz��r��c��I|a�����V>�    �e�������bJ��́��N�u�����
��    T6�    PE���k]�pA ���4�V�SsȻ�����e����܃iݹ~U#},�   ~D�ǩꂚLd4O���3�Tr��zzz���+�
    P��   @��z��.^�( �.�s�+��a��{m۱[�l�x����W/ivrB    ~�aHM��V��BJ�iv>�F>�Woo�^{�5���	    P��   @�r�= <�ˡ�H@��4���E7�
y����//*>?'    O��0�3��\*��Ť�y�܁'U(��G����    �<�   ��}���ꫯ�陆��oq�����jo7�~��$�Ʉ�޼��׿V:�   ���:U�j|9��Kis��r?q����?���I    ��B�    *؅���_�ӳ��;����u}_�0���[�biqAw���[ו��   `u9�� �Q����bJK�� �<+�~��I<xP---    T�    P�Ο?��ׯ��q����}j
z7���ڶ��h��NM���eMie�I   `�\��5����bJÁ�e�WO�:�����jmm    �2p   �
�駟���O �N��VW4 ��ܰ�ö����`��//��v    ���ѩ��V����BR�ivQ~�r?}������jkk    ��p   �
��'����_ ���4������߇��Wc��_�_)�&���֕/�pzJ    6��ahgԯߴ��s~�r?s�8���    �w    � 'O������Ө�[��A;��ںw�4ׯ=�
�����K�8�P    JK�ϥZ�CC�)=L���+�~��Y�1!w    (o�   �B�8qB����'�q��*�u�Tl�޵.�S(�5zg�nl_Z�   ���.�]�#~�&����Y�Ν+�{���    �<p   �
p��q��i
z���al|k�cu�6+���{�Y�뻡����\^   �����=N��ӚJd��YM��ϟW.��Ν;    (?�   �����j||\ ~���PW$�p	��?�u�ڵ�g�)ݹ���\��~   �<9MC�^E�N.$������K�.�a�]��g�4    ��!�    e�p;�d������j}2K���1�˭����:=�L�m�C�����    *C���uA�.�5���!^ �e���B���|��^    �|p   �2T(t��QMOO�O�ꎅt;T�Z;��t�^�|:�P��_ڭ��\N    *��4��ƫ�ץ�I%s��������߿_    ��@�    ʌn�������q�!��������l���;Vg�t��   @�	��W��RF����]V��ڵk�9�_|Q    ��G�    ʈu!������� ���۩�h@Aw���#�6nz��A�   �n�a�-�Q����\R�<m���B�ׯ_�i�4�   @(���     ���v������ڭ���Z��(�v�.�����J�   �
�z�>�1��}9c�z����n�^x�    Jw    (���z��� �0�ӡ�j=.�����O�u�   �k��87r��|Ri�܁oY�>���k{>�o�>    Jw    (===�������=��,����6om����_O�   ���u;��.��xZS�� <b�ܯ^�*�ө]�v	    Pz�   @�����߿/ ��u:��̈́�hk��]H�������ו�l   �d����Z��V��BR� <r��e���;�~g5    ��*ϫ�    P%N�<���q��:�[ۣA;�Q����M[�~���Yݽ�n]�X|L�"   �g�:r5����TV 5����cB�    PZ�   @���?����!�.�i�+���l�]2��Y>����v�=�L
    ��5���4�tjp1E�;���/��r���C    ��@�    Jп��/
�w��=���r�*wm�w~�B��ᾛ�y�����   ���t;uw>��LN@����Ϟ=+�0���.    ��#�    %��O?�ݻw�ߜ��ma���^U���f�o��o�wt��9--.    ֒�ahW̯�DF�S���r7MS[�n    `cp   �b]H�����x]��S��m۱˾�����t��y-��    �S�߭�ǩ���♼�jf5�[�N�S---    l�    P"Ν;�[�n�� H��5xد͡�hm��r�y[���G�����   ��b-&�hl)��xZ@5��˝:uJ$�    ��;    ���/�ƍ����Ю��.�*M(�g~���q   @)0��5�Q��T�\R�|A@��B�O�֟��g566
    ���   ��t钮^�* �4<��0U"�   ���ˡ}u-�4��
�V�BAǏ�_��544    ���   ��ꫯ��p9Lm��    �N�PWا�ǩ���
+�����8�^__/    ��!�    �
�_�xѾXT�Z�S;�Br;L    6^��e7��'����FV�����_]�XL    ��A�    6��k���_�vFql��iK�O�a    P:|NS{c�/�5��a�>����o��p8,    ��#�    �l``@.\P�<�nm��pz    J���%�����'�)rG���r����[o��`0(    ���
2    ����}��'4��������i�    ���ǩꃺ3��\:'����y;vLo���<�     k��;    ����I�8q�p;���4�	�!��`    (7��nGԯ�匆S��M&�ё#G����Mn�[    ��A�    ���̌z{{U(T��ǩѠ|.�     �)����Jd��I*�ROO��z�-��L    k��;    ����e{�bkc�����W[�~    T��Ԟ�_��)M'��I<�C�    `�p   �5d5:���{�f�Ћ��r��*�u	    PY���Z�"��.$�+��sss:~��^}�U    Vw    X#�LF���r�Q�ǩu!yl�    �,�u���>�D��P=&''u��)<xP    ��C�    �@�P��Ç�H$T��W��C    �*�s��hh1��;١z����ܹs:p��     ���;    �������E��i����    �����������BJ����Ν;�x<��/)    ��#�    ����W>Pm�n�vՅ�u:    �^�>��.���J�
��͛7���={    x>�   `?~\�MSЫ��_�a     ���޺��Χ4��
�t+++�r��~����    xv�   `��={V������0��!�     �ɚ3n��4�p��bZ�����>���VKK�     φ�;    ��˗/�����thw}H~�C     ��F�[A�S}s	�������z��W���     ��#�    ��ƍ���/T���jn���     �9��}u�]H�a*'��
�8qBo�����     O��;    <����?^+l��*aRg$�MA�     x�⤲;���rF��8��J�����ӣ��zK�`P    �'G�    ���ȈΜ9C�U��rhg,����	    �g�p+P�c�%�)p^��q���ߖ��    ��pE    ���̌N�<io7T��ϥ��ݶ    ��q;�B}P�sI-dr*U:��|�����2MS    ��G�    �R"�бc��&�������'� �    X=�"�1�F�i�/�T*�|���~��!    ~w    x
�\N�V6�P����hPu~��    �k)���G~���)VVT���9�:uJ    �p   �'T(�p�ոT:�ˡ��!��    ���|���T�\R�|A@%Յ���/    ���   ���������J���[�    �^.����?��B&'�������F;w�    ��p   �'p��MLL�t�5>m���0�    ֟��zg̯�xZ�Ki�feeE�.]R Ж-[    �>�    �3�\����>��a�U�w    ��d-�����4uw!��ʊ�Jb�ܭB��^{Muuu    |w    �	w�ܱ�@%��]���     ����*�UM��%��T�B���Ǐ뭷޲��    �F�    ~���>���Q	�T1�[ݱ��<     �&�rh_]@�sI-dr*I.�ӱc����o��fW=    x��;    ����E����MJ@�j��ik�O�A�    P��E�;c~���_J�$�tZ===v��i�    p   ���d2z������T"�i�;T��f0    @y��fo	y�w�\H)ώ{� �x\'N��_��    �   �wX�����ݜT"�ˡ��5�9i    ��:�˞�ޞK*�g�=T���)}��z�W    Վ�;    ��#G�؍I@%�x]�Y���    e,�rh_]@�&��e>T���!�B!�߿_    P��   �7>��#����DMA�:#�     ({.���X@�I=HfT�k׮)���S    P��   @����5::*�uDjy    @%1�3��ij4�P	VVVt��9;�i�&   @5"�   ��Y�Hׯ_Pi����!E�.    P�Z�����̧TXYP	N�<���zK�PH    Pm�   �jccc�pႀJ�s:��!d�    P�b^�<1S�&�-rG�+
����?��9�D;    TfA    �V<׉'�m�JR�qiW]P.�)     �E���޺���Z����L&�cǎ�o��    ��p   P�r���9b��dSЫΈ_�a    �j�q���B�	ͥ9�򷸸�S�N����   �jA�   @U����L&T��Z_q�    @53iGԯ�xZ�Ki�nllLW�^����    Հ�;   ��s��	���
��Pw4�:�[     ��-!��NSC)VV������׮]SMM����    ���;   ��b5ݻwO@�p[[�ׇr3�    �5�\��η����|Y!��g�*+�
    *W�   T���!]�tI@��B�V��
�    �r;��.���J��ʕr�裏����]^�W    P��   �
sss:u�}��~��cA��     ���:L���7��b��;�W.�SOO��~�m�&�    *w    /����ѣ��x����=�A�    �'�4��uw!��dV@�Z^^�ɓ'�ꫯ
    *w    �P(�ȑ#J��*���_�5>    ��g���>���F�/B�����_|��^zI    Pi�   �h������;�|w,�z�G     ���=r���ZP�n߾�h4���N   @%!�   �b]�xQcccʝ������z��    �Z�.{�}g>��
1w����ϫ��V���   �J��q    ��ݻ�ꫯ�;��Ԟ��]    ���:�+�׭��rB�(?+++:~���~�m��~   @% �   �������������\�m���a
     ����8����Ä����r���u��1����ir	   @�#�   ���R)����P�b$�[��Ү���!     ���S�c��%��������_]    P��   �V������d2�Yc���Ѡ��     ��ihgį����R9����:{��~���	    �w    ���WKKK�Yk�O��~    ��g�#���BJS	JP~U__��۷    �w    ���˚��ٻ�/����㯻�]f�aeSDC�|�6mOlN�tM��&��6�Q������ *"3,�,�ܹ��&]�����<�|��0?���~���ʕ@7{tC_��   ���C����\�=�&�V+'N��ƍ�iӦ   t#�;  ��>����W�
t��:��M�X�	   ���UR.$ߞN������^�O~�T*�   t�;  �����s����C�F�R1On�@�+:   t�ͽ��|���������Di4���~���~:   ���9  е��f����m���Q�\ʁ-��W�   �i�ZΓ#}936�FS�N�h��=z4O=�T   ���  �Z�=�\&''ݨ^.��[S-��  �����v�>:��;]�ټys��   t�;  Е�z�\�r%Ѝ�+��<0�9   ��7�}mS;r���\3�-N�<�M�6�?   �@�  t��>�,��կ�h�֓'7�T,   �.��ڑ�ٱ�L���A��ʡC���3Ϥ\��   �ϛ  �U�����/��@��W��@��   нz�z�bco޿1���;�avv6?��O���O  ��	� ���l6�a�F��l�汑�h�  �����<9җnLelz6���!ǎ�w��   t2�;  �5�{�LLL�̓�����+n  �5����؆z>��|9%r�;�?>�6m��?  �N%p  ��[o��+W��͎�zv�   X{ڑ���zz��|>q7�N�<9��  �N$p  :�g�}�_��W�n�gC_�   X���\L>���Z�V:�g�y&�l  �<�T  ��6>>�_|q���E�P�c����   `}x���R�����}ˢ����������/��/  �4w  �c5�����?M��t�R�������^	   ��<�ۓr!���T$�t�۷o�رc��w�  �N"p  :�s�=����@�(�yrS�j=   ֧M�����|pc*MK�t����g���ٷo_   :��  �Ho��V�\��=�b��e0}=�    �ۆj9�o����ij��p���/�#��7  �� ��s�ҥ��W�
t��b!_�< n   ��P��'6����̩��`�V+�3�<�rYF  �>o&  @G���ɋ/�8�ݠ����^q;   �TJyrcoΌM�!r������СC����   �6�;  �Q����m�0�A��q{]�   ����o���c�����������5���o  `5	� ��q���ܸq#�j�RlH�,n   ~��_G���t��n|��lݺ5   �E�  t�O>�$�Νt��,����    ܋����FzszԒ;��^�O~�T*�   ��;  �ꦦ�r���Z��|���?�:�JI�   ܟ�w�'G���g暁N�h4r�����?�s   V��  Xu?��O�M�����r`��   X�z��'6����d���P7n�ȉ'��o;   +M�  ���_~9�n�
t�v��uq;   �ڑ��#�9=*r�s�;w.=�P�o�  ��$p  V�G}��?�8���+��<�q;   �D��v�ޗ3c�n���LG�ɏ���j�   ��;  �*����ꫯ��j:Y��[�S,   `)UK�<��7g�&3%r���������я~  ��"p  V\����~�����d���r�`J�v   `�T~��>:�I�;�֭[y�������  X	w  `Ž�����Ɇj=��恔
�v   `y�o�{b�/g�&31k����f۶mٹsg   ���  XQ|�A>��@'����M�v   `��G�{sF�N�:v�X�lْ���   ,'�;  �bnܸ��G�:�`��'-�   �������щL5��N�l6�����_��_  ���  ��h~<��s�?�ST�9�yP�   ��v���H_N���@w�ܙ1yꩧ  �\�  ��8x�`&''����oL�(n   VW�ȝv�<��Cٽ{w   ���  Xv�O�ΥK�����4����   @�hG�O����wrw��$���Z6oޜ���   ,5�;  �������o:UoO)_�:4h   �I*�K���K�w�,��9������?��O  ���  ��ir<����?��˥|}ˠ�   �X�R!Ol읏�g�������9v�X���  `)	� �es���LLL:Q��?��J�   �NV+�䦾�w}"�"w:����cǎ<��#  X*w  `Y�6.^��D�C�v�^�   ]�V*�ɑ��%w�;����m۶T*�   ,�;  �䦧�s�ȑ�Z��<���[���   @ש��ٿ�7g�&E�t���������~  �� p  �ܿ�����h:�|ܾup~�   �����#�3c�i���cccy���o|#   �%p  ��ɓ's�ƍ@��)���z�   �n��#�9�;��w�͎;222  ���  K����9u�T�������-�v   `��oG�zs���D�W��ʳ�>�b��  ��	� �%�l6���|�:I;n�������  ��e�R���#ro�.G���ɑ#G�W�W  X(�;  �$���LOO:I�Xȓ��W��   �M����G'"q�|��g��㏳gϞ   ,�~  `����\�|9�I��B��4���W_   `m���w���nM�a�����g۶m���  ��r�  ,ʝ;w��k�:;��l��   `=�T��\���ܲ��k6�9t�P~��  �~	� �E���~����@'yl�?�{�   XO��V2;��gw�Vۭ[��_�"��  ��!p  ��ѣ�}�v����З���   ���}�:�����L`��;w.;w�̖-[  p��  ��|���y������z��   ��=2XK��ʵ���jj�Zy饗��3Ϥ\��   ���  p�fgg��/:ɶ�Zv�   �d�p=s�dtZ���jO>|�p����.   �B�  ܷ������)��V�w��   ��;\�܍Vn�mV�_|��g�f���  �C�  �}9u���at���<6ҟB�    �K�P�c�9;6���ji�Zy뭷�cǎ���  ���  ��Ν;y��7�b�Z���k   ��J�B�Л�F'2�hVK��̡C����O  ���  ��g?���!t���R��y0���   ��)ybc;r���9��X=����#*��ַ  �� �{Ҿ>���ہNP�)������Y    ��J�8���̌ȝUt�̙�ݻ7���  �m�  �t�ƍ���ہN�>�������    ܻZ���7�sfl2�f+�Z:�g�y&   ���  ��~��ٴ���k/������   `A�zJٷ���c�Ѹ�Z�����������  �	� ����ѣ�����b��'6���    n�R�ޡz>�5�VK�������{��lݺ5   ���  ���]��s��:�c�2\�	    �7R��L��������_γ�>�bэ�  ��  �U�����-8�vo�͖�j    X:��*�;�̕���j�����E����n   ~C�  �V�����&V�C�l�   ���s���f+קf��O>ɥK��}��   �	� ���}�p��j��[����    �|��2;�ʭ�F`5���y��gS.�X   �;  �4�ͼ��K��6T-��
   `�<����c������F��W^y%����   p  ���fff&����R��<���   `E���<ގ�G'sw�Xi��y>����ٳ'  ��&p  �Ӆr�ҥ�j���9�e`�P   ��S-�#r�L��
��'Ndǎ�T*  �/�;  0ovv6G�	��R���mH�\
    +�����6����T�-�;+��h��_�?��?  X��  ���~>r��R($OlHū*   �j���g��oNV���hΝ;�}��  X�T  ��a�իW�����P�	    �oS�'�s�|6~7��Z�VN�<�;v���7  ��#p �unzz:���Z`5�����    �9��W3;���ə�Jj6�y�����0  ��#p �u��K����v���`=    t�]C��4�����u��ͼ��9p�@  ��E�  ��ٳg3::X-j=ytc    �\���щL��VҩS��gϞ���  X?�  �N����7���ޞR�o�O!    t�b!y|co޽>���f`�4��>|8?��  �w  X�<�Fõ¬��b!OnH�X    ��R,���9=:��V+�Rnܸ�s��e߾}  ��;  �C}�Q�^�X�B�����{J   �{���g��nLVJ���ɓ'�k׮T*�   k��  ֙���ǎ����2T�:
   ЍFj=�1��g�w+��]��������   k��   ֙�fvv6�vֳ��    ����j��\�򝑕s�ڵ\�pa~�  X��  ��\�t)�/_����Jv�   ��g���F3wf�+���_ώ;R.�]  `-�?  ���µ�jVZ���#�   `m(�}�yot"w�|sde4�9r$�7  `�� �:��K/��ݻ��V)��恔ڧ�    ���>�7���щ�5E�-���J�o�  `m� �:p�ڵ|��'���n��q{�T    kO�\�c������cǎ��g�M��#  �Ew  X��f:�V˂+ﱑ�T�z   �e��r���Ӂ�0333���_�e  ��Ge   k\�#���$V�#C�l�   �����J��|19X	/^̾}��u��   k��  ְ���|�ᇁ�����G�z   ���k����\n��V�+���g�y&�b1  ��!p �5�^H�����J)���   ���PH�m��{��j�.��{�nN�<�o��  ��;  �Qo��F���+�Z*�k�Sj�f   ����Pϻ��i���>Ⱦ}�2<<  `m� ���O�>XI�B!OlH��:`   ���^.���z>�9�VK���j�����K��  `m� ����ϧ�t0+kT�f   �l���P_%���,����������/  @�S  �s�ԩܼy3�����j    �7��W2٘��t#��ڷ��۷/}}}  ���  ֐������[��4X-g�po    ��3T�Tc�Ǎ�,�V���_~9?��  t7�;  �!/��b���+�R*f����    ��V*��p=��&�h���ƍ��㏳gϞ   �K�  k��˗���VJ;j����TK�    ��R/��?�9=��˥��u�ĉ�ڵ+Ţ�  Э�  �F���+�XQ{7�e��   �?lC����*�t�n`95�?~<O=�T  ��D  �5��^���d`�<8P˶�    �W��+�l�el�XN/^�O<����   �G�  ]nbb"gϞ���j9{6�    �מ�Z��_=��ri�v�ꫯ�駟  �}�  ��<�f�a+�R*�̓)
   ��U*��p=��&�h��e||<gΜ�_r  ���  ��G}�����JhG�_�<�j�    X�z��݃�|xkz~i��/���ݻ7�J%  @�� @�j��;v�+fT�F   �xk�<����;3�����~�ȑ����m  ��L  �.��+�dvv6��e�@-    �T��U21;��w���ʕ+�϶m�  t�;  t�7n����0T��ލ�   ��T(�w���F'3=�,��G���g�  ��  Ѕ^xᅴZ��r���yb�@
�    ��+ylC=�G'3�'�dzz:o��f���o  �|w  �2��Nn߾Xn��}#��;    ,��r1;����t`��={6���O___  ��&p �.2;;;�2+ᑡz6�+   �嶹ޓ�ٹ\��,�������J����  �lw  �"����\`�m�U��Po    `���eb����(�ctt4/^�Ν;  t.�;  t�+W����ˁ�V)����    �J*�G��ywt"s�V`9����y��S,  t&�;  t��^z)��
_=�7�G�    ��j�Bv���ͩ�r���������SO  �Lw  ��E��):,�]�2\�	    ���Z9��=�bj6�.\��dxx8  @�� @�k��gΜ	,������    V�ΡZ�4����,�#G��G?�Q  ��#p ���K/��l�S�\��    ������p=�Nd��
,�۷o��?Ξ={  t�;  t��W��ʕ+��T($�7��X    t�j��=C��c2��Z�VN�<�]�v�X,  �w  �`/��r`���П���C    :�p��m}�\��	,����������v  �Ρ`  �u���ܹs'��6�V��@-    Щ����\�g�K�>ȁ���  �3� �5����XN�r1�F    ���ճw��wG'�h�K��j��ѣ�����   �A�  �W^���l`���Sj�    �Z*���ZΎM�ڵk�r���<��  V��  :���xΟ?XN{7����   ��1T)硾J.O��R{��رc��O~  `��  �ü����a�l�f[-    �m�Ts{f.�s��499�w�}7  ���  �A.\������ri_���H    ��z�P�;�'�h
ai������\��  �j�9  t����\
�B�4�r�    �V�b!�����t`)5�?~<���w  ��;  t�7�x#��dX>��3\�	    t��ZOn�����l`)}�駹u�V���  ��;  t�����9s&�\�j=yd�7    �V�����\���Ri�Z9r�H~��  Xw  � /��b���ˡ\,f���    �ZR,${��9=6�f�X*�����g���  V��  Vٵk�����ˣ�R-    kM_O1��+�t�n`��W�O�8��;w�X�m  V��  V��Ç�?��r��_˖�j    `���ۓ[w�5�L����l�z��ɟ�I  ��%p �U��{�e||<��=����    X�
�B�������6���tΝ;����V��  �J� �*i6�y��7ˡPH�����    ָ�b!{�jy��T`����9r$�w  `�� `�=zt��SX���2P��   ��1\-�ޞ\��ݕ�s���\�~=�6m
  �2�  �
�����G���z%��   ����Zn��e��,��Ǐ�G?�Q  ��!p �U���/�_m
K��T̾��    �zT��yt���F'3�j���۷s����ܹ3  ��� �
�y�f._�X�R*    ֫z���*�p�n`)�Z��<yR�  +D�  +쥗^
,�����+   ��nko%�f�26�,�������{��׾  `y	� `]�t)ccc����Sʮ��     �a�`-�3�m�K�ԩSy�'R,�E  ���  V�ѣGK��ճo�?�B!    �(�5X�7�Kann.���/�g�g  ���  V�ٳgs�Ν�R{x�7�՞     ���Z9��z�O7Kᣏ>�7���j�   �C�  +��lί��R믔��`=    �o�s���ىܝk������^�_��_  Xw  X'N����L`)�<>�?�    ����Bv�r��T`)\�t)7o����p  ��'p �e��Ϟ=Xj��{�W�Z    �P����=�br6��?����  ��  �ّ#G277XJ��r��    ܛ���uw.�s��b�����իy��  ,-�;  ,�;w��O>	,�R���7    �w�B!{�j9=6X
�����  ���  ���Ç�j�Ki�p_��b    ��3P)塾J.O�kbb"~�a}��   KG�  ��ڵk��/KiC�'�j    f{57g��m��7�̞={R,% ��"p �er�ȑ�R*�ٷi     ��
�ޡz��H��,���lN�:�o~�  ���  ���r�֭�Rڻ�/Ւ     X�z�8�������b�>}:H�,� ���?k  XǏO�e��������}�     Kc[oOn�m���\`1��f^��<��S  O�  K������T`����ytc_    ��S(�g��S�'ҴW�"]�x1������   �#p �%�^ii����R*    XZ�R1��r��t`1ڷ����k����  `q�  ���|������ʖ�jF�     �ckoOF�gs{f.�W�\���x  ,��  �H{��̙3���S*fφ�     �k�P=�\�H��
,T{���������   'p �%���[ogI��ЗJ�    `y�J�l����Ÿv�Zn޼����   #p �%�h4r�ܹ�R�W���    `el�dt���ٹ�b�Wܿ���  X�;  ,�cǎenΡK�T,�ё�     +��ճg��wG'�jlttt�	  p��  �H333���Keφ�TK�     +��\̃��\��	,F{���?�a  ��'p �E:r�H��f`)�z���    `ul�f�n#S�}Y��7o�/��֭[  ��;  ,���T>����R(
ylc    ��S���3T�{����x�����O  �?w  X�W_}�z;Kf�po�=�     �����m}�\��	,���x.]���۷  �ww  X�;w�����0P-g�`=    @g��_ɍ�F�猜�p'N�� �}� ����+��Y�B!�F    t�R��]C՜�
,���d>����ٳ'  ��� �ܾ};��y
�B`�����    ��U���ۓk������/)p �� p �x��K��RΎ�z    ���p57��ef΍�,���tΝ;�}��  ���  p��_��/��"�X� �؟��     �c������܍��B����w  �Gw  �O���j`)<4P�`�k    t��rFj=��,���LΞ=����  ���  p�����Ū���9�    �;����L#�f+��N��_q/�  ~7�;  ܇#G���rx��=:ҟR�    �;���_���w1;;�w�}7�G  �w� �=���Os����bm�W2��    t����\�j���\`!Μ9�Xq ��C�  ����_,V{�}�H    ��S(�k��wG'�h4�� � p �{����֭[���9ܛj�2    t���b�������B�>}ڊ;  �w  ����Z`��zJyh�    ��=�_͍�Ff����������  ���  �\�v-7n�,֣#�)    t�R���k���T`!�  �	� �8v�XZ-+<,ζ�Z��=    ֆM�r���rkf.p�fggs����߿?  ��$p ������,FO��]C�    ֖]C��s�N�6RX�w�yG�  ���  ~��G�Zog�vo�OO�    `m��
y���Kw�����LΝ;�}��  �/w  �n޼�/��2�C��<�_    �6=�_���l����j��� �� ���ꫯ�������     kW�;�#ռc*p��������G  ��  �[����/�,Ǝ�����    �m��rFj�N7��ԩSw  �o�  �[���[�V`�j�b�    Xv�rkf"��o�ܟ����?>�w�   p ��cbb"��y`1�n�O�X    �>���_���Ӂ����o� ���  �9r�z;�2R��?    ���@oO������\�~��w>���ر#  ��	� �i_z����B����    `}�9P�����:y��  "p ����W_��΢l��^.    X�*�l��s}����+W�d۶m ��L�  �6===�',T�T�Ã�     ���Ռ�m�iO��t�ĉ�˿�K  `=� ��;v,�f3�P�7��T,    X��c�U�ٝ����իW��  �+�;  |eff&/^,�`���}�     �=�_͗S���3�����/~���� ��J�  _9~���v�P(d���     �F��Ǉk���T�~ܾ};_~�e6o�  X��  �{�����z������+    ��X-g�����F�^�Z������ ��H� ��w�ĉ����T,d�Po     ~�G��5�H��g7n����x  �� �u�ܹs��j��R1     �M�\��z%W'g����������  Xo�  �k��^ff*�0�=�<4P    �ﳽ���ӳi4͸s�^�:�Q�T  �� �u���,Ԟ})    �{�����������j����������  �z"p `ݺp�B&''1R�dc�j    po��˹6U��l3p��g�g�b�  X/�  �['O�,D�PȞ�}    �W�B!;k9=jx�{�l6��;����F  `�� �.]�~=7o�,���z��R     ��@O)#�rF��{u��Y�;  �� �u���ぅ�)��`=     ��@57�6�l�I��ȇ~�G}4  �� Xw&''s�ڵ�B��؟R�    �����y���Kw���;�#p `�� ��=z4��i�_��-��     ,ƃ}�|19�Y3�ܣ�x��˗��C  �:�;  ����l>���B��M�`�    X��%�;�9k:p��z�-�;  �� �u�7������Sg~��_��g8
IX>���wk�)W���S�����ڿ|�U�hW�lY�@� 3�l�ȑ% �������K��t�G�;��n�i]��.    ��p�V���vl�{f�ɼx�"���brr2  `�	� ȍ,l���	8�l�=[o    8K��VㇵV�I]�~=����=  `�	� ȍ�7o���^�i]��c���	    8[�B������ĳg�bgg'��j  ��Rh  ��}�]�i�Iį&    p>��w��������;�����o�  0��  �������	��ǣ���     8�R!.U
�|g?�$?~�n7�Գk  ��� �\�������*��d�     ���F+���6�9�l���o��/��2  `	� z������pZ��ע�&    p�*�4>���ik/�$��k����ي;  CI� ���ӟ�pZ�b!��T    �"|4R�������q�x���q�������  ��� �����+++����z���v    �bd�I~8R�ٍ����s�� ��$p `����G�z�n8��J)��+    p��k�Xj����g{{;���bzz:  `�� Z�n7fggN���     �h٩��Vbf};�8��ύ7��c  �0� 0�n޼�N'�4.��1^-    ��p�Z���B4�<��x+++�����SI w  �֝;wN#������    �ٯF+q{�pׯ_����:  `X� JO�<�V��N��h-�%�I    ��5Z.�d�k���y��qt��H�4  `(7  J��N#M">�    @?�d���N�z����t:q�������  ��� ���-������G��(��     ��^�V���cŝ�ݾ}[� ��� 0t���?Y��T
i�Yo    ��ߍVbmg?<��8;;;������  �N� �P�v���ѣ����z;    Ї��4.�J����6��ύ7��c  ��� 0Tn޼�N'ऊi�V    �}<R��;��ur)�XYY���ݨT*  �L� �P�s�N�i|2V���v    �OU
i\�c�eŝ�]�~=����  �A&p `h,,,D��
8�,l�h�     �죑J,o[q�x�?�n�ij� ��%p `h���g�i|:^�B�    @?+�IL�K��x�N�w�ލ�?�<  `P	� 
�r���J�Ie��^�    � ��Q�g���Xq��o�� 0��  �?��O��P�S�t���v    `@�$>h��ɖw�ngg'���bzz:  `	� x�n7=zpR�z�t�z;    0X>l�c���]�/-�q�F��  Dw  �_����t:'��Ɇ�v    `��$�5�1���6+++������  �� ��w��퀓��
q�z;    0���˱�lǞw�q������  �� ������V+���D#     U�D|8R�ٍ���y��q  � � 0в��^�J'3Z.��z9     �t�t�������������>  $w  ���~,--�ԯ&�    0�V��x���6�o�� 0p�  �o��6�]�4�L��~�f�    Wk�Xh�Yq�^�x�f3�F  ��� 0��ݻpR�Zo    �H�D\k��w�q�ƍ��o  �� ��������'�(b�z;    0dVܷ�����277  0H�  ��ׯG��='�	G�    �'�V�G*1��p�N���ߏ�>�,  `� 8�v;���N�^*�T�     �h�V����س��[ܾ}[� ��� 0p����;��n�I��x-�$	    �a����(���n�Q^�x�f3'� ���  �{���D�X���J     �j�x�lǾw��ƍ��7�  �;�;  eqq1���N�Ӊz�n    �]!M�z)��G���  w  ���ף׳@���4���    ������9B�Ӊ����g�}  ���  �v�KKK'�w��H��    @>�w��Iӊ;G�}��� ��'p ``ܸq#��n�q*�4��     ȓ�x�jG׈;Gx��E4��h4  �J� �����	8�O�k��   ��)�IL�J�p�lP�o�	  �Ww  ���b�Z���d/p��T     �>����~t{f�9���\  @?� 0�_�p��׭�    ����\��b��8L�Ӊ����g�}  Џ�  ��v�KKK��^�|h�    ȹk�R,��aÝ�ܾ}[� @�� ��nܸ�n7�8�ף�Zo    �RH�J��Z{���؈f��F#  ��� �{333�)�I|d�    ��G�J,����s�^�w00��7�  ��;  }�ٳg���p�Gk��    �W���T�+�V�9ܓ'O  ��� ���������$I�[o    xՇ����#������\|��'  �D� @��v����p��F%*�4     �?�b��b�h�����w  ��� ��u����t:��d�     ��Ñr�X�s�������45" @�� з��8ΥZ)�B     ��r!�B4���^�w�܉/��"  �_� �K�v;�����w���    ��Z�3�������  ��;  }��o�=X��-c�R
     �6U)�\!�ݎ��l\�F#  �� �K���8�'�     ��$�F%f7v��%��_�5  �� �;ϟ?�V��6�b!��+    ��֊1��D������w  ��� �����瓱j     p2�$��z)�������ӧO�ڵk  �� ����ɓ��)�IL7�     �q�Q��V;�F�9ĭ[��  ��;  }eff�`%�棱Z�$     8�l<�r��Z�������v���i  ��$p ��d� �6�1��Xo    x���X�ޏ^ό;?���w�ލ�?�<  �}� �7��v������H%J�1     �VLc�\������	� �w  ��_���1���Z     ��>l��jss3Z�V���  ��E� @߸w�^��\iT�V*     �n�\���][�N����׿�W_}  �� �kkk����6��    �Ƶz9^���c�;  �� �������h�c�0     g�R��B��n��vwwcii)���  �u  }a~~>�m>�     g#I"��J1���[�n	� xo�  �w>�v�p�R!�+�;    �Y����Is7����y��Yt��H�4  �	� x����p�i     ��b�ĥj)V��^��t�>��  ��&p ���?�8JvL���     ��Z�,p�Pw��� �^� x�~��ǃ8ʕz%*G�    ��F1��r!6۞��s���CEi�=  K� �{������G��     ��L�Jw������~���  \$�;  �M�����p��r1�*n[     ��T�s[���t^u��=�;  N) �{s�Ν��8�G��     �|%I��Z���j}}=����X� pq|� ����R*�q�!p    ���R<i�F�.����|��  E� �{��}����Ñj�I     p�i���X��x�����  \(�;  ��_�������p��k�6j�    �"]k��ass3��v���  �� p མ��	8��z%*�4     �8�b��Bl�;/e�E�oߎ��
  �w  .\����ŋ��|4f�    �}�����ѣGw  .�� �w��̓�8�H��R     p�j���j�n��R�ٌ����V�  p��  \���Z     �~$���K1���R6\t�֭���/  Λ� ��j�bcc#�0�4���r     ��\��b~k7�ʫfgg�  \�;  ��͛G�n���$    ��SJ��,cuw?ढ़����܌���  ��$p �B=|�0�(�Fk    �����yU�׋۷o�W_}  p��  \�lգ�jf�Z�F�     ���BTi�t�/���	� 8ww  .̍7�=�0�F�    @��R+��V;ढ़��X__����  ��"p ��<~�8�0�4���r     �?���1�l��^u�֭��o  ΋� ����������Q�B�     ���&1Y.���~�K  �I� ���y�f�Q��V    ��3�(�������a����  �� p �B<y�$�0�R�K�     ����Q-����dz�^ܾ};����  �� p ��mmmE��
8̵��     ��J�s[퀗�>}  p^�  �����/�)�iL��    @��Z/�|��^�����������  ��&p ������F%
I     ��R��d����/ݹs'��_�%  �	� 8WقG��8̵�j     ���e�;?3??/p �\� 8W�n݊�3K9�D��R!     ���BTi�t��V�u0tT�� �l	� 8W>8̵�    ɕZ1���l��~�?��  gI� ����ߏ����ו�$.�+    ��Z/�|�n�G�	� 8sw  �͝;w��uT)o�nT#M    ����L���������<<*%H  ��. 87���8���v    �At�^��3?��c����}  �Y� p.�������׍��     �g�R<Xr���2<� p�T%  ��l�=���u�T    �����\+��f; ���~�N(M�  �� p �\d�Q��W�     `p]��^�w������&  �,� 8Ϟ=x�T�|pt-     ��^L�־�\�333w  Ό� �37;;�N'�u�#�     `�e+�����  ��"p ��ݹs'�u�4�K�R     0�.�J�xk7z���᣹����O  ~)�;  gnqq1�uӍj�I     �R��D�k����w�
� 8w  ����R����n�Q	     �ǕZI��O�={  p�  ��[�n��^*�h��    �0����&���t:��!����  �_Ba ��ZXXx�#�     `��IS�b,m;ٕ���?� ���  ��f�;;;�J�$�6*    ��R+	��ɳg�  ~)�;  g��x�D��B     ��r!��4Z�݀l��jE�^  xWw  ���Ǐ^��H5     ^�k�x����w�^��?�c  ��� p&��n������&q�^     ����We�Hw  ~	�;  g������^u�^�4I    ��UN���c}w?�ŋ�Hi�  ��;  g";n^7=R	     �_��.p'�"���ŧ�~  �.�  ������WU�i�WJ    ��"M"�{�o�߿/p ��	� �����boo/�UW���    �$1Y)��+�D,//  �+�;  ���۷���W]i�    ��r�$p�@�ݎ���  8-�;  ����|���B���n     ��x��4���Q"~�����/  NKq �/��v8�UW��    �N�$1Y)���^��'O�  ��;  ��ݻw�׳���	�    ��r�$p������PR��  �!p ����	x�h��b!     ȟ�r!Ji{]�8y�$=z�(~��_  ��� �_dyy9�UW���    ��R�K-+�Dܿ_� ��	� xg+++�����;    @�MUKw<�<  ��  ����.�U�RT
i     �_c������N7ȷ���X[[����  ��� ��^u�z;     s�R��-�;w�ލ���*  ��  ��v��f3�$I�J�     p�V���� �I  ��� �w����G��xi�R�r!     h�
Q-$���.!�Z�V���G�(S �d|s ��<x� �UW�     �����x�l��&�������  ��� �NVWW^J����;     ��r�(p����� �� pjϟ?�N��ҥj9Ji     �R�X�z��=��nmm-  ��  �������    8�TE�N���^lmm���H  �q�  ����B�Ki��T�     �Z9��333�?�!  �8w  N������F�K�b�$     �u�B�b��n�oO�<� p"w  Ne~~� r����+     G���e�=�^�x  pw  N�޽{�ʎ�    ��\���=�:�N<�<���  �F� ��,--�4^-E��     �Q*D���n�	�y�)	� 8�� ��v��l6^�R�     �R�O�V��nqq1  �8w  N,[���z/M��     Ǚ�܉���:TJS�� p4�;  '������F+Ũ=�    �x��4Ji{]C:y�)-,,��  p�;  '�����e��     �P�$q�Z��������  ��� ����9����J     �IMV
��
rnyy9  �m�  ��ݻw���L��F�T     8��r1
I�r��j���~��%  �"  '2;;�ҕF5     �4�$b�R��;�A�=|�0~���  F� ������4U+     ��T�$p�`XI� �Q�  kcc#���2�Bc�;     �7Q)F�Dt{A�=�<  �(w  �����G��I3��r�     �.��}�\��]+�y�+���D�Z  x�� �c����t�^	     xW��{�e�J333��_  �N� ��^�x�)�i�WJ     �j�Z�d#�ٱ��,	� 8�� ��Z\\�N�����"I     �Y)Mb�\����y���  p�;  o�	/M�+     ��d�(pϹl`��lF��  x�� ����!��g��    �/5Q)��f�c�^/�߿���  �*u
  o���������     �T�X�j!��N7ȯ���;  o� p��������L��     ge�R����=ϲwQ  �:�;  G�w�^�Kw     ��d�K�� ������nG��  �G� ���<y��Ҩ�
     ge�\�B�D�����Ç���.  �%�;  GZ[[�L�+     g)M�-b}w?ȯ��9�;  ?#p �P�V��XH�\��     ��d�(p�9�K  �N� ���ݻ�I�����    ��7^.�����n7�4  �� 8���|@f�Z�B�     ��j1�Z���� �z�^<~�8~��_  d�  �����K�r     �y�(������� ��;  o��ۋ����̥Z)     ༌��x����J  �Kw  �p����L�T88     ��d��ͽ����|��ގn�i�  � xCv$d�j�     ��$��������bqq1>���   �;  oX^^�L�J     �m���	r�ѣGw  � ������H($I�W�     ���#��_nF�P��   /	� ����كc ![oO��    p�j�R$흿������V  @F� ��<|�0 s�V     �(#�$��^$�Wr);e����155  �� ��YZZ
�LV�     \��F�Zތ��� �<x p @� ��5�̀Z��b     pQ��5��pA��c��  �� �������0Q+     \�4Ib�T���ݨT*A�lnn  � �Iv�#d&+w     .��1��E\�z5ȟ�����ىj�  �� ��<{�, I���
�    �xY�~s�iLMME�P�gvv6~���  �%p �'/^�)�TH     .�d��b!677cbb"ȟ���; @�	� 8�����`�    ��%;etz|$��������Z  �ow  <z�( #p    �}�6>�W�c{{;j�Z�/��;  �&p ����\@�$1^�    ��d��{u�݃����   ��  X^^���&     ��h�#�r4���t:Q(�|���� �� �[[[U��     �L�������܌��� _�={  �� ��P`R�    @�9�766�9���  �� �x��a�z� �
I��;     �_�����ۋ����jA~���F�ۍ4M ��� �����R$     �_�T��F-֚�+���y��i|��G @�� ���Հ���v     �����A��l6���D�P�cnnN� �Sw  ��jL
�    �#�&F㇅���z���A~���  �$p ȹgϞE���RH�^r{     @��:6i�D�׋���{�lmm  ��` ȹ��ـ	��     ��b!���z,o4coo/����V��������(�� @�� rnqq1`�"p    ��d+�Y���V����5����  �E� �skkk�    �GW�?���lF�ӉB�����  ��  9��vcww7ȷb�D��     ��+��H�$z������A>���  �#p ȱ�X��a0�6^)�     �~S.b�^�������i�Z @�� rl~~>`�Z
     �WW�?�{{{����j5~�i��j���h  �w �{��Y�X�m     ���X#~|����Y�,pϏ�D�/��"  �% @�e�ɷB��H�m     ������~��ڊ˗/G�$��3� �?J ��ʎt̎�$�F+�H�      ���ʥ�Vbsg����G�ٌ���`����  �"p ȩ'O�D���m�Z
     �wW�?��Z�{>���  �"p ȩ,p���[     ��ձF<x���ϭV+:�N
�`�e��Y�^�V �|P�  ����r�o�߮��w     �ߕ�7�ڳ����`�e'����o~�   �  9�����h��4	     �wc�J�ʥ�n�����=?�  9"p ȩ��N�m��v     ��qe������s�ݎ��ݨT*�p[[[  �C� �C����9�o�R     ���2���=���܇_��  �C� �Csssc�;     �cz|�ϲ�}jj*�$	����^t��H�4  ~w �Z\\�^*D)��    ��1Q�F�X��~�ϲ��jE������R\�v-  ~w �Z__�m�j�    �����_m�����>�V���o~~^� �w �j6�A����
     0x.���ܳ��N'
�B0�VWW �|P�  ������C^�m�b�    ���-�fkk+��ǃᵱ�  ��  gfgg����UL���     �A35R?����M������  �A� �3O�>�m�\�$I     M�X��Z%6�;g�s�ݎr��l�i}}=&&& ��&p ș�ϟ�6Z)     �K#�7�L��>55���y�; @� rfkk+ȷ���      ���z<Z^{�����}�-//  �O� �#�n��xN�m��6     ��55R?�������ىj��/^  �O� �#O�<�^��W��F��     �K#�H�$�����V��ë�j  �O� �#Y�N��VJ     �,��'�x��f��/_�S�ӱ� �w �YYY	�m��     ��wy�~h������Q�Ղᴰ����� ��n ȑ��� ��*n     |S������d+��ᵼ�,p r� �Ɏl$�FJn     |S#�#��/_�$I�ᳶ�  7u @N�������k�\�B�a>     �o�V�r������v��j���h�'�  7�; @N<}�4ȷъ��     �l����桿�"h��p���  ���  '�|-��    ��x[��l6���E�8�t�d�����r9  N
 ��X]]�m�R
     S��#���Y�>22������O ��$p ����moIz���|�dI����K���Z ȓY�=c�߻�lk3�̮mI�DuU� �)e��BT������A��� �:      ?\�}������� �M� P��b��b2��    ���hg�qܯ7_����H۶QUU��_�5  ȗ� � ���v��u>��    ���?�}3p���qA^�u~  �r (�O?���|�?     ��>��~���w!��=?��2  ȗ� � w�Fu     @n���{�E4Mu�<'���ݫ��   ?w �|��1(W5�\�    @���揾���>޽{�c��?<�ۿ�[  ��; @>����ۻ�     rs6�d4��v������	�3���?� 2%p (�r��uf�    ��]�g��͗o�{���mۨ�*ȇ� �%p �\w`�^��r�O|�     _Wg������������˗   OJ ��Y��|�k?     �z6{�=���V�   OJ �����wP��Q     ���'��"��}� ����&㪪 ��� 2g��l���Q�`    �|]ΦQ����|O�w����Y��O�>ŏ?�  �E� ��ϟ?庘�     rVU���O����w�w/p��_��W�; @��  ��k)���     ����ٓ�n�}0y�� ȏ�  s��:(��H�    @���G�Ӷm�V���/i���	  �#p ������	庘�     r���i�z��D����  ȏ�  c��_�r�*&u     ����E������?y�n� @~�  ���cP��q     P�Q]��tw��w��4����t:���d���b8�@ �ķ; ��}��9(����}     �q=�=�w�w�{�������  �x �ؗ/_�r	�    (���,��G���>|� p ȏ�  c��"(�|X     ��j>{����ml6���A�nn��  �"p �Xw8K��#�;     �x7�<��݊��=n4 ȏ�  S���~��4�QW�     �R\L'QU�h�ǟ�t����u�>7 �G� ���~�I�^�ٰ
     (I��O�q�\?���z��.�C�L��h ��� 2���?�:��    @y.��'�n����2H[�4ѶmT�� �\�^  2�믿��     �Ҽ�M��?o����b!p�D�\�Ç @�  �����5�    (��|���.�����1��}��Q� ��; @����5��    @y�=#p���.r���A�~��   � �L���L�j��    �Ҽ�Mٻx�)����p�1 @^�  j�6��	�t6�5    �2�*�&��[m��~7���� �� @�>~���e�3�     �z7�>9p��v��lb<�r�1 @^�  ��矃r�-�    P���4�߯�O~��-pO[��
  �C� ��_~�%(�|T     ��r6y�������*HWw����]���  �� d����A��F��    P�w��޿\.�mۨ*2)�n8� �A� ������Lê�q�     �r]�=/p�t+���}��)��?�#  H��  C��*(�|$n    �l����x����?#pO���M  ��; @��ۧؒ�����     p9�>;p'm>C �|�_  2ӭ�����L�Q     P���$~�����o�&��uL&� M�� @�  ����SP���     �b6}��t��tm6�   w �����A�f�*     �t�����>����4u+�  �A� ������\ӡw     ��=�}�^?D�u�=U�
�|>  �&p ����]P�I]E5     ��l2��`���Y?��A�����  �� dF�^��Ȣ     t�A��x��ͳ~n�\
��������  �M� ���j�i6�    �o.��g�݂;麽�  �'p ��f�Z�1V     ���lq�i���Y�x<��c �<� 2���2M-�    ��:��/�K�{�,� �A� ���j��>(�l$p    ��\L'�\I_^^�q�1 @�  ��_�r�,�    ��:��w�ݠ�`0Ҳ�n ��	� 2"p/װ���r�     ������.n_��1�N��4M  �O� ��ϟ?e���      ��hX��o�����s��.pO�b���|  �K� ������L�Z�     ��|6���ų��������t7� �&p �Hw�J�f�:     �?��N����z���m��̤�������� �t	� 2�]�I��#�;     �����������Z�,�'�˗/ @��  �l6A�,�    �?��M��nXH������   mw ��4M�if�     ������}�Xć����  }w �Lt�d�m��b\     ��������n��ƅ���LJ��u  �6�; @&>~��i:�b0�    �?��GQWU4�uk����A:��m  �6�; @&>��iRW     |��d���V���q�1 @��  �����4
�    �[f����b�e���f���x  �I� ������L��     ����C��n��6F�Q�������� �4	� 2�Z��2Yp    �o����ӗ˥�=1���w ��	� 2��R��Ђ;     |���nd�ݻwA:�E  �.�; @&6�MP�qm�     �e>9~������  �� db��e��    �������n��e6��� �6߼ 2��R�z0�a5     ���&��j����� �� @��  �h�6(�dX     �m�aú�]s����r)pO�z�  �%p �@w�����L�U      �7��vyx�l<-n> H��  777A�Ƶ�     s6�o6�h�&��ͪ)� �M� ����۠L�;     <j6�;��u�����?F   ]w ����e�    ������r)pO�~���m��<G H��  �rM�f    �1g��ѿc�Z鸿�����   =w �,��L�a     �����/����e��`�����  Qw �X)פ��     �����{�w�df�Y�_�|	  �$p Ȁ��L�`ue%     s69~��#pO���]  �&�; @v�]P���z;     <Ũ�^ۦ9��,�˸���o�X  i� d`����w     x��x��q��[u�� H��  m���    ��M�]&�>�w���X��1�L�~�>'  �$p H\���4�     <�t�2��r��'��  �� $���&(Ӹ�     x���e2��j��v�  �$p H���]P&�     �t/��^���s2 @��  �[,A���*     ����F/�{v���k8�����  ]�i $�5���     O�R�n�]��o��>  H�o�  ���k\�     <�K��󙳳���,� ��78 ��	��e�     ���鿻�����
  �"p H��2ՃA�w     x��^p�����  Aw ��	��4���     ���0�jm�?�w����l61����  i� $�;<�<�     �y&�a,7��]����ߺw  �#p H�v�2���eTYp    �皎^.p���/..���� �&�; @⚦	�3V     <O���t�u+�  �G� ���n�gT	�    �&/�o6�h�6*g���}F  �G� ������k��     �\/������t���  Mw ��5M�gT     x���W����Ƕ�m  ��; @�,��iT�    �^:p_��A�v�   =w ���V�\�     �y&���N	� �$p H�b��T,�    �s��/; ��M�Dm����  i� $���>(Ө�    �s�^!D�V���΂�i�6  H��  a��2(�`0�Z�     �6�|*�^��=��� ��� �X,����     p�q]����w�ɂ; @��  	��^�Z�     뇛R_r�[��o��&��q  ��; @�V�UP�a���2     P�Q]�f׼��k���U�u�?�`��  -w ��u��gX�p    �C�������l6������  �!p H�n��c�     7z����z-p�)�Q  �� $L�^�ڀ;     �[pi]�N?m��   -w ���m�gd�     6~�w+��� H��  a��44�     �^'p���18���  �� $�i��<u�p     5z��N�O&��_F �G� ���m��*     �Ì�����k�{Yp H��  a'�Tp    ����;�#p H��  a��4��     {�w��` @z�  	��iX�p    �C�ւ�����  �� $L�^&�     p��+-�����n�1���h�&  H��  a�A)��     ��R���V���"p H��  a�2��    �p�+ޔ��l�~� �G� �0�{y�AT�;     jT�^��-��/w ���  !��    �8��Ҷm  ��; @���8���     �y��}��=,��u��  =w �D��L��     �RW��6$��n�=���  i� $j�Z���     p�nPf�J��f���t�w ��� ��R�     p���b�J�g8�"p H��  QG�T�p    ���A�_�wo��   'p H���LU      Ǫ��;q��_��}  ��; @������     G{��}��E۶QUfk���,  H��  Q��(�w     8ְ~���*�L&  <��  Q�&�$p    ��_y]}���{b��
 @r�  ����Ay*g�     p���;��� @z�  �j�&(Ome     �&p ��� @B*�;     �~�+S��m   �� $ʂ{�*};     m���]���c`��ڶ��?s  ^��  Qݡ(��     ǫO�(�E��$x{w ��� %p/Sm�     �Vׯ;o6�{Ot�;  �� $�i��<�    �x��4�;�`8
  -w �D9�+��     �w�=��v��( ��� %p/���;     �7�Zp��; @Z�  �j�6(��     �w�A��� @Z�  ���^*�;     ��{��E��(x[�� �E� �(Ke:Ţ     �:�y���<W H��  Q�&�$o    ��2p��5M  �C� �(�;     @�	����; @Z�  �rW�S-�     @�':o��v��3 ��; @��     ��N�[pi �t� e�     ����� @Z�  ���^��DW�    @�N4��Vw��u]o�s5 ��� � �T>w     8����2݊���mYp H��  Q�2Yp    ��:p�N���� �E�       @QN9'��  ��	� UUU      �|Չ�y[u]  �� $�Wg���     �6��p @Z�  ��     �����y� ��; @�,M��,     �7�6Mm�z���  �!p       �Wԭ�O&�   'p H���2���      �Ӟ��]����C� @J|{ H���Lw     H�n�ގ�j  i� @BZ�;     �����&  ��� $��D�ڶ     �8��1Ղ�۪�:  H��  Q�2�-�    ��N}�.p[w ��� 5��w     8���� H��  Q��Դm      �i���m�>�<�y��  �"p H���2�-�    @����x��?,  H��  Q��tq��e      Go1(#p;áD
  %�� $���,Mӄ�     ��{2]��۰� ��; @�,���;�~�E     ��[-�  �� $��Dy��     p��8m���n4�s5 ��� � �<]��
�    �h��a<  =w �Duk���7     ��V�  �%p HT]�AY,�    @��  �4w �DUU��;�v�&     �-eڶ}xy�  �'p H�p�\i���     ���jP�������   -�( �D�F���A{��w     H�����  �� $j2��x���f׶     gۼ�y{�sZw ��� %p/�o�w     8^�
�KQUU  ��; @�\_Y��ܛf     �q��� ��; @�,���w�     p�]�6�2�ӳ� ��; @�������~oѻw     x9��Q�u  ��; @��M���}��    �X����v���x� ��;  $��;     ���}�r�'p H��  a�� ���9����	��     p����w�{]��i��  =w ��u�������     �X����� H��  a݂;e�-pߺ�     ��ց;�3ʣ  R� @ºw������b?     m��K!p H�op  	s�b~�ݴ�      ��{�A��n���i  �� $̂{��[p    �c�堌�Ӳ� ���  fq��?�~�+S     o9(#p?��h  �E� �0�{����,�    �Q���]�~Zw ��� &p/����     p��ݿ����I��( ��� �0�{������     R�Xp/�x<  �"p H���������òL]     x>�{YF�Q  ��; @�\�X�<�����+�=     bۼm���t�6��1�S� �G �0W*��������Wy     8�f�{��g���Nc:�  i�M  a��$��?�]w��    �C���{g��	�Od6�  i�M  a'��]Qڽ~��     �����i  �� $́\��v�����;     ��C2��QUU  ��; @�\������C��֡7     �C2_;���u�;  �� $���,�����V]     �`������Ӱ� �&�; @���σ�}u�}'p    �C�a��1fsu]  �� $l:�y�z����     ��m�����OC� �&�; @ºk��C�|}�][p    ���aHƳ���F @z�  �A����?�߶�-    ��m,�C� �&�; @��F𜭯po-�    ��6۷_p�l�4�  i� $n8�v�����}-p    ��m[��� @z�  ��w�e�     ^�~���9���4&�I  �5 @�\����povw     8Ķ�GX.p?�; @��  �����M�~�`     ��mv�苦i������f�   =w �č�� _�Zp�O��|�    ���4�YN��_�t:  ң� H��=o���;     <W�ܿ���3�� ��(b  7�L�|}�p{�k�<     ����l���uvv  �G� ���l��{��mf      �M�כ�	^�t:  �#p H��=_�������l     x��?���_�`0��� ��� 'p����[V�    ���tC���uu�;  i� $n>�y����҂;     <�J�^��  �� $�ݻwA����7�me�     �m%p/�p(� H�or  ���fW,~/�&M�;�^	�    ��V�b� �� @�+��	����m      ϳ���|�x��L& @��  �(���n����     ����c��g5]�����i  �&�; @F�Q��� /�_p�    �s���^E�m۟�>G��<  H��  ��8���ٛ���n㡯�     �}��[pUggg @��0  ��fA~;����     �4��� ҥ� ��t:�����r��w��     �dݳ��m���\\\  i� d`>��y�`�o�     �g��ryy  �I� �yz�`{��     �4�r��� @��  ��鱃��F�     Oշ����\9\UU @��  p�b�]p���      ��o7�Zp=w ��	� 2��ݻ ?��[�;     <U����g4  �� d�[��^�����{��f     ���x3j�l������ @��  �����}��    �S�q8Ɗ��L& @��  ��(v��-�p���`a��     ��vMۿ�\��:��i  �.�; @&�C_�r�ءvw���b2��    ��,��[o︝�u���   ]J �L�f������Ֆ��F�     ���魨�_���y  �.% @&&�I�����ϭ�     ��,6�\p���; @��  �p�b~�r���+U    �O�=�۶^���e  �.�; @&,Q�婋-��^�
     }�<�,ggg @��  �x��]P�;�     �����?u���QUU  �.�; @&�����,zz�*     ���r�r( ���F �����?,RX���S?�Ū��3     �ݙ�b����s��7� ��	� 2�]�ؽ��	���+U    �/V�]�B�b�f�   mw ��tW.
����w�ӑ��     �5�M?��;�_�|>  Ҧ� ��d2��z��9�݊��     �n��o���;??  Ҧ� �H�Hq{{��;���     ����+�/���2  H��  #)���w     ���%y��}  �6�; @F...��,�     �M���_���u  �6�; @Fؕ��     |���PL)�ATU  �M� �W.��9�-�    ������[pY��(  H��  #WWW�C�r�^     �Ϻg&��.(�x<  �'p �Hw�b�j�&H۳���h�6jWn    �tg�mk���$  H��  3�Ջ��t1�b����C[     ��/�~߂�Vޗuvv  �O� ��n�b�Ze���     �G��MP����   }w ����󸹹	���Ŗ/�u�u      �c��,��� @��  �q�b��~@     o��yY��� ��	� 2��ݻ }-�     p��D�YpY�׮� ȁ�  3�)�0��~4     ������y9UU=�  H��  3>|�sg�     �`���v�D�=w��o��:  ȃ�  3�������,ˮmc���l<
      ��O�/g<  y� d����ߋ$|�!��A��     ��n�	�1�� �<� 24�Lb�Xe�[��O��     Hc���sqq  �A� ��n�B�����-�     �oR87?�y _wuu  �A� ��n��ӧOAY,�     ���n>�?��c  ��; @�����/�KP���*     ���[[p/ɇ �<� 2��?i;�@ۂ;     �ݮmc��e��*�C @.|� �п�˿�Yow��51�     %�[�1
c��e���   w ������~����n����<     �dw�MP��t  �C� ��n�b�Nc���#p    ��<��݂��8??  �!p ��l6��v�
     (���yyI��� �|� 2uvv�?�t�b���5     ��}������Ç   w �LuK��_�����2     �t����?  �� d�A^�n����_     (�r����	��=��� @>�  ��ӟ����@}׶q����t     P���:Ra��x��(  ȋ�  S�����ݚ7e�Y,�     �f�
�1{& ��; @Ɔ�al�� =�,�t�~     P��e:���㝟� ��ٻ���3��/ �)J")q�,K�▇�޻�\��]՗�T�S��$�'�<E�e��'� �igQ'qEX�y��w�<�������� ������sh�2     9��W������d  �_�  }l||<vww�lJ���v�����j     @^m[pϕ�g�  �E� �ǒŊ�ϟ�����w     ��lF� ;��
܏off&  �/w �>f�"ۊ�b�Z�#���f��clh0      O�*��I��x��'  ��� ������u�Ֆ��}�;     ��]�V�n��xJ���H  �	� ���=ێs���ۏS     y��d���x��� ��#p �c�bE�\�l6��9�Q{�R     ț�j-����񌏏  �G� ��FGG�\.�s��=cO�    �Iض��+gΜ	  ��� ��MNN
�3�8G�-�     �L�Պ��zd������� ��#p �sgϞ��O��s�gI�덨5�1<P
     ȃ�j-��vd�q������  ��� ����l�M�]nٮTc���     �<��ۏ,��~<� 066  ��; @�[XX�鸇�M�;     9��ųD�~<CCC @� �����(�J�l6�l9��     �"kw�d��w7>>  �'�; @���D�R	�币�Fe/      /6-�����T  П�  9p��)�{w�e�\�V�Er     �\����Fd���x��� ��$p ȁ3g����r�-�=l7[���ۏ���     �~�����q�n�nnn.  �Ow ��������:Ȗ�Xn٨T�     ������]��nbb"  �Ow �XXX��$ۛ彈ٳ     �l��Yc���  �K� �ɂEK��� ;N$p��b     �fe/�Ƃ��  ���  '���c?{�%yv�-����    �(�V��D�XpwSSS @�� �D��.pϖ�8l���;��ؐ�:    �O�k�Y|�V��� ��%p ȉd�buu5Ȏ�:lo��b���     �~��W�,������  �	� rbff&��� ;
��:�j,�    �S�l�R)8����s��  �K� �.\����+{     �j��Yd���  �M� ���Ӈ��V�dC�@�����c�:ɂ;     ��䆾���;���݌��  �M� �#CCC������J���f�X���~-�V��    �/���7�,������  ��	� rdllL��1'�'�5��j�L�     ����^d���ݜ;w.  �ow �9s�Llll�qR����/p    ��l�ewاT*G777  �7�; @��?>�߿d�I�ɂ;     ���޿���Gg� ��	� r�ҥK����qR��z�     �o�L����y3<<� @� rdbb���f�d�I.�7[�(9�    �'���_oD���ͩS� ��'p ș���(��A6�ԁ��j�F�3��     �`m7���&�D�ٳg ��'p ș��)�{�����nY�    @�X/�EVYp7��� @�� ����L<~�8ȆB�pb���nv�     ���|��]�Ʌ ��'p ș������d�I��v��T+     ��V���jd����J�R  �O� �3�����v;H��<p��עVo��?     �m[��h�Z�U��  �A� �3��tdd$��쮚��I��v+�p�t     @����E�%k����T  �w �����g��     ^�^�D�Yp?����  � p ȡ���XYY	��\�2�h     �5��  ��  �����޽{A�ub�     ���l�N�Y&p?�B��N�
  �A� �CKKKAv$G�f�y"�V�ވ��ZL�     d�zy/��vd���hFFF ��� ������O�^��$���NE�    @f���E�	܏���� @~� rj||<�����+�'��m����ٳ     Y�.pϝ���   ?�  9u��Y�{F���{u�     �U�l����[XX  �C� �S.\��w҇����l��t���     �i{�ß,���w �|�  �.]���y�~�ћ�vlU����X     @���f{�=a��h���N��  �M� �S���V��['����    ��Y/��&�N �|� ����X��� �:q�^�.�{s3     Y�����5�Gs���   _�  9v���{t��͕m��    ȖV��sgnn.  ��; @�%�G��։Cw�v���852     �k�{�l�#��o�P(���R  �/w ��v�Z��w�ҭS����S#��     ��uR�����K�  ���  �&&&���f3H�d�$�i�Ov�fe{7��
�    Ȇd�������d  �?w ������ ݒcw��8�_s�O�n     ���zy/��������  �#p ȹ���{t"p��ۏZ���     ����~4��EZ��ۻx�b  �?w ��[\\�����֩c���n,��
     H�~y��X,���
���P  �#p ȹ+W�į�� �:u�N��    �v�;��������h  �Ow ��:�988ҫs���x    @[�����ӧ �|� �������W���h4[1P�*     �S�E���``@����� �|� ������\�ޭv;Vw�175     �F�;������]�t)  �'�� ��/ƽ{����䓥+�w     �ke��B��v��EN�:  �O�  ���b
�h��A:u�ོ�?�7     ��U�{�  ��S3  Q,ctt4����tJ�u�?BX۩D�Պ�_~     H��A=v�k�/�o��ٳ @~�� ����)�{�%�q6��u�VlV�1=a    �tY��WH�ogaa!  �/�� 8t�x��i�^�ѻ�{be�,p     uVv*�O�1~���b  �_w  ]�z5���?��ɣ��v9n/�     H��>
ܓ!�B�������  �%p ��ٳg�X,F��
ҩ�ϖ&�{��vX     5j�fl��G��䝿�LLL  ��3  s�ԩ���	ҩ���F������x     @<��9g���3==  �O�  �M��.pO�N��m�
�    H��[��'��s�ҥ   �|r �o�~ҩ���[����     i�|[��7�B!fff �|�� ���r�J����{�N�>|/o�F�ՊR�     �K��A��k�O�lxx8���  �=�� �������a��_�~�t��v�ݑ_���_we�sS     ��lk7������;w.  �'g  ~fjj*����t*�J�h4:��?���    �sϷ��o�lii)  �'g  ~faaA��b�񻣁���_��B     @/=߶��GW�\	  �� ��y����C�N�>~o��Q�7bx�     ��ʋ[u?�����!��  8�S!  ?399��p�]�T���n�Wq.M�	     ��[������M  ��O�  ����ӱ���O7��6w�     ��3�{.���  $|z �%sss���J�އ_     ��v;Vw+�o�7�z�j  @B� �K�]�_|�E�>��w����b|x(     ��Vw*�h�����,��cll,   !p �%�ϟ�b��V����[O�>�܉�     ��y��2*p�ӧO  ��� �W������� }�Ƚ�ht��H�@�    �m�;��G�7�p�B  �_	� x�d�]��N�ܟm�     tS�ٌ��^��B�еZ���ի  ��3  ������ }����������FlV�qf|4     ��o���jG���Y�T����  ���	 �WZ\\<\i��u�:�'+�w     �ey��(������  ��� �W*���r�?��Y֭����v�^<     �O�v�	���  O� �k����S�[���N%��f�J     ��S���_~����ͮ\�  ���  �֥K����ҥ[��f�϶v�⹩     �Nz�ٟ��	���%/
���  �=�;  �u�������v;H�B��R)��f��'�w     :N��O���  �H� �k���HT�� ]�7���oG�     �F�����W�כ��	  �Gw  �hzz:=z�K��j���>Ճzl���쩱     �Nx���>}M6��'/��j�/_  �Gw  �hiiI��B�\{y��#p    �c�;t����zI����  ���  �����㷿�m��t9%��ŗny��\�     �	϶�y422�b1  �	� x��8<<���Azt3p_ݭD�ь�R     �IڬT�R�G�������  ^E� �/J�>ң��{�ޟ��_�=     p��l��z{B��zW�^  x�;  �������)�JQ(��nx��#p    ��=������5Y�|Ǳ��  �*>E ��nܸ���o�S�v�՗�����^ɂ{��?98    �I8h4c}w/���W;u�T  ��� �E�b1��ǣ\.�����Vo���^�L�     ��d�����:�k��/���  x�;  o%94~��wAzt{�%Yq�    pR����Yo��ׯ  ��� ��r��5�{�t�0�xc;>�<     p\�v;�m�F?
^��ڟ;w.  �u�  ���/F�X�V��C����^��bl�A    ��Y/��~��L��j���  o"p �%ǭ�� �P(��t˓͝�qa:     �8�n��z{B��jKKK  o"p �-,,�S$�ۓȽ^�w��|��%p    �؞llG���K�Yq���  �7� ��n޼_~�e��q�����͝�7�1X*     ��J� 6*��g����5���  ��'i  ������1��h�����f��6w���T     ��x�����CCC��Ξ=  �K�  ə3gbuu5H�^<o�����    �w�h}+�����.^�  �K�  Irx��G/���[�l��T,     �~���{���/+
q���  �_"p �Hnݺ����t�E�~�h��v9��L     ���h�����/���  �̧F  �d||�� Y�Ղ�K�N�cp����������    �#{��yЋ������	  xw  �lzz:�<y�Cr$�zྺ����a`     o��L^ݍ~����/�r�J  ��� pd�/_��Hr$�V�]�=��X�݋���     ���dc'��v��������ii)  �m� 8�7n���v����W+0�6�     ��Gۑ��_6>>�b1  �m� 8�dydtt4������ա�ǵ��立     ���nǳ����/���  x[w  ����\ܿ?�^����جT���h     ��<�܉z�y p�{�  ��  ��[�n	�S"yҳT*E�_$+�w     ~���ȋ^ӤU����L  ��� �Nb`` �F�{�L�Z������Vܽ4     �:�v;o�D
����ٳ  G!p ��%ɕ�����5�^j��kqjd8     �UVv*Q��c0G���+W�  �� �w�$���˃y��~{�|     ��<Zߎ����ڵk  G!p ��ݾ};~���>-Jo�4p_�    �z�7�"/���x��N�:�$  ��'H  ����`���G�\z+�wQ(z���T�zP�ѡ�     ���QދJ�y!p�����  ��� p,��7������j����IT�pm3n��     ��V7#Oz��j�$�<�n�
  8*�;  �r���{J$+��?��    xُ�ۑɝ�X,/�J����
  8*�;  �2==}x�����hZ�rfe���A�[�    �������8/���\�  ��;  ǖ(�={�V���3�w�     $�mF�?�z�j  ��� pl׮]��@����;     ���v���y2d��o
�B\�r%  �]� 8�[�n������X<00�F�'��zy/v��19:     ����r��{s���?����b�  �.�  [r���������u�^��W6���      ��l�=��$�ᅅ��  �w�5  'biiI��Iྷ�׳����M�;    @ε��x�����z��ݼy3  �]	� 8�oߎ/��2��v�;I��K�{��Y�ƙ��      ��n��A�y"p�I�]���D  ��� p"���bpp0���u���ae#�\��(    @^=\��z{"������	  8�;  'fvv6?~�N�T:�i6{�����F|$p    ȥF��7�#o,���ƍ  �!p �ļ��{�HVb��j�~���A��Vbzb<     ȗ'��h�"O
���+���g��` ��� pb�^���o��V��i��{�'~X��    ���խțdx&	��8}�t��  ��� pb�����Tlll���{������ʂ�>    @���x��y���|Z\�x1  ��  ��d�]��[��ý�K��A=V��q~j"     ȇG����+�###���~  �q	� 8Q|�A�����v�������~��_"|��!p    ȑV7#��0<��N��f ��� p�crr2�����I���j��׶�]��B!     �o�z#�wʑ7�BA���[\\  8	w  N��˗�����I��ܓ/3�n�����    @KFOZ�������s�N  �I� p�>���{���9����w    �x��y��{|�������X  �I� p����xT*��7�rP���F3�J    @��ۏ��^�Qv���  pR�  t�ŋ㫯�
z�X,���@4���u4[�x�����     �)���a��ܹ  pR�  t�ݻw�=��{�'��|]�    Ч��v���yT*�bpp0�nhh(N�>  pR�  t����᳜���Ao$�J��뿌Xۭ��^5N��     ���v9��G��_�p�B  �I� �1q����7�tX���_Y     �˃��ȫa�����?  �$	� �>�@��Cɂ{Z$_p|ty>
�B     ��f<^ߎ�J^�ͻ������  8Iw  :&9h&��z=�O��Z�'����A��Rb�vp�L���D     ��oE�Պ���133  p��  t���\���Ao�%pO�_^�    ����W��O�T���u�V  �I� �Q�o���P�S.�#�n����C�    �u��Z��V"���G��XXX  8i�  :��ŋ100�F#�4؛�V<\ۊ�    �l{��������H����{?  �!p ��fff�ٳgA�%O�
�h�ۑ���     }����ȳa�q���  �N� �q7o���Prd��ߏ4X�.��~-&F�    �*����"��a����b1�\�  �	w  :.Y���o~�V+辡�����q��\     �MV6"ϒ�{����ӧ#w  ��;  �8ϝ;���A��mE�����.^���     ��V<Zߎ<���v�Z  @�� �7n�{$m��J� V��q~j"     Ȗ׷��lF�����͛  �"p �+n߾���o��nݕ,�F�^�������     ��lDލ��F�MMM~�   �"p �+�C�����NU��pm+>�7bx�I     �b�Z;|�3ϒA�R�y���  ��& �knݺ%p���r9=_:4[�x���/�     ِ�Ιwɽ=�
�B���{  �$p �kn޼��y4�͠��xp��ٚ�     #Z�v|��y7::yv����W{ ���  tMr𜙙��ϟݕ<�:00�F#�b{�+;嘝<     �ۏk[Q�����+#9_pOƌ  ���  t��۷�=2<<���=����    ����ȻdLfpp0�*2�r�J  @�	� ��ׯ�o~�ԅ�y���T*�H���������G    ��ک�be�y7::y6==}� @��H  ����Ǔ'O��J�Ӧ�jŃ��xa6     H�/�d�����  ��;  ]�O��O�H�MM�UZ�V�ɷ���     )�j����� ��R).^�  �w  �nii�0����Aw%�2{{{�&�{�çmgO�
     ����V��Ȼd@fhh(�jff&  �[�  ����\���Aw�.pO|�lU�    �B^^^����۷  �E� @O|���H�4z���֗bx�Q     �b�Z;|��|�R)  �E= @O\�p��)σ���{���P(D�ݎ4i���`e#�_�     ���k�����Wɫ�  �Mw  zfqq1<xtW����G�|�lU�    ��v;�_��p8&�/�vï~��  �n� �3~�a|����[�w�3�iܷ�����=}*     譇k[Q�7��^Gͣ������	  �&�;  =3==}[W�ՠ{Ҽ2����    z���������W���  �&p ������K3i\����֗bx�U     ze�Z;|q����<J�K�s�N  @��F  詏>�H��e�A:�����#m��v�_^�ۋ�    �����Z�BrS�k�>44�Ν  �6�;  =555ccc���tOr�Oc�����J��0{��     �Uo6���F�BrO/��G�+�  �w  z����q�޽�{Ҽ6S��㍝X:w:     �+q�h/���F^}��  � p ��>����ꫯ��n�1<<|�8�j�"��z�,p    �o��?�k���}OLL  �� ���ӧO���V�=I�^�V#��o��V�S����     ��m��N���Ť�E�N�v�Z  @�� H���?~���ݓ���5pO|�t%�ύK    @w|�t5�I^���B|��  �"p  �ܹ�����V+莴��<Xވ�./��?�     t�n�v���O��OMM����<  ���(  ��<�y���x��Y����Q*���lF5Z����z�Y<     tַ�ע�n?�k��� @/	� H��?�8��_�%�dŽR�DZ}�d%n/�>�
    @gԛ�x���$���I���\�  �Kw  Rcaa!����V�ݑ���R;��;�t�t     �I�~�H�k��266y4??  �kw  R�ҥK���ݑ��U�z�,p    �o��?���y'ܽ{7  ���  ��'�|�}�]����F�^�GZ=�ڍ�J5����e    @'=�܉���U�Q����3g�  ��� �T����S�N���n���:́{��+�n\
     N�7��_���/��|�r  @���8  �w���������;��=��A������B�#    �II�۟m��>�ccc�Gw��  Hu  �������h�ZA�%�{�5���^^�;��    ����h���ύ��F�LMM���P  @� H�b�333���t^��;9ZD�}�d%n/�F�P     ���lƃՍ�ey�oݺ  �w  R飏>����#9֧=p�����v,��
     ����F���熇��a�$���v�Z  @Z� H��/���`�����FFFb{{;��ޓ�;    �1������Z𲱱�ț����.�  ��  �V�߿?輿.ҴZ�H���Xۭ���x     �n~\ߎ�j-xY��B�w��  H�;  ���'�ܻ$9`'+�{{{�v_>Z�����     ��|�t5xY2����dhh(fff  �D� @jMMMũS��\.�7::��������e����     �h��ˇ/e򲼭�'.]�  �6w  R�ƍ��?�1�$pςv��/���q1     8�{OV�W�c�~���  ��� �j�a������f:�T*>Ezppi��嵸{y>F��    �m�Tk�lk7x���122  �6j  R-	�gggcyy9�d�=�{�Վo����Ks    �����A��HB�d&On߾  �Fw  R��O?��>�,�$p��ގ,���J�Y<�b     �fՃz����Z��ۓ��ƍ  i$p  ������j�t���p��h�Z�v�z#�/�����     �;~�-����}qq1   ��  dµk��/�:/��	*�Jd����Ǎ��(
    ��՛����z�jɚy2 �'}�Q  @Z	� ȄO?�4�ݻ��e��R�^�?�Gk[qi�L     �j~�~��jy[o�������  ��� �	���133���Ag%�{�|�xY�    ��V;�y�����x���۷  �L� @f$+�}�Y�Y�b��)�Z�Y��[��[�qa��    �?�am3*�z�zY~9�R�׮]  H3�;  �1??###���tVr��J������    ��~j��M�{x2��������  ��  d�����/�:+9�ommEV<�؎����	     ^x����j�zccc�'}�Q  @�	� ȔO?�4�ݻ�V+蜡���gJ��fdŗ����s�r     �½'+���)p���8� ��� �)���133���Ag%+��r9�������|�    @�m��by;;7�^8|ɋ;w�  d�� ��IV�?�쳠���7[���x9>��     y��cC1�d||<�"y��ڵk  Y p  s���cdd$�����I�
�h�ۑ�>[�;Kblh0     �j{o?o�o666y����b1   �  dҍ7�O�S�9ɡ;�ܫ�jdE�Վ�/�'W     ���G�35^���K�i^|���  Y!p  �>�����/��j����d)pO|�l5~�t!��q    ȟ��~<Z��l||�0rσ����  �
�  �444333���tN�k�V�{�]�    ���ӣe��o!	������  Y"p  �>�����ς�)�J1<<�Z-���+q{a֊;    �+����qm+x�d�=y�4�;����  �D� @f������H��������������%+�    @~|�x%Z��Q�zi�X�<XXX���+  �C� @�ݸq#���?����5_?]�ۋ�c�T
    �~W�����������G^|���  Y#p  �����9���h[�阁������ȒZ��<]�_-]    �~�������R^�����  ��;  �688�����ɓ�s����//ǭ��(y~   ���ޝ>�Yh�>��-�؀1�;lll�l�Kg��d:==�n*5U���n:@��8x��]�*˖dk�۷�3�tX$Y����qT��*��`]��9/(�����>/��ͩ���?�y�  @%� P�������]X>E�>44�JS�����'}(     eu���L�Xo�����T��e�'�x"  P��  T����tvv����ayK�������J�)Vܷ?�&u�V�   ����ʩ�7���.�@� @%� P
�v��|�Oq�_�"(��-.w��    �l������������]ʮ��f��  *�� �Rعsg>���LLL��Q��{����e]�w    �TƧ���/@[[[���u����  �Tw  Jc˖-9r�HXŲM]]]���SiF�'r�ʍl[o�    (����f��l�j܋���{.  P��  ����?�cǎe�S�˦XqN%��lYכښ�     T�"l?y�z������X5oooOwww  ��	� (��p�xv���?,�J�G���Vܷ��    @�;r�j&����W5���~��  @�� P*�/~�<���R[[[�+�8?���Xq    *���T�Xo_�bټ슅�͛7  *�� �R���Igggn߾�^MMMZZZ2::�J426�׳��5    �T�/]ͤ��y����p)�'�x"  Pw  Jg׮]�����hmm����P��oYד���     T���9i�}A�a���)�G  ��  ��Ν;���gbb",�b����6333�D�����ky�ч    Pi��x%Sz>��TC�nݺ466  �@� @)mٲ%G�	K�X�)"�J^q���@���MC}]     *���DN]�毾�>���)��{.  Pw  J���ϱc�*ve|�kkk���}|j:G.]ɮ�    �R������Ά��������tww  �B� @)544�=�����^��^[[[� 8z�jv<�P���    ����z3,L5�O?�t  �L�  �ց�_�",���֌���RMLM����ٳ�     �t�����>MMM)�b�g��� �2� PZ===s�r�����Vс{�X���|dmZ    �R�˹�Caa�;��۲eK  �l�  �ڮ]�������ܜ���LOO�RMM�����o�     �T��d�z�������jjj�{��  @�� (�'�|2�|�I&&&��kmm����������1     +����\�q+,Lcc��W��_�>���  �ǿr (��y�#G������V����L�p�r�o},     +͗���}���w��  @	� (�����رc���	K���infjj*���������t�6    `��6<����yP��www�} @	� (�"�޸qcΜ9�^��~�Ve?�;;;�C�rpǦ     �_�W��444��jjj�o߾  @Y	� �
/��bΞ=;2��Z[[+>p/��v3?ذ.��Z    ���Wn���+�z{KKK֭[  (+�;  U���z�\�|9,���ƹ%����T���_���kOm    ������8eܟy�  @�	� �Ŋ�����Yq_mmmJ��pchn顮r_~     +[�����ݰp��ͩ�/oS��lݺ5  Pf��=  �'===����͛7��*K�^����yg��     <3�����H����;v8� ���  T��>��կ��*�p�՘���T��Gs���l\�*     �۱�k�S�����.O?�t  ���  T��{,����s�NXZŊ{�B�⾡�;�55    �_&��s�╰8����զM�R[[  (;�;  U��g��o~󛰴����7o�F�&r��Zv>�6     ��.\���Y�2�����d�޽ �j p ��<��S���2>�ץT__���挍����kW����M    ��+�7N\�S��K�e������1  P�  T��۷�СCai�e	��'��޳�     ,�/�dfv6,N��^[[��z���  �B� @U���Çgz�S�K��3[�K����d��k��d    X>7������a�:::RV===�^� ��L� @U*V\�x≜<y2,��	���֌����gf��������     ,�b��ū��OKKK�j߾} �j"p �j8p �N�*���JQ<[���p��`v>�6=�    Xjn���[�a�ʼ�^���Y�&  PM�  T����<��ùt�RX:��X˙��J�����y�m    XJ���W筷߫2�{��	  T�;  U�^�����3,����ܺu+eqyh8�7o��U�    X*���֝��x��JCCCʨ��6n�  �6w  �ڪU���ӓ7n��S<�Z����Y����=;SSS    �{55=�?\��M��۟z�  @5� P�^|����K���>MMMOY����+�ٲ�'     ���+�;1�$)Wʨ8g߱cG  �	� �z�֭�[xK��T(S�^���<�fU��j    �Xw&&s��Z�7mmm��-�y��͛K�� ��� ��ڿ���1,����fvv6eQ\:�x%�l\    ��:t�r��g½)�kʨ۟{�  @�� ��ڴi������hX�|���w����y]Oښ    �P��w�wu0ܛ����3�2�� @�� �������{/,�2~h`zf&�����;6    `�~�w�T/_>(e^o߳gO  ��	� ��mݺ5}�Q�޽�FKK�܊���t�����l[ߛ���y�    ,���n���r��<(e�7nܘ�F/� P��  �<��s�����)V�o߾�������ճ;RSS    ��353�/���{���T��8o޿  ��	� �?عsg>��3+�K��������ȝ��|=�֯	    ��9|�JF�'ý+�z{}��  ��  ��ݻw�w��]XsK:)�/����5����    �#c�9�5ܻb�V)���z���  � �/<�������3>>�Fq�088����ʡs����G    �m>?۟��p����RWW��y�G��b   �;  |�]�v�O>	K��o޼����]�뿚-�{���    �����p.ܸ�FgggʦXo?p�@  �#p �o�{��|��WVܗHq8_�ꌌ��lffg�ɩ�y�m    �����ߟ�K���>---)���ק�و
  ���  �œO>�/��",����R�[`ʆ��     �щ����FWWW�h���  �D�  �b�޽���399�]cc�����D���������    `bj:__��F�Rh1�R6�֭�{  ��;  |���ڹ����*,���������s���`ú     |q�?�S�aix]]]ʤ��8  ��	� �;�۷/����T�wE�~�����Φ�������!    @��9z7���s��A���L٬Y�f��  �sw  �Ŋ�����"w�]�FS�쌌�����g���Kyi��    ��gg.�v��A���OKKK�f���  ���  �G�<���ǭ�/�����+7�m]o�vY�   �jt���\�U�3����+e���[ʟ  ���  �G��e˖;v,ܻ��ƹ�����է}����s��    @���W���*�S��?�a  �o&p �yx�r���LOO�{W\Fܸq#eucx4'�g��k    T�C�rgb2,������եLV�Z����   �L�  �P__�'�xb.r��������MY}~�R6�v���!    @�����������J�8p   ��� �<�������jjj�"��������t~�w1wl
    P~�������z<��LKKK��z;  |?�;  �Sccc�mۖ�G��{���Q���p��`�X�:��.��    �'���ȵۣai�q���^  ���  � Ŋ�ɓ'355�M��kbb"eV�6�������    (���|yn ,�b(�L֬Y�իW  �nw  X�����ر#_�u�w��č7Rf�w��������p    ����̥�OEYjmmm���K�8p   ��� ��߿?'N�(����P\Pfvv6e��������jm    P�n����`Xz]]])�u�֕�g ��"p �*Vܟz�|��������E�###)����|r�|�|f[    �r(��>��^CCCZZZR&/��B  ��� �"�ݻ7����d�7�����C�9{mpn�    �|G/]��ѻa���e��#�̍�   �#p �E(Vܟ}��|��'��K<���K�}z�b^ՙ�z�   @%������W��Y����y�� �¨*  `�v�ڕC�UE���:::���xwb2_�Ⱦ�    T���.fjz&,�"n/Ff����y  �O�  �`߾}���½immM}}}���Rv���eӚ����-    T�����XeZo/B����  X�;  ܃;v����}�ܹ�M��~��͔���l>>}!���>�4-    P9�ff�Yߥ�<�1���ƔŦM�J��  ��"p �{T����?�s�7���������hN\����    �89��aytuu�,�������  X8�;  ܣ͛7�O>���HX��ֶ����=~q�?��v���!    ��74z7�������0��^[�lI}�,  ÿ� `	����?���T���r��쬚�}bj*����W�|"    ��V��~�w133΀�K������  `q�  �{�ttt����a񊅞��挍����~3��-�    +ױ��v{4,�����3��عs�ܫ�  ��� `����������{S\bTK�^����<�՞��   �J4:>�C���)^�,K^__�ݻw  X<  ,����g�������:w055�jpwb2�?s1/l{<    �������	˧���駟��v  �7w  XB�/����Ά�+V�o޼�jq��<�fu^U�K    (�SWnd`h8,�b����1eP�E�  ��;  ,��kצ��7׮]���ޞ��������N��}��4��    x����8��WWWW�b���  ��  �ث�������W��/^�|k[[[FFFR-F�'�����ۼ!    ����鋙��˧��an��ZZZ�cǎ   �N�  K���;6l������uvvVU�^8�-{WemW{    ������0x+,�2���߿?  ��� �2x���������LX�b����9ccc�����N��O�<��ښ     ����t>��WMMM:::RE�_�   KC�  ˠ��1۶m˱c������n�ˡ�y��    ���]���TX^�+����)�_|1  ��� �2)�O�>���ɰ8���sK���;<|�r��NO{k    �����휽v3,�b��z����  X:w  X&����ݻ�駟��+V|nܸ�j23;��?��zv��T    `�MM��Ӿ�a����ύ�T����<x0  ��� �2*����:w�����֖���LOO�����#����    X~_�����DX~eYoߴi��K�  ��� �2+�[���1���a������Ƚ�|y�?z����    `�\�=��W��%����%��ͩtuuuٿ  ��'p �e�q��tvv�֭[aq�����Uۇf�����sy{����    Xz�9�G�.�H����ݝ2xꩧR_/� ���_�  p����������8���ioo���p�M�u|�Zv<�6    �����@n�˯��1����t�ϱ{��   �C�NU�  ��IDAT�  �Aooo֭[�˗/��)V�1p/|�w)�;��Z���   �JRL����ٳ'  ��� �}��k��o��o<s�H�S�mmmM����ɇ����۵#��5    ����L>:uޙ�}RWW7�Rg�+~�m۶  X>w  �O�C�M�6���/,N��^��{����x%O?�.    �����K�}w<��z{MMex���  ,/�;  �G̹s�2==���1���K5��|^Ց���     �704�SWn���Ë�J�z��_�>  ��� �}T�O=�T:�����}ff6�9q.�����V��    <(�������p�tuu���6���_  ���  p��۷/Ǐ����o���e��FC�w�չ����H    ������ܙ��O�W�G}4  ���  �b����?��ð8Ŋ����S�_��GVw�.�)    �o�쵛��)������S�s�^x!  ��Q�A  @�ڹsg��⋌����kmmM]]]���S�fgg����_�>�����    �����puww��mݺ5���  ��;  < ̯~���p555s+�7oV�����x~�w1�o},    ����ԅ�OU�hƃR��466����ū�  ��#p �dÆY�vm�^����=�n����L���ky��+���
    ��N]��K7o�����{��Im��4 �~� ���o��?�yUGڋU\(�����})����_�>���   �7���g�����Ԕ���T�����ر#  ����  ��x�u�֭9~�xX����gvv6����d>9}!wl
    �犳�ߝ<����p�Z�*����&/��R  ��O�  Xq@~�̙LLL������[q/"�jv��`����5�}a    K����\�5���ƴ�����[�.k֬	  p�	� �����������������HU��>:u>k�����     �}w,_��_�����  �`� `ؾ}{����ܾ};,L��^,�{5���G'�絧6    ����l~s�\�gf�����0��f%{ꩧ���  ��� �
��(��n�/�/F��>::Z���7�r��Z�?��\    �ۗ�28z7����^���>�l  �G�  +Dooo}��\�p!,L}}���Y߅��jϪ��    @5α�k��+�j;::R����  ��� �
����g?�Y�����+��dzf6���O��L]mm    ���ON�w'��K�F����^�:�=�X  �K�  +Hccc�y�|��aa���>::�jw��X>뻘緸�   ��|t�B�NL������kjj��+�  x��  ��<��s9~�x�ܹ�Xq��������l��
    T�c��rq�Vx0����"�J���Wt�  e"p ���_ί~���0imm����g�=;���    (��U�/�����.����T����/  X�  �mذ!����~�zX�b�]��o�'����y����    �ezf6�9q�_�;�J_o߻wojkk  �w  X��x�����?2;;毱�1---�{�nH����+���u   �2�����u������H�jkkˎ;  �w  X�:::�e˖�<y2,L�$p��/��g]wGz;�    erq�VN]��J_o?x�`  ��E�  +��/���g�frr2̟�?73;����O��LC}]    ��NL棓�ÃS[[����T����g�ڵ  V�;  �`����������)�������x>>}!/m<    P�fgg���3>5�b��8ǮD��]��   +��  V�;v��/����p�����477gll,���+7�pwG�x�'    PɎ\��˷��>HE ^�T��۷ϝ#  +��  *�o��w�}wn���+.W��S���ٞ�7    T�#wr����`篕����ؘ�{�  X��  Pz{{����̙3a��w+�njz&;��wmOmmM    ���[�=q.33�@�"l���N%����K/�T�q>  T�;  T��_=?��O399毸d�|ٚ�t}x4_��ϳ�	    T��O_�����*�]+5_�vm}��   +��  *DqY��/�׿�ufg��WSSSZZZr����'�p9������    �'/_��k7ÃU�UwuU�b���k  V6�;  T��[��СC�W�		���oO��O��L[Sc    `%�9z7�?��U�VU�z�3�<��F�  ��	� �¼��[�ۿ����̄�).,Z[[s�Ν�'�S��Ѿ���m���)    �orz:�;�ig�\]]]Ů������  ��'p �
��ё;v�ȑ#a��w��_�~{4_���s�    �D�;y>#c���[�zujjjR�^}��   �A�  ���������X��������ett4��#��dmW{��    �$G���[������`�D7n��� �� p �
T[[;�6�_�*��W�gggß����j��_�   �����h�<�V�J]o������  T�;  T�6d����S,+�###��MNO���}y�����    <HS�������X�2+q�����΍�   �C�  �7��_��_gzz:�O��>::j�����O�.f���    Jqv����+C��^����[�  �,w  �`���ٻwo>��0?�s�����D����h��    �×�f`���J���8w�Zi����^{-  @�� @�۵kW�9����0?�jO������>:u>��[���    ����ɡ���Q���۶m��0  � @)���y��w��T[[����ܺu+������h_�yvG��    ����T~{�s����)mmm�4���o߾   �I�  %��ۛ�7��ٳa~��}xx8333�/ݺ3��N����    ˭�ڋ����dX9zzzRijjj��/��   �I�  %��(?��O39�h>���>44�ٙ��y��=�֯	    ,�C.g`h8����iiiI�Y�vm}��   �K�  %Q�����|��o߾m��;|z�Bz:����    X�7o��ūaeY�zu*MqN�ꫯ  �lw  (�;v����߯x����+7o��lzf6�r�t~�gg��		   ����oO����lX9Z[[+r��駟NSSS  �ʦN  ��y뭷���V�穣�#��Ù��
߬�d|�h_�xz�܇    `)L�����g2>�ln����I�iooϮ]�  T>�;  �Ll��?ȡC���+�����\�~=|����|q�?{6=    X
�;y!��w����ٙ���T�����_  Pw  (��>}}}	߯��mn�}||<|��/\����<�fu    �^�t5��+K��^]y�۶m�2  �A�  %���8���������ˏ+W���������Ҝ���    �b\�W���S����ե�477ύ�   �!p ��*Vv�՚cǎ��W\������]O"�陙�����ɞ�ij�'%    3:>�O����lXY���W�_{�   �F  �{��s���ܹs'|�U�V	�硸�|�h_�xz�ܓ�    0�x����d|r*�<�hJmmm*ɦM��f͚   �"p �+.#�|����̬E����А��������604�/��gϦG    ��ѩ10�g�����$���s#/  @�� ��֮];�b����_�������.gu{K_�:    �]�^����n�����'�楗^���y  `~�  P^{�\�t)������ե��+CCC����Ĺt�����%    �M.��saejnnN[[[*ɣ�>:�  ���  �@�b��������+�����t�nS�3���O�'{v�����    ����|x�\f���b����������_  P^�  �Ś͆r���jjj��ݝ7n��W\R��/o<�u�w    ��ټ�L�'�����ޞ���T�^xa.r  �˿� �����[��O�����݊��۷o�]��@�����<��    @��28r7�L�X��իSI֭[��<  @�	� ������W^�����7|�U�V��իa~�p�rV����5�   @u;r�j�������+�uuuy��W  ���  �̦M���C�ʕ+ỵ�����9ccca~~{�l�Z����%    T�?����U��tww�Rk����Kccc  ��� @z����,����+�a~��g��_��_�ٙ�r   T��w����3������Y��s�b�R��m�  T�  T�b��������w+~Wmmm�3:>���T~�k[�kk   @u���ο9=�_V����tuu�Rk��z  ��!p �*�s��=z47n�߭X�s�Nfgg����o���+;�    �733�����[pge��驨u�ݻw���5  @�� @{�����<333��O��FCCCa��]��C�yf��    Pn����˷�����Ғ���T������?  P]�  PŊ՛�{���O?߭�H���T��/�����)�֮    �t��՜�V����T�be�G?�Q  ��#p �*W<���ח7n�oW\��Z�*׮]����"�ގ�    P.�7o狳�a�+F<S)v�ڕ���   �G�  �w����s��ߣX�onn���X��陙�w�t�yvGښ*�   ��v��X><~6���ae�����Օ��bwww�y�   �I�  �E�/��B����݊K��~�Tuwbr.r{�����   ��6>9����ebj:�|Źf]]]*A���  ���  ��}���8q"�/_߮��a�Y����0�#w��3y��'RSS    *���l��h_F����W�ivuu�����{M  �^w  ��y���������d�v�󸣣����	s��P�8۟=�	    ��S�s��h�������Z��   �M�  �?Œ�+��������l�f��E�>88�����ܘm��   ��r��@�\u.V)���*f���.?�я   p  �̦M��裏���uttddd$a�>9}!�-�Y��    *���C9t�r�555���I�8p�@   p  ��[o�����g�nժU�r�JX�����������t�4   ��mp�n~{�\��+�ū����G�O<  ���  ����y��������577�=�{�Ν�p�S�y��鼽k[��y
   �Rݙ��{�Ogjf&T�����������W^	  �)  �o�裏f���9}�t�v�W��ݻw3;;nh�n�;җ7�ޚښ�    ��L#�O���d����sC&���_���  ��_  ��z��W���?p�͊%����ܺu+,Ε��|x�l�x<5"w   �cfv6�;����+I��d{{{*�ƍ��V   �#�;  𭊅���~;��������Օ���LMM��9{m0mM����,   ��⣓�304*K��^	�����  ���  �w*.Cv�ؑ�G��oV��www����a�_��֦��|dm    x�>?s)}WCe)^�ljj�JW�����ks#+   ���  �^/��R.^���akMߦ��-###��Y�Ŵ55���    �`���#����R��W�N%غuk֬Y  �o"p  �����/~���̄oV\dvv6,N���ؙ���֬�l    �ץ�����b�<===����J��ښ���  ��� �y�����ݻ��矇o���0��[���M��佯O���;���    ��w���3*PSS���d%x�7  �]�  ���ݻ7}}}
߬��+������
�7>5���d�yvg���
   �܆���ޑә���c%Z�fM*�~���1  ��   �w������df�E�7�����իs���poF�&�"�?�=�u�   `y�ON�ç36i���x���� {��	  ���  ��֖W^y%��^�f---imm͝;w½)����Ѿ�������   ��553��������Py���jժ�tuuuy��7  0w  `��lْ�'O��ŋ�+�ccc�����[����غ1    ,��������\����7��+������ύ�   ̇�  X��������ܽ{7��b��xr��͛�ޝ�����<���    �4>�7n��T�ŋ�+݆�y��   ̗�  X�b���λ�;���_������h&&&½��l�\����    po�ȉ��2���̭��t���y�W  �w  `ъ�ݻw�/��l��չ|�rX�;y.-�yxUg    X����9tޙU%[�jU����o�97�  �w  ��<��s9w�\�_jjjJ{{{FFF½���Ϳ>�7�ޚ�]� ��ٻ�/9�3��w眣��X�!
!$�P ���?p�Ú��0��$�s@����\������P���:��>�խ�9����} ��|:4��,_I������ʅ�   ߖ�  �iO?�t���G����%�8�����f��������������Z_    |3�����";7,_�������-���   �.�  �M�����<>��do��c6��_~r&����h��    ����d�{�|d���嬡�!jjj"������ݻ  ��  �b�ڵ�~���p�B�����cbb"�����1�J�[G?���*   ��665�;�L&X��A�d�|��#�De��:  ��  �&�������Bn�Qkkk���Ɯ��f|z6���I�U��   ����T�u�lnX �[�'����ƍ�[n	  ����  �7���{��K/��l6�����hll����`��LN�[��ƞ;7GyYi    �T:~�ə����������b>�����z(   n��  �W---q�������555�&ܧ�&fͧ�c�5ۻ���%%   P�R�Lnr���L�����Dggg�d�ɓO>   �A�  ̻��;.^���%�Q�*����`~����{��ǎ;6��  ����f���chb*X�������2�Ur����?  `>� ��o߾�����F*�
����:���c||<�_WG�w�/�C��   �b���ůN\��1gO����"�53�%����   �/w  `A$/�J�W_}5���/K.����"����\�`T���}�   @�����:<�$/��m��9�]�  `>	� ��bŊؼys�:u*�����hkk����`���:5��mMw    �?��������Ԕ���v�����  `~y�  ,�G}4z{{cl�Ԩ�WSSuuu111̿#��&�o^�    ��K�q��0�B�D㭭��϶l���L   �O�  ,�����?�t:���jjj*��l0�~�J.r_בߗ�    7�T����J_P8:;;s[ �UKKK�w�}  ��  ��K&�?�����o���\�W�%U�_�~=����oO]��X��    ��l�`��ܕ�p444��T�U2]��'�  ��"p  �ڵk��n��'O_VWW����/�_&������wl�   �|�`�^�^P��ʢ��=�ٮ]����2   ��  X4�<�H������p�e������f����"r|��X��    ��������LGGGn�c����;���+   ��  XT���G�J���J&3577���P�0��������m����!    ����G�7�.FV�^P���s��U�o߾=   ��  XT���ݻw�k��f���ihh�����$wF:������]�6EW��   X~z����(���������"v��   �A�  ,�U�V�V�~��������EOO���3I�~.vo�5��w"   ��K���N���$nO�<棒��x�'r�K   ��  X��\�z5��*//����N*��_=���m"w    ���܈�N\�LV�^hjjjr��Q��{ߋ���   X,w  `�8p ~�����l�W���199333�M�s��w�m��   ����s��3�lPX��<��񮮮�6N  ��$p  �LEEE�ݻ7~���Ŝ��_���}}}~.l&��_~r&����h��   �|sml"�9v>�q{!jkk˝�棪��x�'  `�	� �%�����sO��O
����2���bdd$XXI���G��ɻ7GSmM    䋡��x���He2Aᩮ�Ν�d���={���4   ��  Xr۷o�+W�D�W�����T���k:7��l�{s4TW   �R��_=�iq{!J򮮮�W��{o���  �R�  ya�������s�������鉹��`aM����NǓw��Օ   �T�'��-q{A������L6V�^[�l	  �����  �����ݷo_��'?s���+��444,�\���\�^W%r   ���L�}�\̈�Vmmm444D>�����{,   ���  �ɴ�x ���௒ˮ����o|z6���L��֨�   �hlj:���lLͦ�����|TRRO=�T�5  ,%�;  �W�n��.]��W����===��f���\&������E�   �������(++�|t�����dy  ��� ���L	�я~db��H.�ZZZbpp0X3�q��S�����P]    eh|2�:v.fR�p�����Ѻu�b���  ��  @�IV�:t(^x��d2��˯$�������l��t.ro��   �ohb*�:z6f���
Y2����=�Q2���G  �|!p  �Rr��k׮x��7cnn.�\kkk����Q2���OƓw�M��   0_���<z6f�����3�����ػwo   ��;  ��֮][�n��G��K.����ڵk��N�㍏NŞ�6Gs]M    ܬ���x���H��^ccc���F�)))�'�x"��u   ��  �k<�@.����>�\�������D�xr��ǧ�m����.    �����x���Hg�AaK&����E>���r��  ��  �{����^��7�)���ӑɘ�fR�x��ĝ��]�   |=�c�މ�ɊۋA����F�I�g�~��  ���  @�K.�8/������$?���v���l:���L��vkt4��  �o���|d�sA�knn�����7�cǎ   �Ww  `YH.]v��o��f�͹ LTWW�~.7n��l:o~r:ߺ)��   �_�:�yܞu�U***r[�Myyy�ݻ7   ��  X6���[�n��G��kii����H����Jg���ѳ��6�;   ��.]�ߞ�(n/"]]]QRR�$y=O<�Dnp  @>�  ��<�/>��joo����`񥳟G�m�+[   ��]�6$n/"�������7��{otvv  @��  �΁�?��?brr2��eYsss����/���9v.ݲ>ִ5   �.��g.ǜ��h$�ѓ���&َ�e˖   X�  ��SZZ�^x!2�L�����ӹ/_&������wl�   9�{���_���ܲ��+�MCCC�ر#   ��;  �,%�2;w�z�%�ioo�����f���K֌�{�|�ۭ�ĭ��   �c���_.�ť��#���+�H^�޽{  `9ɯwV   �����c�֭q��� ���,����ڵk��H>l�ӗ"�����oZ   ���\�ǯť��1���#����Į]����:   ��;  ��=��100��"���6w�6>>,�?��4�S����U   ���?w%��ť��"�]1�|�{ߋ�.C  ��G�  ,{���G155D������L�R�`�����LܿiMnZ   P��ss����HP\�s����;�Y�fM�y�  �	� �e���4:/��Bd2�(v�eZ21���/79��s��Z�>��|h��~O��   ��L6~u�B��ŧ��-*++#�444�Ν;  `��  !��y�����u&�Tknn����`i]�Mr�qǆ(/-   �p$���9~.��Mŧ��6���"�����޽{  `9�  cÆ144~����3���1==SSS�Һ:4�?:��m��
o�  �Lͦ��c�bx��K1*++�����'�f�={�Duuu   ,gn� ��r�����`\�|9�|Eroood2�`i]�1o|t*��ks�VV   �|�O��[G�ƍ陠8uuu�"�|���F{{{   ,ww  ��<����/榹��-����729�x2vߵ9��   X~F?{��퓳��8577GMMM�-[��ƍ  �� ��t����������t�䲭��!nܸ,�d������w��u�u
   |�������1��-�XUUUEkkk�U�V�}��   �B�  ����x�g�^�LƅcKKK������l���fS��ǧ�񭛢��.   ���7r#�=q>ҙlP�JJJ���+�g������;w  @!�  +�Z�{��x�7bnn.�Yr����===E���3�t����x쎍���1   ��u��p��Rd��U�Yr�VQQ�"�q���(--  �B"p  
ښ5kr�y���?D�+//ϭO�C2���g����Ǻ��    ��ɞk��W(rɤ�d�F�H����z*w�  Ph��  
��wߝ��ϝ;�.��������� ?d���W'���䊸{��    ��Ǘ{?���[2�=�ޞO}��hnn  �B$p  ���?���q���(vmmm1;;�T*�]��t&�ݰ:JJJ   X:���?}).^�[rN��Օ���/����rK   *�;  P48�?�|LMME1K.咉S���Vk�Wbbz6ٲ>����   �I��wO������������|�v��\�  P��  @�(//�C��/��L&�Y�V9��n�}��<8o|t:vm�U޶  �b����w����������룱�1�ESSS�ر#   
��r  ��444ľ}��W^)���uuu1==�㦑��7&���'��5�3!   
���T�}�\LΦ*++���3�E2E~�޽  P�  @���z(~���}��������/�ˍ��x��S���M��P   �����:y!f�Ž��ϕ��DWWW��|PVVO?�t.�  (w  �(mٲ%�������Q̒K�������l6䗩�T���xtˆX��   ��;�?���lqB௒�|�ɓ�;wF}}}   �;  P��)����Ŭ��<����ڵkA�Ig��αsq��5�yeG    ��dϵ���O�����/���X�re   �;  P�����?�|LLLD1����]�ݸq#�?sss����1>3�_�*   ��������O�t���/$S����#_lڴ)��  ��� ��VZZ?����?�q���D1kii���٢�9䳣W�bj6ܺ���ݒ    ��d[گO]��Cc_H�	�����$?�\�����  �b$p  �^uuu<x0^z��d2Q��˻������l6�s��193�ݱ1*��   ��fҙx����6V����G���QQQ����>v��   �J�  ����طo_���Ew�����0��w�F��t�ܺ)j+���   ����t�}�|�O�^Ǘ%g�uuu����r�8���   �J�  �_��;v�w�}7���X���Dccc��Yӝ�oL�/����[7F[C~\�  @�J>,��c6��[IP���� >���(/�r   �ͻ"  ���iӦ�q�F��O�b���333�/���l*^��T<�y]��̏�X   �7g�����l�4�%Sғ�%%%K�Rr�婧�ʛI�   KI�  �w�oߞ�^~���(f����l6�_��\���ܚ��׮   �sɆ�/�ƱO��JWWW^LKO�Gy$���   �;  �WڱcG.r���b��D������܅0��K�165n^e��   �,���oN]��Cc_���5jkk��e���{�7֮]   |N�  �O<�����/���H����hii���� �]���عuSTWx�  @qJ��s�|�NN|�$lOμ���͛c˖-  �_��  �'JKK�СC���8����X544���l�������D�z�D�ܺ1Z�~
   ,��}�{'��t*�U***���+���5k����   �L�  �5*++�?�A.rO�RQ����I�|��&ff���N�#���5m�   �����ݙK���|���������Xj��ͱs��   �	�  ��de�����_�l6�(����쌞����,7�L6�=~>��[��t   ��/�~���u����@��VSS���   ���  �H&��ٳ'�x㍘�+�)`eee�Ƚ���h�M��t��ո1=�o�%JKK   
I��ߞ�WG�NKKK���-�ˈ���8p�@^L�  �Ww  �oh͚5������_��wUUUn}���p�|��c�������Q    �ar6�?C�S_'�И�XjIԾw�ި��   �9��   ��w�7n܈�?�8�Uccc�R�������Ň'�񭛢��%*   ����d�{�|.r���LL���Z�%%%��O�G   ���   �����###q���(V�ī�����Ǎ��x��S�����!   `9�pm8>8s92�l��I���������~<�@�   �	�  ��'�|2^z��b�\�uttDoood]&/+3�t��3�}��ضƥ*   ����\|x�7�}��MtvvFee�R�����cӦM  �7#p  ���y�x�bll,�Qyyy��?w����}�p5�����뢼li��  ��2���oN^�ޑ�DKKK���/��ȅ�w�uW   ��	�  ��d���>���'''�UUU�.������������[7F}uU   @>J>����b|z6��������֥~�f͚x��  �oG�  p���=�\.r����b������1>>,?�S��_N�#����-�   �$�p�g.G:��&***���k�_Ftww�Ν;  �oO�  p�����?�A.rO�RQ����r����L��̤���O�Ķ5�����   �Zvn.>���>���JJJray�yq)%���   |7w  �yPWW���_~92�L��򰣣#z{{���/G�����t<|ۺ�(/   X
��}�b���6�����ť���O?�t   ��	�  �I2�i߾}�ꫯF��f���Gggg������\�<]�_|x2�cc4�V   ,����x�ą����6Z[[sC(�R��1�ۗz�<  �r'p  �G�
�ݻw��Ç�2򮪪�����~�z�|%Sܓ�����ǚ��   ��p��p����H�� nN}}}n��RJ&�'�z�<  @!�  ̳[n�%v����^QF�Ʌb*�����`�J�3�α��mMwl_�2JJJ   Bvn.>���>�������V��TVV����   ��	�  ����333��e�L�J��111,oG���&�?tۺ�,/   �O3�t�������m����6*.���駟�}   `~�  ȶm�r���#G�����"��g��vep$^��d�ܺ)jL"  `~�O�{����l*��J��+V��RZZ�w����   `��  �=�����q���(6�%c����7����LN�+GN���ƺ��   ��q~`(~�Jd�ـ�+*++��5<��c��/   ��  `�=��C111�.]�b�L�J.����"��z�Ke2��o�#�۸:�JK   ��t&���|W������%}?�p�^�:   �w  �E�gϞx�Wr�̋M2I+�t
���k�5�;�l��꥝�  ��165����UCCC455-�󓭅۷o�6   C�  �H���/��rE��������6��Pޘ�W���o_�Z��R  �����P��ܕ�w��������cI_�w�۶m   ��  `����Ƴ�>/��B���E�I&k�R�
�L:o=[Vu�=�W�;^   �2ٹ��ūq��Z�ͨ���+V�&�/�M�6�=��   ,,�;  �"J"������8&''�ش���"�����p��:C�S�Ȗ�Q[Y   ����_���S7#9SK���ϥ�v��x��  ��'p  Xdɴ��{.7�}zz:�I2a���+z{{s�;���F��������ʖ�   ��]��\��t:�fuww��ԖʪU�bǎ  ���  ,����������ܓI[�����=���c&��_~r&�����V.��p   �Fvn.�\�'{�̇������Y��'q��]�  ��#p  X"I���$����(&�ĭ�rr`` ����r�J_ޘ�G����
G   �bb&�>y!�ߘ�����ظt�����cϞ=  ��r�  ��jkk��������Yt�{2y���%������;2�9���;�  �����h��R̦3󡮮.��ږ��ɳ���   ,>�;  �K.�I�/��b�E���L&���Aᙘ�����;o鎻nY%%%  @a����6y}r�ߖ6�MUUUtvv.�󛚚b�޽  ���  ����8t�P���ˑN���$Sܓ�}||<(<I��ѥ���o_5�  @aH>���S�b`�{z�Oyyy�X�"JKK���I�~���%{>   w  ������<�L���?�T*�$Y��D�SSSAa��?���x�u���)   X�._��^��t&`�$Q�ʕ+���lI��l�  ,=�;  @I��<x0~���bQRR������Aa�N�㭣gc˪����UQ�  `�Ie2q�BO��0���dr{E��l���˝ˉ�  ���   ϴ���.�~���U�\vuuEooo���p��:�[_���룱�:   X��'�7�.���L�|K΅���� �۟}�Yq;  @��  ����ؿ���?�l6�"Y?�E�^L�w1�1?���$�d�;   ��dϵ8r�jd���[r�D�K!��:$n  �#w  �<���{���^{��b�du����ǜK�������D��x�ֵQU�   �L�����K�3<�ZZZ���iI�����<�L��;�   �'ޥ  䱕+W�SO=���zQE���b2��ڵkA�|}$������GWS}   ����g.�L:���룵�uI�]UU���+++  ��"p  �s�V��'�|2��D�d-u:�������O���O���]�+���$   X��\����8���,��������D��  �)�;  �2�z��صkW���[E�'�3�L��Y�^���W��o�F<�e}�WW   �ktr:~s�bOL,�$,������{���6  ���   �����2rO�T'��'''��p��D��ȉ��-��si֔  ��C�W"��,����X�bE���.��+**rq{mmm   ���   �H�?���_���"������닙���8�ҙ����?z#�۰&����  �X̤��3��ӡр��D�+W�����O��   ˇ�  `�ټys����.��=YW�������J���q��z���÷����   `~���g.����,��|���;*++���3��   ˇ�  `ڰaC�R0�ܳE�6<����ٙ���d��113o||:���{6����~�  �9��#{�L���Ő�����,�s��   ˏ�  `�Z�~}�ٳ'>\4�{�J:��D���=�W'��&>|��h�w)  �]����N_��3����-�����I���3�Duuu   �|�  ��5k��޽{��^+��;��L"���������x�/'��]�+���4w  �o*����/���177�Z[[���yџ�D�Iܞ�%  ���  ���+W�����W^)�໪�*����ڵk.�P����W��o�F<�y]4՚�  �ޘ�ߞ�cS���x������eџ[SS��  ,Sw  ��L4?p�@.r�d2Qjkk�;r�8]��W����׮�������4w  ���|H��Ձ��rod�>$��ihhȝ�,�$n��g��\  �\yG  P :;;s��_}��H��Q���rS�������ȅ����h<tۺh��
   >7:9���>4>���3��j���������   ˜wu   $�8|�g�'?�I�D��4�dj���HP�F�s���Y�*6��  �bw��z����Hg��)���l\lIܞ�����   ˛�  �������0����E�777�&�����+���g.Ǖ��x`�ڨ��  �b313�������*������dQ�����  �;  @J��db�O��H�RQZ[[s�����bwuh4~������k���   (����>�T&��***bŊ��'�`����  �;  @�J&�?��s��K/���l����\�>99��T:�=~.6t��}�DU�#  �p%S��J��l��(//��+WFYY٢>W�  P���  �������gff�tttDLOO$�����u+c�   (4g��Ǒ=���d��=�ۓ�}1%����   �;  @�����E�/��bQD�%%%��ٙ��g�$���%��?8s9��ƿ�zK�UU  �rwcj&>8{9�G��J29}ŊQQQ���M�ݻ7   (Lw  �"PWW?��s����d��r���+z{{#�J$�����|<��veܾ�#�a  ��&;7'��Ǘ{#��X*���$n���Z���  
��  �HTWW�&����gLMME��"r���t:�H�3��sW����x�ֵ�T[   ����T����/���ߒ����;w޴�V�^�?�x   P��   E$�tL&����Kq�ƍ(t�����g2��/���+GN��kW���]��  y-��~�Ӿ8z�?7��R����3jkk��6l��~8   (|w  �"SYY���_~���BWQQ������E�|I&��#���k�����V���   ����x|p�r�M��������_��%A�����w_   P�   E���4�}��x��Ws��]�1�=�������x�/'��]�u+��4w   �?{����8~u �Lm'OtttDcc�=/�۷o�۶m   ���  �H%�������q�ҥ(tI����-r�+e���蕾�28ݶ.��  `������^���T@�H&�/fܞ�������[  ��"p  (r{����{/Μ9S�ᾘ����/r�+�NN�k��[��������4   �l:��g��䓶��hjjZ��%��y�X�n]   P|�   Ď;���>��|�^UU%r�k%�N�^������n�խ�w�  ������=1�J����hnn^��%[�x��&>   ���  ��{�'����w����>3>=o=kښ�lZuU�  0�Ʀf��D�ȍ�|���---������x��'���=   (^w   ��֭[s����[�{GGG���͹28��c�uMWl[�e��  p�2�l��?�^鏬���dj�b�����hhh   ���  �/ٴiS.�>|�p�O7������N�;�R��]���G��n]�u  �]]�MmO6GA>jjj����E{^ru������   �  �֬Y�����_�"��t�$rO&�_�vM�ο4<1�}x26t��}VGU��  ����MŇ�z�|�`@�J�����E{^�<x0*++   na  �J]]]��3��O��H�RQȒ�T�;�F�\��nY��숒��   �g����<�{=�*������E���СCQZZ   ��;   �TKKK<��s���/���L�$rO.p�_�.r��I�������q��k���:   ����T|p��gN�$6O ,����ػw��  � p  �k%��?����_���¾�������I��T��x�r�xܶ�#��[�e.� ���t&>���z}���W__������+V��ݻ   ���  ����:����=7�}ll,
Yr����md�sq��Z\�{7����-  ��Cq��՘N��]r��յh�۸qc<��C   ���  �o����#����(d��n2]opp0�ۘ���_��kچ㾍k���"  ��1:9�?{%����Ŏ۷n���sO   ���  ������s�=o��v�;w.
YCCC��M&�[%Ϸuep$z��b˪θsMw���  P�f��8��@��:Y�!Y&3n/))���/n���   �E�  �����Guuu;v,
Y]]]�O�;�E&���W����Pl_�26t�  PX����ǑWc:�X.��wvv.ʳ��=�X�^�:   ���  �<������|�AA��"wn���l����8�?�mX-u5  ,��������T�r��������سgO���   |Sw   ���[���Y���[��f�P%�{�J�ڵk"w������_N���ָg����p,  �Q�!�/�������f1��d�߁���6   ��p�
  �MY�vm<��3���<R�T��26Y�=00 r�;K~w����hܱ�3�X��%%  �L6'{��'W�"�)�yS�������mQ����IܞLp  �o˻I   nZkkk<��s��$����P��Ԉܙ3�t��bO��Ms_��  @��:4<%Ƨg��Ōۓ��'�|2JKK   ��;   󢾾>����_��}tt4
U�wuu�"�l��>n���t�}�\�nm��6����   ����t�����X�3n߰aC<��#   7C�  ������Mr?|�p|��Q����s�{�ȝy���h.�ټ�=��neT��  �tfә��ro��n��Z�u���eQ��}���뮻   n��  �y���~ꩧ�wމ���lPUU%rg^e?��r��Z\�>�ׯ���  ,��������K�1�J,g��'gA?�p�_�>   `>�  X;w��8r�H�$r���>�;�fr6�=u1N^�{֯���   ^�ȍ��121�ܵ����eZ�?���bŊ   ��"p  `�|��ߏ������]�xeee.rO&�g2���28>�?9+��ލk���:  ��7�������t<�,V�^QQO?���<  ��"p  `A�z뭹����_�t�0׻�'��E�̷d��GN�Ʈ��{튨��  ��%ۓ>��g�cnn.`�+))�����9�B�������D   `�	�  XpI�}�С���~�T*
Q2�L��B���ř��q��Pܾ�3��銊��   ���t&�}�'{"��S3nokk�}��Eiii   �B�  �(ZZZ�?�a����199�(��W�X����ҙl����㮵+bSW[.b   ��䃣�>���zc&U��(N��®���T��~Κ5kb�Ν   I�  ����������w����M:/D���I�I�>;;�&gS����q�Ӂ������%  �����8r�'Ƨg
I2E=9�H�\ڝw�۷o   Xhw   Ur������݉w�՝&���}߽bv�I�b�	�@�!��Lz�O�+g:�L���B;�m�b�1��}�U�kL�ɮ*=�9�|�RUI:ǖ�[�{����q���(GUUU_���'�<S�q䃳�?8��]͍  ����8������������u�{9O<�D�ٳ'   �fp  ��x��'���#�y�X[[�rs�Amhh(���6���t�z�����mۣ��6  `+��_�?}v!7�C9J;�m۶-jjj6��������  ��E�  �[f߾}������Z���D����������Ym�l�φ����Dܻ�7����jo�  ���/-�{��K�Q(��Ԑ������@�o����x��7�!   ��UN   n��6���������oY6���{OOOnt����l���x������Hܳ�'��苚�  �r�����σO_��B!�\����p{U����҂��>��   7��;   �\KKK����9����QWWWnV��WW������H������*�  ���j!N_΋<�VV�YCCC���oz���{�G}4   �Vp  �(�������x�7�̙3Q����r����X�Ͳ��'>��b(��������  P�R���K�yQ���9/����������+l��{,��   �[I�  ����3�Dwww=z4��֢ܴ���0���hY�|��/��^�v�}]��  ����<�K��޹��_Z�
��w===�nO����?�C�:   p�	�  Pt���������B�妹�9�܇���ܹ�f���ˍ��v�Ǟ��Mo  �U(�ŧ#��޹�1���U��GR�f������?�G466   w   ���ݻ�����������Qn�E㴵���PY��)~�s��ӟ������bwOG  @�I��?��?}v!���onߥ��=���6�k����O~��  @�p  �h����/~�r����r������ҥK���p+�����F�C�]���5  �|16�����[MjmO�����o�'�|2   ���  P�jjj���������ܹs�������~r_YY	�UF�g��?������mۢ��9  �V�81'>�"�f��z***���7��7oN���������   (F�   ��M�s�=G����{��B�)�?00�C�KKK����L��އ���-��=�M  7Å�x��`^|	[Qz����/7�kTUUŏ~���>   +w   JFj���#G�D�P�r�.0���CCC1?���[�<zۚcߎ����  �����>���s[Uuuu�᭮�nӾFCCC�����d!3   �M�  ��r�wFwww��W�����('W�!�����b049oL~��ͱo��;  #��ua|:�=w!�f,�ek���͋�S�}�������   �N�  ��������J���188�$��S�?]Ԟ��(CS3���Ggsc����{:  �U
�>:��bL͗עe��U=5�of�����Gy$   �T�  P�҅ߗ^z)�~��x����ܤ
��6� �b163G>8���;�bOOG^�  ߥPX�OG����y���b ��͹Y}��T齓ÇǮ]�   J��;   %��������7ߌ���('�Bw�=<<,�Nљ���ߟ�4�����z:�R� �o(��e>��Z?o�l�������6Kj���O~��[   �R#�  @�۳gOtuuſ�˿���|������*� ?�arn!����B����%� @�ri4���`�--pYjkO�a���fI���?�|^4   �H�  �����/��r���188央�.�ҥK��,Bq�YX�?|t.����w�DU��; �V��Z��/�Ʃ���R�=��7�U}߾}���   �2w   �Fj&{饗��ߎ��?�Iuu�W!���ŀb5��<s>����;�����*  (o��+q����ɷ���Z������7��>;w�   (u�   ����ƿ��o�P(D�H��s���\@1Km�)��qGog�7��  �%�������xp4V�h����&/ZO�͐B�/���6�  ��$�  @YڳgOtuuſ�˿���|��+ۙ������T@�[^Y�.ǇG���ط�/�7�� ��glf.>X?��th,
kk�muuu9�^�I;[������(   ʅ�;   e���5^~��x��Wcpp0�IgggTWW�;��z:si4�����o{_l�l  J�ŉ�8}a8ΏM�����o���<�@<��C   �F�  ���."���K�?�!���X+�f��Op###e�sQ�R(*���Ƹw{o���Ȼ  P��b�O�����brn!�����-���7��{���;w   �#w   ���{,�������B�墩�)7����j@)���ߟ�4���bܻ�'���Mj6 ��-��1>�4��_���� ���x���+�7C}}}^ȟ�   �r%�  ���gϞ���_��W��P>��uuu�m۶�t�R,--���������_���==QW�m+ �[e~i9>�.����J W'�"��766n������s�=��   �3W
  �R����W^��^{-���X[[�r��'���ᘛ�(E��+������ξ��o{o4��  7���|���p|:<�By̕�f����������
�o߾x衇   �w   ���t��/ĉ'����erO�{{{cbb"(U+�����p��8�m�q������  l�4������_��&�v���9ܞ�o����x��gs3<   l�   lY>�`�ܹ3~��_���b���R�.�����Mx��)���81�GkC}�=�w�wGuUe  pc�WV㓡����P�,,p}Z[[���;/:�hy��f��  @1p  `KK���_ƫ�����Q.������CCC���P���g�ǻ�.����ս�^� �Z��/��ǗF��9��K����My�{�����   �"w   �����x饗����q�ĉ�i=��������t�R,//���4����8}q$�ۚs�}{gk  ���gpr&N��G���Ƥ�z{{���i�_���*�z�رcG   �V%�   _z衇r ���^+�@xuuu�����c~~>�\���ŉ�<Z����;��* �����O���C1����K�������|����Ə�㨯�   ���  �/�0��/�����s(��f���������r35�<s>�=w1���̭���� �U��/��ǗFce���H��nO-����<    w   �+����ӟ�4�z��������Aggg����{��L�RC����ő�ok�A�흭 ��s��ə8�~>t~l2��������QQQ�������]�v   p��;   |�Ԝ�.0���뱲�堥�%o����M����81�G[c}�=�{z:���[a @��_Z�O.��G��1����koo�����4G��O~���  ���   |�;v�����կ~���т���144����lrn!�~�y;s>vv��]��1��  ��J[�G�#���P�Cl����������m�����SO   ���  ��H�������~;���(5559�>22sss宰����Z�o���aw�� @)Im�g��r[���b �'͛������vC_7��ӎqw�qG    �+x   p�<�/n��曱���.]T���������[Eju?��x���Z�����n����<_���������)��   PN�  ��ٳ'oO��_�*fff�����f���^(�
�� @1���F{{{tuum���޽;:��   ���:   �F�i���E����q�ԩܨX�R����@���r�V�� (����I��}�����>��q��w   pu�  �:<x0v��o��FY��S�{
��&������蛭�w��f���  �,sK��ɥ��xp4f����|���?jkk7�uSX��^����    ���;   ܀�;w��/�����cxx8J]j���������R���O>�cg�Ƕ��t��վ���"  nTZXwq|:>���c��K;�������F����{�'7�   �N�   nPjx��OǏ�'N�ZS����ϕB��B!`+Ka��c�y�&���qWwt�4 �����3C�qvh,WV�u��ۣ��kC_3��?���y�4   ���  �y衇���o�W_}5����544��CCC���@���j|48�G[c}nu���;�k�� |��ť8;<�\���� n�+��555m�린�/����   p#̬  `���_����o�ٳgK��=5ϥ����HY��a#M�-ĉO/ğ>��m�q{_W��n����  X-��c�qfh,���r��	�A������]�6JEEE8p ���    n��;   l����3��'�|G�����(eW��&''c||<��Ka���y��:��o�����  ��t^0<=g������X.� ����������܍�Z����hii	   `c�  �&��;r��������h������p7<<�B!���������X��t�}]�T�q� @�]\�O�����ј^X���׺��6�5w��O=�T    K�   6Qj����~G����{/7:������O!���� ����B����x��`����ή����� ����872��ڇ�f(NWv%KM����*:�v�
   `㹚   7����s�[js_\,�Fǚ��r���� �[Z�ra|*�ʊ��������TU P:�n-�Ǧr����T
����]]]]����y�F���^x!�p   lw   �IRc�/��x������Q�***���),���B!�������&󨪬���)쾫�=��? ��������L|24�G'��s�����DOOO��n��:�����?�A    �K�   n��5zjz;u�T��(�`xsss����R W/�宄ݏ~R;����z��ܘ p}R����t|6:�F�ce����a+I��lO�ՍR__�>�l^�   l>w   ����;w�W_}5�����������ctt4fgg�vK+�q��h���v��Ѳa�� �w[[[����8;4�����@i�������|�(�v�Ç��<   ps�  �-��K���G����{/jJՕ�����t/�n���7��Ʈ��������@	 \v%�~nd">��� JS�cwwwoX���:~���m��   ��%�   �������;�����_�7��-�SS���P�����[\�.��R_�����jn�� ש��C�3qnt"ΏN���r �+�wuuE[[ۆ�fooo��G?��&x   ��	�  @����m����⣏>*�� ضm[nr/��>���x���<�j�c{g[���-Q)� �i����q~l2>���e���&���7,����}�Ѹ��   �u�  �H���{�'~�����B�������D]]]����t`����J��4�G
����Ďζ���5UU D�����L|6:��L���j 壩�)7����FHϟ��<�   n-w   (2}}}��+�ěo�gϞ-�pxkkk�ʊ�L�)����xU��1���])���5��`kI���s#qa�XX���MEEEtuuE[[ۆ�^
�?��ñw��    ��+\   P���g�y&>�����oKKKQ�R�}۶m9�>??��Y-���d�|�y��6Ů������u� �hvq)>��/�����v�v(_���yQx}}���^sssnmOG   �x�  @۹sgnsO!��>�,JU
����DLNN�t+=����lhr&�cg�����꾳�-Z6& ����\^Е���Q�V������y~y�R�<>�`    �G�   �\j�{��⣏>������������=r�{)�PjR�}xj6��g�����ho]-���-��n<$ �i�P��RK�����[Z`kHa����hkkې�KA������   @qp  �q�]w��ݻ��^�K�.�lz]]]l۶-FGGcvv6��ofa)>ɣ��2z[�r�}Ww{4�� ���Ÿ81_�MŅ�(������ڼX:ި������'�   ��	�  @	I�_z�8y�d���g
�(EiK������>66V�?�����)<��Ϝ�������;�ڣ��9*+* n���ZM����ߤ�G'cj~!��+5��yc������Ǐ~�����   ��	�  @	ڷo_n�����܄^����s�`xx8��R[��󨮪��������;Z�Q�; lay%�������ӱ����VUU�����ظ!��cǎx���Bk   �4�  @�J���������ĉ�������:bbb"�x��r�0�Ԝ��ܘ��;:��o7lH�& [K���ӳ���ߖ/ƧbrNK;���._)ܞ�7*���SO��&   PZ�  ��=��Cq��w�o~�nsooo�m�###���@qI�hF�g�x����������-1��]-Ӱ	@�I��\���cp},�hi�.-�Ls����y��۷km  �&�   e���9�����{q�رX]-��P
��v�ԟ���x�v�+a�q!jk���9�[b[Gk4�� [���rO����}n�c�oSSS�[��|�F��l���	   �t	�  @�������_���RTUU�����166�[������4���{-Q[�H�r���#�s�����T�����hii����iZ��;�����   e�U%   (3��^�ӧO��o�+++Q�R�!�,��ñ��@i�YX��������ln�����oo����\��ҴZ(���l�M������_,J��;�;R=�Ӽ�F566Ə~�����   �<�  @���{bϞ=��o�_|Q�M�i��������� JS��3:=�������2��Zrؽ��):���X
��L����l\����X-�޹%P��ꢯ�/��nD
��ݻ7~��    ʋ�;   �����x���O?�#G��dzn~���m�###Q((m+��8?6�G��͍����U轪�2 �5���ٹ�����}6��܈4�kooߐ���������i�   ���;   l��v[�ڵ+�|��8{�lI���m�o����177@�HA��L#5��6����ii�z�h��� `s,,��]6��f���ͭ� %�������7"��?��Cq���   P��  `�HA�g�y&���_����(5UUU9133ccc�ܡL�Pe
Z�����|_s}]�v����[Mu����_Z���hj&��g��[�����]]]yNz��������   �O�   �����x�W�w��]|��Q��v�)�022R�A}���,,�G�i��[��r�=�����(�𷤝{&��
�M����R l�������ɻq݈������;�3   ��A�   ��Ԝw�СػwonsO��&�%RXzz:�����uL/,��ɥ��qMUUt47DgSC��6G_{K��x��zR;���|��\nfO��+p3�E����9�~#�^�=�\��   [�w   `K��_��q���x��J2$����U����b [�����v������|_cmMt67FWKc��6�������r��Z��ٹd��_�83�ف['�Sk{SS��N
�?���gϞ    �w    ���w�uW��7�����(5555100��������$sK�176��.�^����ֆ��ji�M�)������P�
��7��1:���=5�;��Ecccn\����ݻw��*-L  �-K�   �����������s���;�������-r��Ғ�R��Rtrn!�3_�WSU����Ҕ�񽥾. n���jza1�G�fcd�r�}�P�b���]]]���zC���O=�Tn�   �6w   �k����~�ȑ8{�lɵ�����6���>55ZM�ﲼ��&g�"��[뢭�᫦�|��"
l�o6��������Uav���Pz
�WW_�e����������    p   �J
'<��3188o��F���E)��������Hm����p�R�}tz.�+M��W�j���>޻��r�{CmM \��啘�_ȿ_R�=ڧ�-�JN�suvv��nDj~��g���>    �p   �U���+q�ĉ�ӟ����QJ���b۶m1>>����WjX�YX�����W�7��D[c}]-M����u9�l])�>���s��}�򢙙��_��(})����55׿�/�՞x�رcG    |��;   �w=���q�}��믿�[�Kɕf�������� �(sK�y\��^�h8�W]Um���P�U�=}�\_������L�/���|nb���|�\?����e#Z��k�~�����Geee    �-�   �UI-}/��R|��gq�ȑX\\�R��۷o��������Ͳ�Z����<�ReeE4��F{c}�75\�7����������A������[�;:��ف�`#Z�[[[��g�����    �.�   �5ٽ{w�򗿌w�y'N�:kk��Jm����###��� 7K����i���B��ښ��ޯ��;֏5UU�<K++1=��C�s1�����t��QR�z�C�Hk{uuu8p ��    ��   �5K!��ƾ}����_����(%uuu�m۶�䞆�p��--�qqb�k���TGs}�������߷/�k���3Ky��t^tr���# ����===9�~�v��O?�t�C   \-w   ລ�����ş����農��"�����H��E�6��� n��s�����c�u�_��S����1��������斖�
�� ����'L�-���j ��R���+Z[[��5�<멧��y   �k%�   ܰ��/o7�ȑ8{�lI5�������@nr���m�@�(�����2������ʊh������M��9��T[�o7��)U�)����w=�M����ا�����\�������������~<�@    \/w   `C� �3�<�������6fgg�����}�澰� �,5X��oߦ��:��Gcm�W�)������6��fJ7ҮWB�)����q
�ϯ�N��P� ;�ƪ���m�)�~�����駟΋�   n��;   ��R���_���?�=+++Q*jjj��?==���Q(�\�q�siQ��_}���"R �.�kr���.ꫫr8>�S@�^<W!��/,_����������]LA���ʞ���jii����r�i���Ç���7    6��;   �)�����{�ȑ#q��ْjZM������>?? [Q���ڳ�����������h���������>௄��ǵ�I�Uė�Z�_Z��F�W
�ǥ���K���_������ (*i�ojmOs��������   ��$�   l����x�gr#�o����Q*��������9���ۭR��pU!����Z�k�*s�&�禀|uUU>��k�/�_[U���iԬm����K+��c%ԗV�o�p�j�?���r`==���Ws��PB�� �������^YYy��M�v������   �=�   ��K��?��O�̙3��[o���B������������v�ƤP�\j����W�O����c��J𽺲2��t_���]ݗ��5_�_��c��</=��2��ؤ0���JnL_Y-��k��j��K���5O�IǕ��Ǥ�.�ϥ�/����W�})��b���SWW�[���Z���in�1���   �fp   n��o�=�'Nğ���X]]�RPUU�C )̑�ܗ��~C1 �#��WV�n��K�o�������7�V��W]��-���_o:_K��o�˯�`3���J����A�kU[[��n�-    6��;   p�=���q�}�śo��ϟ�R��ܷm����y��" �mq��C� �#�J������~i8���8p�@�   p3�   �D
����122���Q
R�a{{{�������|   ����loll���yO���駟�s7   ��I�   ��R�����ԩSq���X^^�R��"}}}177���  p��pzkkktvv^W�z
�>|8z{{   �Vp   ��޽{��{����w��G���Z���H�����155   �JCCC^D\[[{�ϭ���Gy$��    ���  ����:>�`���1<<� }ߩ���9FFFbii)   n����<'I���*5��ڵ+�Ů��   `�	�   E���%~�ӟ�g�}����cnn.JAjIܶm[LOO���Xɴ�  �+͟���r��Z�����Ç���)    ���;   P�v�ޝ�ɓ'�رc���� Ls�}vv6   6Z]]]twwG}}�5?7�>��OD___    w   ���۷/��ݛC���_��B!�]jOLm�)�>::Z2�|  ��UVVF[[[tttDEE�5=7�:�����w�    �J�   (	)ı�����������Ν����(v�Mq۶m199�G)|�  @qJ��]]]Q]}m�y��{�7y�    (v�   @II���=�\LOO���K��>4�Z���se||<fgg  �j���Ewww^@{�v���ʋ�   J��;   P�ZZZ⥗^��/Ƒ#Gr�إ�Ş����������R   |�Լ���mmm������8|�p466   @)p   J���@���?��?�8���?���B�Ժ�m۶����A�B�   W�]�������r���=��S9   P��  ��p�w�q������+++Q욛�s����d   ����������������k׮    (e�   @Yٷo_�{���[o�G}kkkQ�*++s�b
��6����   ������؞دEMMM<��Cy   P�  ����!�����Ĺs�>�B)}}}177����@  ܸ�赭�-/|�������ٳ'��|   �\�   e���>�{��#G���x�kll������������  �/����Օ�^��ߵkW����   @�p   �^www��?�c�����b�+�����ԔC����  �����<OI�r�Eoooޭ*�    ʕ�;   �e�0��~������㭷��-�Ŭ��*zzzr�=�򗖖  (]�?5����\���\��'�̍�    �N�   �rv��?�����O?�w�y����q۶m��}||<VVV  (���y�jGGG�}5��N���9؞�   �U�   [�m�ݖ��ӧ��ѣ���Ŭ��)s bb"
�B   �-��wvvFu��_�M��'�x"?   `�p   ��{�'��'O����cii)�UjqL͏���199SSS���  @qI�S�����������Ӣ��<   `�p   �Ҿ}��HA�cǎ���r������� ���cvv6  �[���.7�����J�ݿ�a
   `�p   ��r߻wo������j�������ɭ�)辰�  �͗�������ժ���Ğ={   ���   ��Ԑ�~�����������������n� �r��)����W�����x����{�    �N�   �;\	����[o��q
�(V�}����������� @�kii���Ψ���������~���c    ��;   �U����C�Ł�w��]�;w����)h���SSS9辶�  ��hjj���X��q<�@    |7w   �kP__�>�l,//��o�]ԍ���֖�����133  ��K󁮮���������������   ��p   ���15�?��cq�ر8}�t���F1�������vOm�  \�T������W����_�   �:�   ܀\9x�`�߿?�=~�a���D1J��������sss  |�t���y�������#�ĝw�    \w   �P]]���>�hnt?u�T��S(���7s�}~~>  �������ۣ�������?�p�q�   ��p   �@�����=�[�}��8y�d,--E1�������t����  ��,�ӎG)�^QQ�M�ohhȍ��~{    �1�   6A
�?���y����'�:���ߟ��SнX�O  �,��=5��p��ۛ�����;v    K�   `��۷/�ӧOǱc�r�����4���bbbB� �����)ԞF����f�G}4�o�    lw   ���{��#�S����l����<����WVV  �IjaO���������---q���    6��;   �M��A��Ǐ���b����U�=5�� P�RX=���`{UU��}lWWW<������    ��    �ȕ����~��crr2�M
�477����t�WWW  Jɵ�SS{jlO��    �\�    ��m�ݖ���x���;q�X[[�br%�>� (W�c��ڢ���/�VVVƮ]�������    ��p   (��/���\��f�B���/�� (V���^SSw�qG8p ��   ���   �Lccc<��ӱ��ǎ�?���B�W��i\	�///  �J)�~%�����������   ��!�   P�jkk�����裏ƩS���ɓ9L^lR�{�y>�S0  n�fokk�㻂�i�fKKK�߿?v��    w   �"�:������ٳ��}rr2�Mj�LC� �����*7�_M����3~���#    �K�   ���ٳ'�������������(&W�����9辸�  ��R��Jc{
�������lO�   P��   JP����?cjj*�y�8�|
�(&y,,,�{: �����Ρ����]����;�3y�|   ����   ���=�=�\����ٳgcuu5�I}}}�� p�jjj���=����3؞X����o߾    �4	�   ��"?|�p<��q�ԩ<�����\	�/--���d���  |����������;���?�p�ر#    (m�    e���2�U�q���8~�x\�t)��֢X���FOOO!�~�B!  �����hkkˍ��&��n߾=8�w�    �w   �2500/��b���űc��̙3���Ţ��:��Spiff&�����  [SEEE455E{{{^�m�����x衇r�   ��"�   P�R��O>?���ԩSq��ɘ���b�BI����u3}_)込�  l�|0����i�I�#S�}�Ν   @�p   �"Rph߾}y\�x1�?�.]����(�����9��:��� @y����S��ۚ���۷o��<    �O�   `�_|1ɏ;gΜ����(�u>�p���*��y  nLmmm����i��=���΍��~   �<	�   la)D��O���8u�T�<y����uuu���9�>==]4��  \����hoo���&���P�Ν;   ��I�   �܊�o߾<.^�Ǐ�K�.M����::;;s�畠{�P  �[jhojj��������s��۷ǁ���%    ���   �����x��cnn.�;gϞ����(UUU��3�R�|
�/--  �%����zkkk^����F�;�37���;    $� �����X]]��}��t��jjj�   nLccc<��y�9s&�}���b��@����H�tO�w  n����lO#��}S
�www�������'    ����TW�&i����Z Ә����15B.,,��z�/��7"rR>]TI�ߦ�{���O����k��I�Bi�0��,  [��ߞG1���s��������<�(
 �͑�������jz��o��   �Ւ�ຬ�����dno�����������P����-�>S�&I!��q�L
���LGGGy;�� `�(�V������=���r�{1�I  �Y:�J�P�VY��v    ���; �*5������p}uL#��WVV��]i���Ǥ�tq&����<��N�  (W���D�B�4��*��  l���N
���ν�I[;    7B��dO��.�ŋ�1���b�Q�����Mi;ށ��ضm[>^�  �E1����UZ������N)��@  \���ޝ@g]������$d���"��	�E�E�}��V��ڱ�e��z�̙qڞZ���.ETv
HQED�N�	KH H��^�FDH����ޯs�yB�&3��w���ύ��wm��y.��     �-� �TVV���ڵk����ݰ`�W_}%x߉'\��FU�d��֭[�ѪU+5mڔ6#   �@mu���t7,%%%�6w�3  �8{���v�ׯ�ݭE��  ��a�V�gE���io[�r	gΜ9��<�_�=�۳{UVb���_��3tt�  �7� �lc-�(��u^^�kg����l��}�v7<l�زeK�i����  �`U��ݞ{7l���JHHp��ɓ.�na��@   ���Â���n�PUY8�
<z�꥔�   �O	Gii��=�n��[���x^-�^Wl}��U_=�JDl�`���� �[�@�ӹ۶ms�O��އ�`�sC�6�ݭ)33�I!   �N�v�ܰ֠��׻g^���7;dڸqcw�>�<��  �3�[���%���h�;u��m�   ��ٍ�TQQ�>|vX����׆'`_\\\�����d`mX����4�k!x  ���; 1�[;{nn������$5c'�?��37�m*edd���m"�kTT�   �``ϳ�{�v�6w֭[��{��kt���Y��!;xj�I6hu  ���y������۶�تU+��?Pll�    ȕf�����ڰP��9r$,���ކeW������.��ym֬��6m�� ���; ;�kA�/��҅����#���$=-�,P���]��ݳ���Fӹ�   ��Q�F>|�{�n�ڸq���{�c�.�,D�;  ejk�߳�^�z�I�&   �WZp�����s�v������q׮]n�+99مݛ7o�^[�hᆭ� �w p�w�>h�p����0o޼ٍY�f�)�gee�K�..�   ��mۺa����tZ�ܟhu  ��Bm����;�5F{   ��[��ؖ��f÷��ކec<lNbn�{V�g���  �>� `<-�6lp��C�	�.�Y��c'��u��6�lc�M)   ���(���ۍ��b7/�$���  ��kk�P�=�dff���/Wll�   �pa�j���矽I�u��a<������ۼ�}����֭[��L���  �� ��#,���矻ӨL��-��ނ\�R׮]]����-<   ���4:Խm!w��M��  ��kk��Gzz�z��ƍ   u���w�^mٲE[�n�Ν;]����ѣ���O�0�}�vw�_v�e�5..N ��F� ��B�_|�{����J�d��V�X�M�սW�^43   �y�����6�({������ǏwAw�*  ����			.�~nɅ=�dee��  �Pf�vkf��D۶ms�x=v���������e˖.�ޡC�j7Z �w �Cv�w͚5.�n��i�����0m�&Wvv�ٰ��t   �@�ZFm��jݺuڳg�_o����٨��PYY����   u���4h��~��Ђ�ڵs�:��   �������{vhOv�a׮]n,^��͗����Z���`0  �� |�&L"�P�ƍ݃4H,�~�z7<�����S��ݙ�   `%''k�С�m۸������'O����d��IIInX���ݭٝ��  �W�fF�a;;xW������֭��   ������Kw룽8���Z��kx��?�[`׮]���. @�!� >`M}j_�z���܇`Q��ݚ�z�쩾}��}���T3   �5jt6�~���<�o�>���,Tf#55�|�Vw�  \*+��@{bb�ق
[���7o���vc�   �Pd!v������@M����ؘ>}�[_���6hw���wc �"P�Z�J+V�p� �Y������HIIQ�>}4x�`���	   TM�4�����ۻw�v�M���Wee�_>���Q��f��6_d�  Ԅ��[������ξ�B�-Z�p�1�   �v�ڥu����>s�����%K��a�Ν;�2�.]�(::Z  � � �Ȯ���v��ٳG@(:|����kѢE�ԩ�����/����   hn�[��5�ە��`��֦j�Z�,�ns�ӧO  �|,�nm�6<7,�3Ezz����>    Y���O?�'�|���`�qڿ9v����z�r󯪇� �G* j)??�5[[c��S���X�;�l�aÆ�Y�f   �'�nϴ[�n��͛]3����111nXӪ�m�8qB   �hM�j���t��ڻv��Z   BV^^�>��cl?r� �,���ذ9Yvv�~���2@[� �w ����rwJ�>��a�N.�!�?�PYYY4h���y6�   �@T�^=u���O���/�t��#�nM��VV�|�9��;  �ǚ=�����;סC��   ����b�Y�F}�M�Xg��f�~���fw� ��� P���ג%K�z�jr���溑���������L   ��j�����r��URR◰�}>�`[ee�������ɓ  ��B���n��ƺ�YyD�F�\��]�v   Bѱc�\S�e0�������6��V�+��Bmڴ �{��l۶M,���k�`b�Ľ�3g���>\-[�   袣��3�O���͛UTT������Шk�4�v  ���x;�V5�nA���t�o�^m۶   �l�mӦM����׻5/ �ٚ�e��hڴ�������6 ��p�sXkߪU�\c{AA� Ԝ-F�ב���,6L]�vUDD�   �@W�������e�wE�?6�,�f"6��ۦ�5�[S  |�lѠAl�W[#���7V�ΝբE   ����>��C��~��Q�j����9s�f͚�.]�h���֭�� j��; �����裏\c;�*�{��k�2d����JEEE	   ��`M��6�ݻw��[ۘ�G���ᒒ�ܰ���naw�  ,UC�qqq.�n7�4o�\ݻwWJJ�   �Pe�7ntł�����6lp��q�����+--M ��#� 암����/^�'N�oj���?��_}��ns   &n{���/��_��OZH�Frr��[�����J ��g�v[���n��Z�r����   eV&h�|��:t萀pg_V��p�BeeeiРA�ѣ�� P��-k۳���L�P��P��ٳ�t�R:TW]u�{   JvK�cϹv���w��u�J�Fjj��fw��:uJ  �w<M�e����H%&&�P�]I+    �mݺյ���g�����zqnn�M�4q9�+��­� Ώ�;��STT��}�+��,lcA�E�i�����԰aC   �ȞemC�Fii�>��s�޽[ǎ��ϥj�����ݭ�  \����0{�P{JJ�ڵk��h�  @8�u��������v��! �c��S�L�;Ｃ����ꫯVZZ�  �F�@� �&��i~��$�  �P���p6�n�Ok�ڶm�����Q�x�|m�6O�8���
  ��~�Z�݆��GEE�q��j߾�233	�   lX��|�e˖�[�Nyy��J����_��vp �5� B^aa���}}��'u~E<��t�븮��w�3   �,�ֱcG7����]�}�޽�U�.Y0/11��[��vg� �wY���Y�ݮ��ז-[�K�.��   @89t萻���s�)�[�]�v�p���kյkWEDD �w !ˮ�����ŋ]K��`�!����?��O:TÇw�X   @(hڴ�櫯�Җ-[�ζAXYYYg���-�g���r����r�  ��:Tզ���T0���hi  @X�R��K���[��om߾]/���Z�h�J{����H@8"� �؆��\t]_��{�ky����j;�6�5N   �"::�5��0�����w=m]��[�ݞd�>�}lO�;�� �Pg����8�s�B�v��y�����v�v    \���kΜ9ڰa��u�n ����{������O^@����aavkk�?�ۄ�6��3gj���=z�z���U\   IU��-dna���<>|�N���a,�naw�9 
,`av�/��m�ֵ��4    ��ٳGs���ڵk	�~V\\�I�&��I+���+% �=�P����EEE�<�q��)33S��r�ڷo/    T��ƺÝ6N�>�;vh۶m����������6t���v�܆�+++ @0�\����Ҟ����eee�q��   @�dV�2}�t-Z���;��A�@P۹s��~�mm߾] 5X���U�n�t�m��Q�F   BY�z��O�!OkR���]m>v�Y]�p���6--��=�w�� ��iٍ$�s�j�Ϯ֭[��   �Â����6l�  ��j�}Ĉ�߿�[?�PD�@P��3f��� -����jذa����#    Xm�.]�0��a�wی<r�k|��a-��1������  @UU[����բEu����   ��Y�b޼y�裏X����	���[�օ뮻Nt% J�*Z�l�;=|��Io�T9�|�Z�J7�t����ˤ   a'%%E�{�v��߿_[�nUAA�JKK��Jik	��`BB���5�{��� ��ii��Av�_��͕��ō   �;v̵?/^��e0 /;�2q�D-Y��5����K *���<m�4	 ���ʜ�}�ᇺ���ղeK   �iӦnk��������u��A<����5�ڰ�}r���}|� �ڲUh�a7��P�6mԶm[   �0[����\㳭� ����+���}�|����� ;� ^aa��N��/��B p!�R���k���5j���   -��	����m۔����}���ׁ��aDSYY���w��  ��n�S�3$99�m�[����.s?_    \����^�Z3g��ѣG tmڴ�e&z��1c�(--M ��X��m���}�]�� T��C.]�T�~�������O    �f!�.]��a�6$;(ZPP��>u��?���H��ǻa,��	�۰gz @����9hoѢ�Z�j�v��)::Z    j&77W3f�О={ <ء�K|���:t����z�. ���;��dmr�&MrW� @m���(''G�|���NN&   �a��޽{������6=:��V�~}%&&�a쐻���^}�0 �/�9РA%%%�u��n�iӆ@;   p	
5m�4mܸQ ��W_}��F��>}����  XpP�������]+V�`�Wآ���iĈ��꫹�   ��sޭM=//O���:x�JKK}>_��^t��o!wϰM�  �EEE��������왙���    ^�	�ڨ��� >����^Ӓ%Kt�w�98 � �]�3q�D�` �d�vx�N&�;�m�   �8�m��c��{�����\ི�ҧ�Z}m����݆}N ��e�v�>n�v�D�ܹ��4i"    ޵a�M�:U����sٚ���g���W7�|��5 Pp�wǏ�̙3�|�r�/�ٳ�Mج��G?���   @�Y�<##��4ݱc�{�>v�***|���
]k��a�ƚ�,�~��	x�e� pa�}:::�m�7j�ȵ�ggg�aÆ   ������ɓ�y�f��X�ȪU�\	�1cԿ7��@D��_}�駚2e�� ��`a���&l����[   ��IKKs�w���ׇ�Ν;����f�s_� �'Li,`�iw��u� �;v�)..�؛5k�:�P�D   �[�����C���O ����2���Z�b���_�E͛7 � ���&N���k�
 �a߾}��_��믿^7�p�ې   p�RSSݨ���z?x�JJJ\뺯�MM			n���w���c@�������n��ܹ��6m*    uk�֭�4i�


 ��m�6������o�Q111�@A�@��k�rrrt��a�?�>}Z�g��ƍ����L���   �}~������]������� �������<�B�6,�n��w �.+�&���$�fҩS'7(	    ���P�O��իW�̙3�Ke�A,Y���&��=++K ��3�@4w�\͙3���������\7�|�$    �e��mۺ�QZZ��{��ё#Gt��q��x�6<l��v�໵�[ �EDD�����a���4]v�e�޽����    0lذ���ۺ	 x[aa��~�i���W��v�4h  �'� �]E>a��� ��,'Nԗ_~����]�   ��X��s��n��z���<�cǎ� �/DFF����6�(o�O��^9� TDEE����n�Zݺuso   <�&2c��Z�J �K��i�krss]��~ !�����g���>ۄ oZ�v�v�ܩ�����С�    ��5�7o�܍�����{�n8p�5�Y�ؽ�Z�-to��控��z?u�  �U�gdd(;;[͚5   ���駟jʔ).� u��ѣz��իW/t� �?p�36�z뭷�~�z@09|���|�I:Tcƌq�    �������j�޽ڷo�:��Ǐ{=|���X7<�e�>�O�݆� �}����vs5j���Lw+FJJ�    [ۘ4i�֬Y# �;d�}�v�s�=��� �%�Z |®�y���]� #kg\�d�����g?S�&M    0Y��cǎnxTTT���@{�����]�B����-�2ㆧ���-��	�۫/Z��/��cn���\{۶mթS'p   �v�ء	&���H �o��z��)P��n��l������zs� �%??_�?��n��v���_    ��m�ddd��a��v߽{�{���N�8���}l4����4�[�݆�[�����(w��^a���0O�-\c;   ��aks���ܹs�@@�nڴI��{�[�  _#��klSx���ڼy�  �X��7�p����.��    �X���t�Mָn�h���w�G�uW����u��Ӷl��6�-�n�w{�: �k_�� ���q��.�ޡC�o�   �l=�Zۭ� վ}���?�I7�t����*��)� �b۶mz�W�0 ��U�V�	�����Z�    �k[oڴ��*..v����B��QZZ���`����7��P�'�n!{O �^�1n��k�ݰ7�[�V�v��   a�� 'O��J�  ��:������_h�ر�> �w �l���:u��p�P�k�.������v�S�N   ��p��Ν;��t߻w��>|�l��W�[ ֚�m��j��3��qx�� ���SRRԼys�m�V�Z��f8    ��%���Z�~�  �X������]Ƚk׮ o#���l�N�X�B Nl���g�Ս7ިk���k�   �0�����;�Q��,�n�����Ǐ�u�_j����8�߫��W}���O�=>>޵��a���teff�fv�}    8�M�6)''GG� �cǎ�^���u뭷��� j��;�Z���q��iϞ=�pd���3gj����{'    ��kj>�5�:tȅ���ą����]�R������&6����s#pa���ns֚���m�7m��5�[3��>    T���g͚��r @H��e˗/�Ν;����� o ���6nܨ	&�X wve����'����q    �>��`��s����UTT����~d��'O����e���>��B��f;B�}}DEE��!��n�u��l����ccc    �`��W_}U����Pc%��?��~򓟨G��KE�@�ن��"~�w�܄۔oԨ���PPP  �8p@��_4v�X���S    PS��P�����n��eeeg��{���ǵ9��]�	�WVV������ EDD��u;�a�boذ�[�JMMu-��j    |i׮]z��ݼ B��T9n�8]s�5�����# �w �b����nM�-��g-U6�m��ܳ�mo{ެ�*>>�]�nv%�m�m޼YS�L�l���+��nЈ#�   �Uj��E���O��B!x��m6���]Y˺�m��q��JKKs�����   ���Z�J'Nt��@��u�(//O��w��@mppQ�!����+??_��gmT�a|���m���_l��:��k6Q�={���ۧ{��+_c    P]�	�;v̅�m?~܍'N� �'o�tS�P�5d۸�oYӻ��=�j;����~|�Oh݊<ֺ�Y�JIIQzz������	�   d6ǝ:u��/_. 7V��������Wff� ���� iZ��k����/��2eeei���:x�ڴi�m���&�m,�ƣM�|m�ڵ:|��~�_�w    ֘d�u�����F��G�����-o���	�_,ok�	�{T�����@`��ok��a�vd��ຕ/Xh݆�-Y�zrr�{��j    ���
Ǎ��;w
 }/|�'t�wh���� ��{mڴ�M�l���6 -�n�m۶n��t���/��m:������P �a�Uv��P�V�    ��:�����._ZZ�֒��6,_�ޮc�\7���$_��{� �������'$�ayO(�^=o��<A���m�ʚ��՚���ڍ���+    [�l����URR" w���o�����Z�j���Z�b�&N�ȕ��6-�ޭ[7l���/5jԈ�;pG�����7����:w�,    U���n4iҤ��[�����`��Z(�jS���m#�jx�s���V�Wf_���ws����x�/��<�s�����ϳn����������{�����������R���Ն5�[P    pq6�[�d�f̘!n?�y���z�ܹs�T �-_�\�v������. �b���p͞=���m@�o�^]�vUǎ]V���;�����^w�y�$    ��Y�ښ�mx���[���������m��y���sٟ;7�na�s� �6�{�/�n!����?�	�WekD>��������~�8�W�D�߳p:    ��ٜ��W�^-��ۺ��=��ږӰ���ڼ�s���y{�� ���IOO'�����|����/~�eff
 .��;���p���4j�ѣ��7v}�>g ���&Mr��#G�    ��<��6     �b�_z�%mٲE<�g�ԩ�Z�h�iӦ��zFF�Z�n��V藒����Di ���G��'�Џ�c���G �}�p�p��M����ճgO�j�J��q��pa�2:�������         EEEz���~!p4i�ą�m����k��^5k�̧a��!�|۩S���k����1b�yoD � \��g�a�����.�ޫW��^Y�l2f��^��V�X���2�w�}罢         @�۹s�^x�;vL𿤤$h�޽����2-[��?X�<�o�Z�}�ر�' |w ���'�t��Q7l�ԦMj��U(�8[}bb�JJJ��֯_�g�}V<��bcc          x�[�ε��W��X�`�Νխ[7eddl��)��O>q��_�򗊏� xp5�?��S:r��{vҰG��ׯ�kn5��N���-[����>� �4          H,^�Xo��6ae?����٭�݂����l��6�ѣG�v�ء����.?��* �C�S�w��3�<�UYu����{�V�>}ԠA�*��'�������O?�_��WJHH         ��t��iM�6M|��P��Vy����3(��� �|������ֿ�ۿ�C, @�C�|��gUVV&�NJJ��&X�pb�R�d@��ڵKO<�z�!%''         @`9y�^}�UmذA�[�Z�R߾}թS'իWO��2۷o��g�@,?���\�����af�֭z���U^^.����=z�䪦��g'���~��%          �Xy�3�<���|�nԯ__�;wV���դI����4�8˴������{]�
@�"����7��_֩S���`��\���o������         �����p��={�kذ�kk�ի�bccJ�T �WQQ�W^yEw�}�;� <p������~{ �w%''k�С�ڵkX�=�fP;�rM�=��Z�h!          �a{wO=��
߲v�>}��`����"�@͜>}Zo����!Y.@�	�' ����+''�����4h����ׯ_�N�j"""�M����+ �g-O<�|�A�i�F          �ݾl�v{��n�ZT���]� �Q�ܙ3g4m�4W�:|�p/$2��z�jn����pX���+�Ptt���w?~�]u����E          uc���.�~���7Z�j��:tP�� �5��۷O ��2o3f�бc�4z�h܁��g����_'��%6��֭�;��� |�M� xǉ'��s��7����5k&          ��{�nWDeAJx�ۇ��m�*Yi w�v,X�2pr� |��;�rss5~�x�>}Z�t������kմiS���d������O?����w|}         >����g�}Veee�wY�}ذaa{5{���Y�p����u�wr� w m߾]/���***�K����k��F�:u.�q���]v�����7�����         ��nݪ��'�=�!�����l¨���^�����t߫��իWO Bw ��ܹӝ(>y�P{����ݻ����*EGGՓ����9 �C��mroذ�          x�ƍ���/�ԩS�w$%%��+�T�=�VA�;����&���?u/ ���;B��٣�{�ŗ(33S7�pm�`��z_\\, �UXX�B���o/          �fӦM�۽�
��﯁�~}bi�wJ�X�f��Z���8H�(�$�q��=��3*++j'11Q�^{�:w�,Ԟ�8&���޽{��SO�׿��4h           ��c���⋄۽ ""Bݺu���Õ�� ����������p�֮]�7�|Scǎu߇ ��@8x�|�I����c�vkm'0z�,�y�f��ݻw���ׯ~�+���         @�؞�s�=��'O
��u�֮L�Y�f��Y���;�=+W�Tll�n��v-܁ g�O?���9"�\rr�F��v��	�a�1 ��}�v���Kz��%          ճo�>wk���ǅڳ�aÆ�gϞ4'�@ZZ��n�* ޳t�REFF�[n��A�b����DqQQ�P36��ӧ��lEGG�C���������}��ǂ         P����D���L�ۛ�֭�~����;j�L����?����뮻N Bw HUVV��_�޽{��IJJҍ7ި6m��׸qc��~�������4          �����.�~��Q�vZ�h�n�A͛7j��;�;�f�rM��\s� ?�@:s��z�-�ދ��ܹ�F����8�7bcc݉���R�y��)99YC�         ��*))�SO=���b�梢�4x�`���_���j��;�[3g�t٥+��R �w ͞=[+W���\���zwM|�&d܁�3m�4����=         8��]?��:p��Ps�Z�ҏ~�#��^b���a)// ���ɓ'���>}�@�"��O>�Ds���/33S�G�VÆ��aۼ�<��O�ք	����N-[�          ����z��UPP �LLL���^�z)""B��T�ٳG |�B�999��X��� 8p��֭[��믻¸8�ˮ���Yu+--M ꖝ�����#�(%%E         @8����+���ݻw5�����n���"�Lw���(p���z��ծ];>܁ a��_|�EUTTgW:�d���j2�?�9�g�}V�������8         �Ȋ�z�-���
��A�Q$�cd*��q��)��������t.܁ PZZ�~���Y�����k���jР���7 �طo�^}�U=��,:         ,͞=[+W���V$جY3���u�rwVh!���D܁ g'�^x�
�誫�"��gIII���r�~Խ�7jҤI���         ��O>�Ds���ǲ}����W_�������@�:x�ƍ��z��s@�`veք	�c���bbbt�7�S�N���8--M��� ����]��-D         �`�֭z���]���#G�s��B�IMMuō�O���a?rrrt���\��G�`���Ӻu�kڴ�n��V7@�����1c��٥K         ����@/���***��kѢ�n��f���u+22R���:t� ԝ5k�(==]�F���G�P�6m���/\X�4f�����Z��yny��G�$         E���.�~��q�¬�x���:t�k�X���;P��Ν��\y������X�Ǐ�*��	׀4l�0��	P܁�`�x����#��+        �Pr��)���*,,.����8;;[�/�TlٲE ��ԩSոqcu��I w ���kܸq�t1ί~��9r��w�..�@��srrt���s(         !�s��;��=��n�ͅ:�d* ������/�����wjٲ� &�@��<y�����KHH�wܡ-Z�---�imA��}��g�?����:         ���w�Ѻu��ڵ�+����e* �Oyy�^|�E=��JLL��C� ˖-ӊ+��KMM�]w��^��������Ç@`x��w����5[         zV�p�B��Y)����5d�!����_qq�^z�%��׿V��Di�@�W% 캬�ӧ痑���4h ��p���?��� 
         �8���n� kk=z�������20Ǐ �پ}�f̘��o�] w  ����W^QEE��]��ٺ馛\#8��ܷn�* ��رc7n�~���*22R         @09y�k�-//�/))Ʌ5�5k&���4�@ X�t�Z�l��
@� ����ӧ5~�xZ��G߾}u�׺k�|�RLvkȻ��         �`a����


��kժ��[;8�e*v��- �7y�d5m�T�۷��@��Y�fi˖-�w٩����Z^v�@`Z�p���u��M         @0X�`�֮]+�_vv�n��&EEE	��L8*++]I���G%&&
��p�h�֭Z�h��m��~�5��+���@�v���=��cJMM         �6m��n)�����O?��]���LX�9�B�=���ի' �E���Ǐ��^��ӧ�o���ȑ#գG!�%$$�k���;��c_�r�ᇙ�         `:tH���*��}�k��V}���w �l޼Ys��q�5 �E��I�&�	���o�Y�:uB�]�E�\[�l����u���         4�N�Ҹq�t��1���ׯ�1cƐ�R))).+SYY) ���mڴQ�.]��~��Gi͚5�7���[nQVV�Z����ݻ p�����ر�ڵk'          �L�2Eyyy·EGG��nc�/�YV�B�EEE8Μ9��^{M��\�' � �Ա��BM�6M��=��z�.\��ÕZ@೫'L���{Lqqq         ��U�\� ������Nedd��2܁�SVV�r���oU�^=�{܁:d��<yR��]�e��:���;��������'         ��B��ގoKHH��w߭&M���L��o߮��_�F���G��C�oǎ��<���C�1 x�\�R]�t�~�         �b�������˅o$''k�رJIIB�
 �͛7O;vTVV� �-�@�]����fW��=�p{���5�WTT@���.�LIII         �aΜ9.g�onMiii�Μ9�	&��SÆ��p���'�:;a����7�t�:w�,�>��NMMUaa� ���R����z��!         �.����\|�p{��|%%%z�7��_��P��u`�ԩ*..�~ȏ1B]�vM�����/�ԇ~�A�	         �+���?~�*++��Y÷��iMqqq���WYY� ��7jٲe2d� �mذA�V��v�uשgϞBx��1|f̘�nڰ         ��0e�	_������'JLLB�e*���r:tP������>t��	M�<Y�����էO!�؉r ���1슭�z�+�         �sk׮�@����$���?&�,����/ ��ԩS����#�<���H�-�M�6M��^�zi�СBx��N�6m�ʕ+տ         �bي�'
_KHH��w߭��d!�Q�]�vi�ܹ9r� �w�Grss9Y��u��Q7�p��,�n�gΜ��2}�tu��I)))         ��������L����5v�X����@p��{�.]ԦM������7� ��Z�j�[n�E����WLL��6���D �ˉ'4e����         �m�-��͛)66�5�7n�X܁�r��iw0��STT� �w�f͚��
w��{�m��~}����	w 8�_�^�֭S�=         xˁ��{�	Rdd�+lڴ�^���]����B ����z���5z�h�R������kٲe
wqqq�뮻��Y�����; 8Y�{VV���         \�3g���7�ԩS���ի�1cƨ]�vB������T
@�X�p��w���n�G�^d׏L�8ѽ�3;U|뭷*--M�Wj���ѣ�=�n�          .��ŋ�m�6A�����l!|YƆ�;\��[o��?����� �"�x�M�v�ڥp�Q�F�M�6�"���K��w��j۶�         ��***r�J����}�
�L�


4o�<��G? �"�xɡC�����+�0@ݺup.&c@��Ǔ&M�����:         ���=�7�xC'O�T��ҥ�,�L��ϟ��={�e˖�=�/�>}z�O�ڷo����J��$&&*&&F,R �mϞ=��?���C�
         ��+Vh˖-
w�[�֍7ި��܁�UYY���zK����U�^=�����jݺu
g��}��7�C��&���d�޽�f͚�^�z�aÆ         ����L���]jj�n��VկOt_#����<W8d�����Kd'��N��p�;�C���.��;���]���?��         ��>}��;�p֠A�u�]�������İ�� �����˕��, ���;p�/^����+\Y+��Q����&�b�w��:rРAjӦ�         ��ٲe�V�^�pV�^=�r�-��8�e*�����~�m�w�}p������Ds��U8�pcVV����J- t�9sFS�Lѣ�>�;         ߧ��B'Nt{L���k��@
��2yyy�֬Y�+��B]�t�KC�����u��	�+�t2D@upBK~~�V�\����         �>.ԁ�.��r���G��!S���S��?��?% �G���ݻw���Y			3f��>�.�N��͜>}Z B�;Ｃ�={*66V         ��>����+�eddhĈ.��;<�E������#��Ҍ3���,(�z�.��Ddd�RRRT\\, �����M�F�)         �\o���N�<�peي�n�M���pB�ܹsշo_W
�vxrj��>ӦM����V�Z	���pB˂4p�@w�         �غu�֮]�pe��G��@Ւ�����(�:uJ ��}Ϝ9S��w� �w��N�>�Y�f)\effj��j��7o��a���{Ocǎ         `,_1e��9sF�jذaj۶��ꈈ�Pjj�8  �o͚5.g���- 5G���e˖���@�A�3f�;a�Wj�i�ʕ�ꪫ���!         ��{��U��С����/�&,SA�o���{�1�v@-pj��ɓ�;w��5j�\
�@h��w�yG>��         ގ?�ٳg+\���h���.k��
 ��۷O}��$ 5C���E����D�w���ر��K�d]_|�6o���        �0g健��
G��k����X5���& ���w�u�;~. 5C��&�xY�=����ꫯ�qqq���WYY� ���3g�G��         Li�ҥ
WC�UFF��ڠ4=ǎӂ4j�(�>�@5͛7O���
7��������&d܁Д����?�\ݺu         "UTT(eff���w��Y�w��_W� 	�@���D�S9��֎�t���m����{g���1{k���tvg����*�(g-�H�� B!�����QAr�|>���gƙ�`5\��}]������~7��J=E&���@q����?�|6hx8wxW�^�w�y'�(��>��Ciƌq��� ��W^�e˖��     P2ǎ�ݻwGM�0!~��_e���J(�ڵkǝ;w�w��]��?�c G���C�&S6�gώ���C͕ZPlgϞ���?֬Y      ��o���N����~����RS!p��ٹsg���K1gΜ ������˗c���Q6�Dq�|UWW���� ���W_�U�V�P     P���q���(����X�hQ�PH�{�(�t ����}�˿�K �L�����_����(��>����w(�.Į]�b���     @��h/Mo/�����я~0T��ڻwo=z4�~�� ����ƕ+WJ9�=��)p��2eʔ����;w�P\���Z6ŽR�      ŕ�:u*�&}����,�������Pl���J���k _O�_����6_55^>��,�8��O(�s��ef��     �b���W_}5�h͚51����$p�b;|�ptvv�ҥK�j
V�
iz��mۢl֮]O>�d�pK2�;����x��gMq     (��۷���ts��/�0�cܸqq��� ��w��],Y�DK_C�_�7�(������x�F��Pi��|+W�      �%Mo�ӟ�e��ğ���Y�C-�|555eߵ�t���طo_,[�,���|��g������8Ə0�P�И�     �xv��.\��Y�bE<����%5w(�W_}5���Lq�� p�ظqc���D�̟??/^0R�P'N��ĢE�     �b(�������������&�Ŗ��wvvf�;�ew�O
�7m�eR[[?��OFRڌ�����_�pS�     P;w����G����?������dh �����X�t�)�� w���͛��>�2����S�NI�`Ŕ)S�ʕ+����>�;wn      �oiz�믿e�`��X�xq�p�C9��b���Y�|���{�nlذ!ʤ��1�{ѐ��ܡ<�|������       ����?ǅ�L��4�FB�)�D���� �����@���X�bۗ^z)ۄ�h�1cF9r$�rؽ{wtuu�6      �si�Q�|��ߏ�S�����L�<9�^�@�>|8�=O?�t ��� o��V���ٳcٲe�%�8�#]U��;�į~��       �����O��2I�m�;�	Iip����7ވ���sw��)�'ND�����mv��S��|�}����O~�Ǐ      �'Exe��ߪ��Y1�RSq�ȑ �o�޽q���hii	�+/�6n�e�dɒ�;wn�h�C�tww�����?�a      �/ip�C��L/^���#-� �C�������#p��_��gϞ=Q�����/��I�&E}}}ܺu+��x뭷�^p�     @���O�2I}�K/�0�ry����?�yL�:5 �;dRhw���(��k�:�ɘ�6d�O��<.\�}�Q���      �p�ҥ����L�{�9}�F���ŷ�~;~��_ p����m۶EY�i��?�|�X!p�rz�w�      9�q����닲H7��{�-QWW===���͛�'?�I�g�N�N��ڵ+�_�e��/d�;�NC9uvvFWW��      ����.�����_2������_(��7o���۳��N�N�	�e1mڴX�jU�X"n�r���-[��/~�      `lۺukܺu+ʢ��9�/_0ښ���P2�Ɣ��Q�T�L�N��9s&�=e���?�����;�W
�_~�娩�$     ���2L^z饨��
m�
(�.Dggg�������R{��w�,��������f�ԩY����@�\�~=����v     �1l߾}q���(��s��3�<0ܡ��z�-�;�'p��zzzb�ΝQiz��ŌE��2E�/^�|Ҵ�;     �صiӦ(�4��
�;������I����e%p��v�����Q)6���,m��PN����Ϙ1#      [._��Eve�hѢ�3gN�X1mڴlp`___ ����[�l�_��e%p���m�eaz;c]
[?��� �'mʶo�?���     ��%��[���R��/�0������ɓ�ʕ+��֭[�?�i�������R���#G�DL�2��vƼ��� �+:{���     Cz{{K5<pɒ%1k֬��f���w(�7n�|k֬	(#�;��N7���e���WWW�ei3�W�0�����x��      `lHQݵkע����W�X���ÇP>�������S:)l߱cG�A��h���c]ڌ��r���t�L�     0v���,���b�̙c���P^�p˹s�b���e#p�t8�/_�20����������Ҝ��lϞ=q��͘0aB      0����J31���*~���Uw(�m۶ů~�����S:;w�2H��;::�"m��P^w���"��{.      ]��ݲ���n3�555P^;v�_���R:wJe �+�u��yS#W�ǎ���{�=�;     �(Ka{������n�X6iҤ����[�nP>i`�}�b���e"p�T���[��޸q�bŊy�D<p����z�jL�2%      �;�˗/G̟??ZZZƺ4��̙3�Ӷm���RI�aˠ��#Ə�'w MٵkW���     ��غuk����?����Cy���i�{ccc@Y�)��7ofWu]�R�5k���H��}�;     �(���={�D<��1w�܀<�T@�����)(�;���Dooo]�>ˢ�<jhh�������	���?/^�3f      #k���q�Ν(��}�{y���@����{wJE�Ni�ڵ+�`ݺuy�nH��g�Pn����G     ��J�\L�<9�y晀�0�8q�D�?>fΜPwJ�֭[q���(�����Uڐ	��;     �Ȼ~�z)ڊd͚5QUU�ӦM����{�n �������/�PwJa�޽���E���|'��y��1��<y2.]��=     �������E����Ɗ+�$��S�LɾG�K�N��)�4	����룽�= ��@���{��_|1      )p/�e˖ń	�&5w(�O>�$N�:O>�d@�	�)�۷o������V�\�ƍ�3�;0 N�     �������2X�fM@�������۟��g�;� p����ۗE�E�����S�N�555EUUU)����ѣG�ڵk���      �4|(ݲ[tO=�T̚5+ �RS�k׮��/Ptw
��?�2x��c۶m����W��!#����c�ԩ���P?����w�      �>� ���v�,MpH���>}:�̙Pdw
-�q���Q===�	�����ĳ�>���Q[[�iC&p�;     ��z�j?~<�.��p�����+w�N�N�;v,�_�et����Y�~},]�4֮]���c]ڐ<x0 ���w��qP     `���i�`ѭ^�:�U�j	�s��� �-����Pdw
-M~-����/LuO�{[[�Mc����t3ɡC���Z      �4��*�J,^�8 �RSq�ԩ �����q�ܹ�={v@Q	�)��{��K�_y�l�{GGG<��1u�Ԁ�D���	�     �Ǎ7�ȑ#QtiB���ۿ��V���5 ����t���"�SX�/_����/����-[b�֭1o޼l�N*WUU�6�;0X
�����>      z��틾��(�������̞3f���˳^���> /��� I=ŏ�〢�SX����^:�|�ر�ihh�6o�W��ɓ'�����ĉ��>�����p�B477      Ck�޽QF/^�6��͛���-k%f͚0�8~�x\�v-�H�Na}����û~�z6�}۶m��SOźu�b��Q�TFZڐ	܁�=]�     0��޽[�����'v�ڕ=---�D�����������4�6����s����BJ/�]�zl`���i�b�ʕ�bŊl�6���!;y�d $����     ��9|�pܼy3���ٳٳ~��X�ti6pƌc�ԩS���:;���G	�),�;�t�ԩl"9�����ٕ\�6m��f'��͛g�;�Ήc`���h�5      ��{�_��ݝMt߽{w�H�VbѢE��bL����V^�x1 ������QS#�x�TSH酛���;;;�'������>`8܁�҇��V����      `h�۷/�j���q�ر�ihh��˗��իc����)5w I=ő#G��XP4w
����������T��k�ƓO>0������5�;     �иt�R�?>x8ׯ_�-[��֭[����֭�D�R	iMMM0��?�SHw
'M?z�h0�Ouoii�&�/[�,ƍ�L����q�Ν H</��r      ���p!���ӦM��+Wfτ	F����`�=������F�N�?~\;�Ξ=�=o��f���Ś5kb�̙�V:�N��'�����/      <�4��s���ذaClڴ).\�t#1#A�v���즑����"�S8�FGOOO�ڵ+{�������V҆L�Hq�ɓ'c���     �������s�����ٙ=3f̈�˗g�D}}}�p�������ի�D�N��ǆ����ׯ��K�ƺu벍<,2�~��     <�S�Nō7��w���l���͛���-�g͚0�Ə�&M����t3�����S(}}}q�ر`�����&��޽;�͛��R^�hQTWW|�;p?��      _��^===Y+�������hoo���ڀ����$p�j���E#p�PN�<�Ռ=�*�t� =�iGGG�Z�*�L�� w�~G���w�:$     �ҭ����g�f����c�ҥ�nݺ�1cF��HME� �+W�DWW�ފB�S()|c�K'H�l�[�n��T�ŋGUUU��tڸR�d�# �4��̙31w��      �����i+FIؘ&��޽���ĢE�w�[��Kؼ6P$w
%M'?Ouoll̮�Z�fM�א�f�<yr\�z5 ���;     ��s�ԩ,�f�n%b���z����qxX"V�~���{.�(���=��]��Mu߾}{vB9�TN'��o�+m���`Ǐ����     ��K�];�_���[�n��u��ł�|���� �{<E#p�0>��Ӹr�J�ow�ލ����I��+V�ʕ+c	A����ȑ#0 �      |;i�+c���ӦM�:��KL�81�A�N�555��� IWWW�O��(�;�az{�\�t)6l��6m��fS�[[[��p�p��/f�,�u�      <�Q06�]�|Y+�7JS��a�.��t�m͚5E p�0Lt-�t�t`�{
�;::�\}}}Plw�~�������      <�s���͛7�|�J�M�υ���ѣw
C�Na�8q"(�t���I�K�ƺu�b���A1	܁I��w     �Gcp`~��7o����X�zu̚5+(7Mp?�����BH�\O�>�G:���fOKKKvJyٲe1nܸ�8&M���>�u�V �     ��Do�����v�ʞ�V"����ʧ��) ;s�Lܾ}[CG!�)�K�.�F��Ξ=�=�ׯϦ��kVfΜC:q,f;u�T      �h�;���ĺu�bƌAy�����ݻYS1�����SB7���n'�H����իq�ڵhll      �Y�>�ܹsA���w�y��e�ĢE����:(��ST*������@���"�S�W�7pRyÆ�|��X�vmL�:5�Wj���Z�dI      ��N�<}}}Aq��9E��ihh�Z�U�VŔ)S�b����I�&����`�����@�N!���W�u�V�ر#v���rN�Bx�t�M�     �pR�Ny��y˖-�u�ֿ��/�����X�w�;0؉'�@�N!���7qR9��f�~��     �����ӦM��+WƊ+b�ĉA1��´f`�˗/Ǎ7� ����g�}�~�i��rR9_�N�555��� ��      �� R�aÆشiS,\�0k%Z[[�|kjj
���9s&-Z�gwr��ٳ����ʍ���I�իW;�<Ƥ�)r�x�b �p�B���9�     �zzz��V I��:;;�'M�����b���� �C���:uJ�N�	�ɽs��<�k׮e��7oޜ����[��^�T�ї6dw`���[� v֬Y     �WK��� 8�_WWW6�=�mmm�P@߿��x7�Pwr�w��ݻw�zR9]�bŊl���	��cC<HZ��     ����&i���]�����%
��������6y���ӝ;w`��~�@�N���p�t�RvR9Mv_�pa��kmmF��xk      �o&r�Q�!S�Y�~},]�4֭[3f�ƦJ��p��O`���糃/*�gwrO��p�����T��i[�jU6�}ܸq���b      ��R�����;��{��7o^6pѢEQ]]�-�������e�s��	�+�;�v�֭���OF�ŋ��c���[����W��Y�f�+m�ҩ����  p     �z�;V�+�#�;v,{b����`�)S�c������nw�L�N�]�p!`4���d'����Ғ�Tnoow��0����6�׮]���Q�@-�     �ˮ\����p���زeKlݺ��S�/^UUU��ijj
��H�	�ɵ��hK��ҳaÆ����6pN��t]N�s��<�A�a��!Zccc      �e�6����ӦM��+WƊ+b�ĉ��Ө ��"���	�%������cǎ��SOeWr-Z�(�����w�������ȑ#�f8� _%��      &pg�]�|9�iӦX�pa6���59i�{��:< `@�	��5��҆�����3iҤ�r��M�2%x����СC�k׮8z�hܽ{7 F
��ϟ      |�魌�������̞4Q���#k%����5nܸl(ا�~ ����Ν;Q[[�GwrM��Xw�ƍؼyslٲ%0�T�DUUUY���Ķm۲S� ��Z      ૝?>`���2MuO�D[[[�^�:f͚�t�@���ח5---y$p'�Dm�E�P~����<yr�\�2{�����7n�+W���e-      ���m�0Zzzz����3gΜl(�ҥK��F�6�nݺ�Mq�_Z��+�r+]m��!y�~n�~��x��wc�ٕ\���Q�T�Ҥ��^{-�= ��ҥK     ��������c��ӧ��7ވ���,v�6mZ��]�G��cǎe�N�S�WqЍ<��[W�^ͦbC^ݽ{7��ߟ=iӖ&��X�"&N�E��fq��۷`(�     ���M��
ƚ�7oƶm�b����0����UUU�WK��޽{㣏>�S�N��<������[i
4E�yްaClڴ)�,Y�Mu�;wnE�q��C�ٳ' �R�F�UWW      �3���,�����466fCӓ���ݸq#;�{������G!p'��䖉�Q
�Ӊ��477g'����c���W�������Z,����חE�/     �"Qyq�ڵl �ﾛMsO�D��^�T��zzzb˖-�s��lz;���y&p'�Lp������_�7�|3�����i�'ׯ_����������pIk�;     �	�ɛ4���?Ξ��_��bŊ�8qb�ɡC���^�}<�4D��ݻQ]]�7wr�w�"Mu���̞����r[[[�7.Ʋ������?����:     �e�g��wÆ�d��|Tw�܉�7Ǝ;`(��C���>}z@��ɭ�W���ٳg����}6ս��=�ݛ��c��y�f�����^k      �L�N
8s�̬�H�D]]]ɥK��׿�utuu�P��Wwr�ڵke�����^�����r����֎�?Z����o~�p�B ��tc      _dHEs���x�ײ��˖-�b�Y�fEޝ8q"����;nݺ Ć7�J�Nn	��4�==�ׯ��K��ڵkGu���o�G�	��bM      �E)�M�Ӡ�zzz���s�����������?��?q�Ν w�J�Nn��
_�>�صkW�<��Y�hѢ�����C���͛`$Y      |�����P��7FGGG�755E<x0���޽ �Ś����K)�}�v v�ԩ�ihh�+Vd�ɓ'���駟�+�����0�Lp     �"�Z)��7oƶm۲g��>�3g�������ہa'p'���I��pҟ�w�}7��>o޼,t_�xqTUU����?�1��`�Y      |QPe50���1V�\�=�Ǌ����Wܹs' ��իW�H�N.	��Ѥ��ǎ˞4�}���z��!��~�ȑ8p�@ ���.H�s�J%      p.$����M��w����+Ml��o~c� 0b�	�+�;�t�ƍ ���nٲ%��k��ٵ\i#�m�����lz;�hIuwwG}}}      `p 6x(�iӲ��+V���'��?��������0R$����͛7x<}}}q����ijj�U�Ve��'L��H��֭[�ҥK0���@�     p�i��`�/_�6d��.\�Mu�����СC�s�� Iih`j*F�P<�;��Z)P�7b�ƍ�������۷�h�6      ����^�����3{fΜ�loo����a��������o�)� #-Mq��7wr�w�7pӧO����,v������~tww�h�6      �\
ـ�s���x�ײ��mmm�z��5k֐�o����4�Q����7�;�dJ+�����^˵t��X�n]̞=���{���������A      ��ãK���ڵ+{ZZZ���i�{mm�c��.\�~M��b]@	��%��4���?̞�ܲe�b߾}���k     �����ٳg�g����P��k�Fss���^�������b]@	��%�at����x�k     �{��t#7��������w����X�jU,\�0���������ĉ0���:�\�}�v �'m� �k     �{Dl0������ѣ�3iҤ����b�)S�|�߷u�� m��GwrI� v�Ν      @���ƍ�e˖,^�7o^<�쳱x��/Mu?y�d�9s& F�g�}�7wrI� fm      p��FF��~�ر�6mZ�\�2V�X'N���m۶�X`�;y$p'�Dl �`�      ���`�]�|96l��6m�%K�Ă�СC08�F	�ɥ;w� � k     �{�������w���+��#�;�dJ+ 0��     �=�7 �6 ���R:� 0�w     �{Dl �`����\��� ��      ��� ����#�;�$b �6      ��ͷ �`w�H�N.�� ���      �� �Y�GwrI� fm      p�� ���7����R����\� �Y      �s���  ����UTWW���\J/�  �      ��� �������K��; 0�5Z      ����Y�7wrI� VUU      � �/�{�n@��ɥ�ِ �      ��) ��(L���% 0��     �=w �~&��7wrI� fm      p�	� ���#o�䒈 ��      ��J�  ��*��;�T]]  �      �� ��> o��RM�] �s���     �� �2��F%L.�7.  X      �S�T `0�;y#p'�Dl �`�      �TWW �`����\� �Y      �cB+ p?7��7wrI� V[[      ��
 |Q�ۭ��;�$p �6      ��`  `������;�TWW  �      �1 �ڀ<��K&L ��      ��� &p'��䒈 ��      � 0��y$p'���� `��     � 0��y$p'�� �`w     �{Dl �`���y#p'�&N�  ~     �g��� 0@SA	��%/� �`&�     ��{ `0k�H�N.544 @�����X�     $"6 `0��#%����  �u     ��� �`����\�4iRT*���� ���      �3� L�N	�ɥ���,r�~�z  ����      �SWW�u}}} ��y$p'�R�&p Lp     �\�R�&�޸q#  Lp'���V��Ξ= @���     �E���; �H	��-/� @bM      �E)p?w�\  H	�ɭ�S� ��i�     �� �. ��䖘 H�	      �H� $UUU1a����[&� �5     �544 @:�V�T�F�Nn��
 ���9i     p��ġ7�J�Nn��
 8�     �e�'O  k�J�NnM�81jkk�Ν; ���     �� ]y%p'�*�JL�>=Ν; @9��       _$f ���+�;�6c��; �XZ      �E&L�������	 ��z#���Zsss  �e-      �`ib�'�| @y	��+�;�fj+ ���      ��	� �;y%p'�Dm P^�J�Z      �+� ��RW1eʔ�<��k��� �Sڄ���      _6}��  �+u552a��O.���Ԕ� ��� P.��     |5C�ܬ�3�;�VUU���={6 �riii	      ̰  (7�;y&p'�R�&p��={v      �`3g� ��v#��䞸 ��w     ��6~��hhh��ׯ P>w�L�N�	����      �^
�� PNw�L�N��
 �3iҤl�      _m֬Yq�ر  ʥR�Dsss@^	�ɽ�"\SS��� ��n      �,� @�455E]]]@^	�ɽ���lCv�̙  �aΜ9     �כ={v  �c@�	�)�'�|R� %��O      _ϭ� PN� ���B0� �%n     ��555E]]]��� P&��ww
A� �QSS�f�
      �^�RɾW9y�d  �!p'��B���6e��� [�F+E�      |��	��<RK)p'�AB�Nkƌq�  �-l     ���Vv�� @9477gM%���;w�� J��'�      ��V �\��Ƽy����� ��Z[[     ����J���� ���"�Sb7 (�q���O<      <����GSSStuu P|w�@�Na�嚚���� ���ΝUUU     ��KS�� Pw�@�Na��=mȎ; @1��     �ѥ�b��� ��ɓ���1 ��ʼy�� P`�     �G�n� �逸�
(�;�"z�b�^     ���w,�J%��� (.]E!p�P�y�  ����9�L�      <�����5kV�;w. ��jmm(�;�2y��,~�p�B  Ų`��      ��I]� P\UUU��SO����I�� ��M-      �^
ܷm� @1���D]]]@�)��oݺ5 �b1�     ��kmm ����S$w
�tW (��S�FSSS      ����Ǐ����  �'��E!p�pR�6mڴ�|�r  ��      �㩪����~::;; (mE"p��-Z۶m �/^      <�����N�ӧO(
�;��d��; H:�     ��1� ��{<E#p��Ҕ�J���� �[KKKv�     ��3w��7n\ܾ}; ��H��@��)�I�&�O<�O�  ���,      <����hmm� P&�S4w
+Mq�@���t      �F��*p��hll����"�SXi��o� @~�)"��     :i�Ы�� @1���J�P$w
+�p�Ǐ����  �)�����      Cc޼yQ__�n�
  ��0`(�;��&���I|�A  ��lٲ      `�TUU�cϞ= �[�ܞ:I(�;���8�; ��     `�N� �����'O(�;���ޞ�P���  _fϞ���     ��Z�dI  �gz;E%p��b�ܹq�ĉ  ���v     �ᑆ555ťK� �/��(*�;���8�; ��     `���b6m� @>�7.�y晀"�Sx�ꫯ �'N����      ã��]� 9�x�⨭�("�;���O�̙3���� �C:�VUU      �����㣻�; ��I��@Q	�)�ɽ�� ��ʕ+     ��SSS�-�={� �/�JE�N�	�)��	� &L��}�
     ��Ja�� �gΜ91eʔ���S
s�΍����t�R  c[{{{61     ���4���? ��0���SQ
i3���7n `lK7�      0�&O���͋cǎ �+V�(2�;����
�`�?~|,Y�$      i��� �c���1gΜ�"�S����{WWW  cS� ���6      �����������;���?��a���c AD���QA0"���hS��[�&�$�MbV�ny$�dc��^+I���w<QO0FQ��>_�嚣g���z����-���3���TUU ��Ұ_h��䍂��2dH�q� 䦡C�      ��u�����_= �ܗ6�AC'p'�TTT� G�h�">�O�  n�IDAT��      �v�PN� ����,�t���	��+:t�N�:Ŋ+ �-餕���      �v80n��  r[ڔVPP��	��;C��@J�;      ��}��@=p衇��;y'�i��m� ��ڵ�8       �@nkݺ����!p'�EϞ=c��� ��Ç;B     �����o����  rOEE����!p'/��N� �!]|6,      �;i`��K�.  �2$ _��K�f͚���� �[�{��~`
     @�JS�� �{:u�;v�w�RqqqvQv�=� P���*      Խ�����Ɩ-[ ����o���	��n���f'�      P���n���O>�d  ���� ***����եK��ܹs,_�< ��1lذ(*�      W���w ��{������|�&"�~��q�u� P7F�      �C9$��g�x�� �{i���;y-�q�7Ć �]tPt��1      ����YO�hѢ  �Viii���? ���k%%%1lذ��{ �]GqD      �{�)�w �{C�����|#p'�5J� ��E�1`��       ��������J  ug����H�N��СCx���lٲ  jǈ#���GQ     �\UYY)p�:Թs������בG)p�ZRXX��@     ��5t�����~�ׯ ���5* _	��4(��w�x�w �Y�}�M�6     @�*..�aÆ�]w� @�jڴi2$ _	�!>�$�v;���� �f�3&      �}GqD�}��QUU @�I��JJJ���Oeee�v�m�q��  jF�.]�[�n     @�k߾}���#�,Y @�9������O�f͢��"���  j�رc     ��#Mq�@�I��:v�����	�G������Z P���bРA     @��~��~ϳf͚  j^�!�	��:t��rH<��� T���:*5j      ����1jԨ��� �Y�[���;�;��c�9F� լY�f1r��      ��9������o��7 Ps�<��ls�;�;��8 z��K�. �z��&M�      �OfTQQ��{o  5���$F���vh���w �&���ٱ�      �_GuT�w�}QUU @�>|x�������7:w�˗/ `�92Z�l      �_���ѻw�x�� �^1z�� >"p�Hocǎ�+��2 �=רQ�l�      �߸q�� P�ڵ�#w�C���n�-�z�  �̰aâM�6     @�׳g��֭[���� T�����ww����q�1��UW] ��K�G}t      �p�;6.��  �G�^��K�.�����СC���o7� �@����,     ��e���ѡC�x��7 �{���g	���ɳ&L����: �]gz;     @�TPP�Mq��/~ ���ܹs���3�O��NTTT�w�a�; �4����<      hxRKq�-�Ě5k �s�sL�y�4�;�D�@��D���  v�Q�F�{'      SQQQv����  �Lǎc���|��vA�y��?�!V�X �9rd�m�6      h��������w �C�&M2�>��vAz�<yr\r�% |����0aB      а�)��Ǐ����7 �:��_@�����ѽ{�x饗 رѣGGYYY      ��UVVƝw�i�; �c�=��v�w�S�N���� |VӦM�)      �S�`�u��1����n�ѣG���;/^ ���7.JKK     ��������U�V �s�'O6�vB����㏏^x!�m� �GZ�jGuT      �_���'�5�\ ��ҥK0 �/&p��ԩS�8��� �#S�N�ƍ      �gذa�hѢx��7 �|��0�vN�{�㎋�<6l� ��:w�     @~*,,�ɓ'�e�] �����#z����	�a�l�2Ǝ��rK @��>}���      yn���q��+�� �gM�6-�]#p�=4~������c͚5 �*���gϞ     @~K��L�?�� ���Wt��-�]#p�=T\\�w\\u�U ������b      >֫W��۷o<�� |�Q�F1u�� v���BEEE6�}�ҥ �f�رѮ]�      ��N8�X�xql۶- ��Q�FEyyy �N�{!�5s�̸袋\��W���b	      �Ծ}�9rd�{� ��Y�f1q�� v���R�Ν]��w�O�%%%      �h����裏Ƈ~ ��R�^ZZ���C58���'��>�  ��;��c���      ;ҢE�?~|�t�M ��m۶1jԨ v���A�a5eʔ��� �F���'�      �g�ر����ʕ+ ��	'�EE2]��s��TVV�C=/��R @Cu�QG�~��      �ER�7}����K �M�^������;T�4�v֬Y�����u�� ���u��1q��      �]�¾�}�Ƴ�> �/�&��N:)�='p�j�&ڎ3&-Z �Мx�QRR      ��fΜ/��Blٲ%  �����<�='p�j6iҤx�'bժU š����      ��ڵ�B�;�3 ��kٲes�1��;T�ƍgǋ\|�� AӦMcƌ      {b�ĉ��#�Ě5k ��W4i�$��#p�зoߨ����~8 ���>}z��>      {���$fϞmX  Z�>}bȐ!�=�;Ԑ�3g���?k׮ ��z��#F�      �iX`���㩧�
 hh���㤓N
�zܡ����f��/�� ��h�$����      ���¿_|16l� АL�81ڶm@��CJ;��?�x @}3u�T_      T�����4iR\�� EǎcܸqT�;԰�O>9�,Y��~ @}ѭ[�5jT      @u=zt<��#��k� �w1{��hԨQ �G�5�y��Y�~�e� �%%%1w���"      �Saaa�r�)���~7�l� P���[ݻw�z	ܡ4(F�<�@ @�;��]�v      5�S�Nq��Gǭ�� P_�n�:�L�@��C-�9sf,[�,�z� �\էO�9rd      @M�8qb<������ �71gΜ())	��	ܡ��7�y�������غuk @�i޼y�z��E      Ԥ���8�S������z���2z��@��C-�ҥK{�q��7 �Y�fE˖-      jC�Νcܸqq�w �eee1mڴ j��j��G�/��K� �#FĠA�      jӤI���矏W_}5  ���ٳ�iӦ��;Բt�ּy��_��_b��� u�]�v1cƌ      ��֨Q�8��S㢋.�M�6 �ѣGG߾}�Yw�鈒�����/ �KEEE1��hҤI      @]�СC����_�:  W����S�P��PG��� ԕ�ӧG�Ν      �ҨQ�b�����SO �����đ��� j����I'�˖-�իW ԶtdV�A!      �9s�ī����^ @.�4iRt��5��!p�:Դi�8����G?�Qlٲ% ����q�i�EAAA      @.hѢE6��?�iTUU �=z��G@��C�֭[�p�	��_�: �64j�(�`UZZ      �Kz��Gyd�u�] u�Y�f1w��(,,���!�5*^{�x�� jZ�Xս{�      �\t���ǒ%KbŊ u�K_�R�n�:��%p�q��'�o���� PS=��l�      䪢���7o^\t�E�y�� ����0 ��'p�Q\\g�yfvq�� T����3gN      @��رcL�:5~��� Զ�>4}�� ��rH:���N��/�8��� �K�&Mb���-      ��G��%K�ēO> P[JJJb�����Z�n�!����'&O�7�|s @u(((�SN9%�]      �E�=�ܹs�{��^��� ���O�:Pw&L����z��/	 �['N���      �7���:+.��ذaC @M:��#cذa�-�;䠴��SO����ov �W����{l      @}U^^�Mr���UUU 5�k׮1}�� ��rTځ�`����w�k2 {$����N�6N     @}6`��;vl,Z�( ��5k�,�8�(*��B.�9�}���$��.��d vKiii�}��Ѵi�      ��`�ԩ�bŊX�xq @uI��͛mڴ	 7�!�80�L�7�tS ��hԨQ̟??��      Eaaa�~�������z�� ��0mڴ�۷o �C����	����/ `gN<���ٳg      @C�N2NÞ~��Ė-[ ��СCcܸq��;�'�tR�\�2^|�� ��3~��8���      ��]�fC����� �=թS��3gN �G��D�F���3ό�}�{Y� �h���1u��      �����2^y�x�� vW�-b�Ѹq� r���t��W������k׮ �.M��;wn      �Y�f��o�K�,	 �Ui��g��[� 7	ܡ�iӦM�s�9��(6n� жm�콡��$       _�@q����}/V�\ �3ip�)��|p �K��P�.]�d�\rIl۶- �_�Ȭ/���-      ����8������~�_�> ��L�0!�@n�C=u�!�dGm�� �S�ƍc�Ѯ]�      �|վ}�8묳�'?�Ilٲ% `G�'O �	ܡ9rd�Y�&n���  �řg�ݺu      �wtP̜93��� �t��i���>�;�s�&M�M�6ŢE���PXX��zj���7      ��~����;��w� �]۶mc�Q\\@� p�`ڴi�aÆ���{��-�$�5kV2$      �O�2eJ���{��� 4o�<�=��hٲe ����;�|�ɱq��x����k���1r��       >+5�g��"��{. �_ib��g�����/wh �ک��[�n��{, hx�N�GuT       ��Q�F1����˗/ �Oaaa�~��ѭ[� ��;4 �My�ܹ�$�g�y& h8�=��8��      ع&M�Ĺ瞛E�+W� ����<@�$p����(�<����OK�,	 �ѣGǤI�      �u��O|��_����z��  ?��1bĈ �/�;4@���q�9�d���e���k���1cƌ       v_YYY�w�y�$���{/ h؎;�;vl �������,r�����믿 �?��9s�dGg      {�]�vG��֭ ���:*&L�@�'p��iӦ��/9~��śo� �)n?�3���0      ��ӱc�8���A��ׯ �#�<2N8� �;4p-Z��o|���$^}��  �2$N;�4q;      T�Ν;ǹ�?��c�ƍ@�p�a��̙3h8��5k��u���K/� ���ʘ5kV      P��u�.����g�y�� �~4hP�r�):h`��}۶mU4hM�6��|�+q饗���? �Q�Fŉ'��      jPϞ=�3Έ�.�,�n� �O}��y��Eaaa ���}[ ^III�s�9q�WēO> ����Ǵi�      �y�����O?=k(�S �Oڬt�YgEQQQ O��]����=�B���+��� �V�֞��q��      P{_�җ�k���#|p,\�0���h���>�AI�{څ�&�?���@�Hq��3b���      ԾaÆEӦM���/�-[� ��o߾�`�q;4pY�m�6�!��)���]���O
 jWz�3gN><      ��ӿ�8묳��?�yl޼9 �M��z���ـW�a����yh���&M��m�� Ԏt�5o޼��C      ��_�������cÆ@n:th̝;7(4|Y�y�f��@�<yr���č7�UUt �IiSQ�MܧO�       r�A�~���?�u�� ������O>9�
�,pߴi�������m۶q�W:n���l�2�9��ҥK       ��k׮Y�����$��� �n��m�ԩ�v�3Y�q�F5+��V�Z�%�\�"���k�.�=���      �]�;w�����o��o��� u#��ӦM �l��.p2ݺu�/�0.������� ��ںp��hѢE       ��}��q�d���U��ړ����1v�� �S�oذaK ��6m��7��l���e��=7x���;wn      P�~�k_�Z��\�2 �y)n�5kVTVV����}�ƍ&��RZZ�~�����~8 �}�G��3fd_      @����ƅ^�^zi,]�4 �9EEE��C=4�������� ��?0�m�6n��� `פ��ٳg�a�      @����w�yq��Wǣ�> T�f͚��G��=p� ;��O�4)Z�n�^{mlݺ5 �|�[,��:(      ��!��7o^���P�R�v��F� ��w�}wc |��ÇGYYY\q��nݺ �:v��&N'_       ��!����կ~eH @5�o����=��l�}����Q�F�yz����ַ��K/�7�x# ��~���i��M�6      ��9rd�j�*.���ظ�\Q�=շo�8�3�I�&�IE��|��Ѽy� �"i*�7��͸���'��|��4�7.�N���      �e�~��/�5k� ����2N>��(,,��q�~�z�;�KJJJb����hѢ������* �Q�A<w��0`@       �e����/�0~���������KA��3��#����q�nݺ �UiJ���㳋�+���k�w:v�,����       �S�V��.�+��"�y� ��A���~zr�!�E>�׮] �+����|'.���x�� TTTĬY��-      ���~o�p�¸���㮻�
 >+<묳�C��3w`�����׾����\�ZQQQL�6-ƌ       ��̙3��_���y�� �#i��y�Y�f�+>���� �S)��~�v���ƍ�!�w�}c�����      ��:4�N|饗��ի �ĸq�b�ԩ�}�]e�;P�҅Z�.]�+���˗@C0p��8�S�$      v�s���o}+.���X�dI 䣒��8��ScРA���@�+//�/�0n�ᆸ���* ����l�1c      `W�h�"�?���馛bѢE�	 ��~��3ό���/ ��ǁ�{� ե��(fΜ�rH\u�U6� �N:6��3�p�      ���6mZt��-���X�~} 4t�/}�KѴi� �S�k֬	��ֻw��������+��_�\WPP�F���?>��      �7�غ���cŊ��M=�w\�?> �ƺu�����m۶�E�:�j�*;v���������iӦ �E-[��9s�D�~�      ������7��͸��⡇
���u��1���ڵk �w�y���֭[c�ڵY�
P��D����8���i�z �A�ŬY��y��      P�7ns���n�򗿌?�0 껁f�KKK�:|*p�����I�ȭ/�0n���l��# �R�&Mb����&      ��6x��l������/� �QqqqL�:5ƌ �i͚5��� 5�Q�F1iҤ�ݻw\s�5��[o@]H�Ci���       ��u��q��m�ݖ���� �/Ґ��O?=:u� ��3�W�^ ��{����|'n�����`�;Pk�6m�|�92


      ��f8��l@�ڵk ����#���ӧg�j�g�U�V@mJt�M�C��.֖/_ 5�o߾1{��(++      ���~������q�u��_�� �E-[��9s�D�~��&���۟�W�\ u�s��q�f�n�y睱u�� �N͛7��3g�СC       ��h�",X�?�x\{�~�� ��ʆ	���@MK=���EEE1eʔ6lX��W��^x! �V:���";+�P       W<8�v�W_}u,Y�$ �R�&M�ޢ��2 júu벍~�
��y�زeK�ԕ���8�����믿>>��� ��ڵ��O>9z��       �A�֭�_�j�u�]q�M7ŦM������7��^VV �����n?U�WUUŪU��}��P����4ɽw��q�7d�{z���5���:*&O�l�      P�nb̘1ѿ���//��B Ԇf͚Ŵi�Lm��ʕ+�ۢ}A�䊖-[�ܹscĈ���&�x� �"iZ�̙3�C�      P��i�&�;Ｘ����w��]lذ! jJ�~�b֬YѪU� ������ً@.9蠃����v�}��q�-�ć~ �Զmۘ:uj<8       �4�=MR�ӧO\w�u���@uJCH�0�C=4 �R�ؓ����_ f�o6,n���,v���
 �5n�8ƍG}t      @C���ƹ�O?�t��W��5k���Hh***bƌQZZ um{Ǿ�	� �,}�J;��_}������Y�w\���      @>�ׯ_���#���+��ضm[ ����/f͚ݻw�\�>Ӭ\�2����=MDN�@.�֭[|���v&�������~;������O��"      �KM�6�x8�u�]+V��]Ѹq�8qb�;65j �⭷ފ-[�d�?�oڴ)V�^mڴ	�� �L�ӧO�+��[o�����0�k�.��>h� ��      �����}��ߎ�~8������������O�֭[@�ICڷ+����׿
܁z%�&3fLTTT�����{ol޼9���e˖q�1�Deee       I����rH60ܶm[ lW^^�������ԯo��B���_�v� �7͛7�3fdG��v�m���h�z���$F����M�4	       v���4X;���o~/��R �-u���0a���@�[�|����v������,fϞ�}@K��Q\UUU��*��eʔ)ѢE�       `����q��O<����cժU�t�CEEE��Ѳe� �Ҁ���@���י;wn�3&;��駟�C+..����?~|�j�*       �})n<xp���/��l8��h�z��ӧO�N�:@}�~��X�f���a�z������y������.�7�x#n��l���r�����{��      ���!ci�؈#�^�{�m۶��t��!��~�!�@}�����,��'�)�i'@C��~������}ѢE���ݡ	�      j^t:s��8�����o�'�|R/D�֭cҤIQQQ���P����>7pOO�U
��Ν��R���;��G��[�P;�4iÇϾ��       �#Mx^�`A����D���~:��)m\7n\�=:;��>K��?�s�W^y% ��;f���ɓ��c<���q�� jF˖-�� cƌ�f͚       ��k׮q��gǲe�⦛n��K�P?���ĨQ��c��4/����,p����IGqM�81����{�>�z�o�>ƎÆ����       ��x�����=���,tO�݁ܔb�#�8"�>�hC����ߏU�V}��-��}��X�fM���@�HG�L�4)&L��=�X,Z�(�x� �L��ݳi�����        ����+[)t���G�"l��ޞ|��� �&M�N���J�q�u�]��%�m��K�?�zh�7.��o�       �~��?��q�m��08jGiii�=:,شi� h�v������@�K�q���[o�����ğ���X�~} �ֶmۨ���#Fd�!       P?���7[i(��w��<�LTUUP�Z�l�~xu�Q�v /��w >R^^3f̈iӦ�SO=��w_v4䳂���ٳg�80
      ��a�P�+V����x�Gb۶mT�4X��#������� ��s�k����ǿ0pOaӦMѸq� �#EEE��i-_�<���裏Ɔ�ž��Mj9rd�j�*       h�:u�s�΍I�&e������ظqc {�G�ٴ����g���믿�����-[�dS��dV >�s��1{��9sf<����T�^x��\4HisG��6lXv�i�       ��M�6q�I'�ԩS��?��O�z�� v��#��ݺu�|�dɒ>���{�t�R�;�N�c��Ou_�jU�S9-q4]�v��Çǐ!C�Y�f      @~kҤI�3&F��<�L�u�]�����Ś6m�vX�7.��� ߥN}Gv�^������H��^{�x衇����k���[��C=4F����       ���� ��뗭7�|3���l��ƍ��.]�DeeeTTTD�ƍ�����x饗v����Jl޼9�N��IN�:���_�b�'�|26l��kZ�j��N"�޽{��       �:t��3gƔ)S��G�{�'V�X���IC��#�8":w� |�o��֭���v���=E�tP �g
�W�^�J���X��<�z�����J:�o߾�n�t���      ��JQo�T�ֲe�����'�x�Tw�F�n�b���1t��())	 v,�<;ܓb
��G:c��\۶m��_~9��{�X�vm@Mkݺu���ߤv       jԁ��Y�f��O?��w_���QUUА���ƠA�bԨQѩS� `�}�����.�/Ύ��z�i��/�N8�X�|yvA��3��k��Pҿ�t��!��m����E�       Ԛ40aK뭷ފ?�������;�P_e-�a��ݦ>�]�y��X�t��~}���_=֭[��2�f��]�t�֤I�����B���#��:���ݻw���o߾��      �	���q�q�e+�{衇��G���? ץ��ݺu�6kTTTD�������/~a�K���m۲�aҋ2 ��m۶1z��l���?�����q�x�.>i����={F�^�⠃�F�       �� �O��/�Gy$�aÆ�\����]�Ɛ!C��C�}��' �;�>��~}��$E�w�����J�rZ�ڵk?��S��r�� �l�{��E�)h/))	       �o� �tByZi`j"R���O��N�HQ������L��۵k T��{���ˁ{*�Ӵ���@�jٲe��9�$�K�.�b��^zɄ�h{�޽{�8����͚5       hH��~��e��O�_|1�x�,xO}Ԕ��"8p`�Lj�i��Ά��r�f͚X�bE��[R�N��~�F:��W^ɂ����}ݺuA��.��1li7p
�S�޸q�       �|QTT}���V�׿�5�y�xꩧ��_6���VZZ={��xS�a� 5/]ߙ]ܓ��@����4i�M�N+It��߲�=�˗/�6-����6(��״R�~�DYYY        ױc�l�?>�}�ݬgK�\�����LAAA6l�w��YО�� �����sv+pOǼs�1@��>�w��![Ç�K���o����)zO���Z�z��5$�,o׮]v�ݩS���vGZ      ��iժUTVVfk۶mY���/���?K�.�-[�$i�`�=�A�)j�i ԝ͛7ǒ%Kv���
�_}��X�vm��@����[�5x���ߴiS����J�{���B��қ;���j۶m��v�Ƃ��?       P}���Ӊ�i����D�ϥ��˖-������6?t�AY�~��Gyyy ���sjwf��4�7�}�/ O�ƍ?��������J��ʕ+���;�|��{ｼ�,..�����w�}��6m�|����͛       P7�4i�M�N+I��K/��MvOa]
��k8R�ѽ{�����n ���{�]z�n��O<!p�Ci�{���J�(��)rO���5k�����V:�#���׭[~�a��ߗ&��h��㕎�J�z:�$�O;|SԞ�       �)x�ӧO���8��S��&����kٟ��?r[IIIt��)�x��f����xꩧv�y��/^�8�KKK �K�}m�w&]��}����Ziwt:~d�ƍ�u���9�o?i��?)MUOk��7m�4������4�>�O�����o_�b       h�R�бc�lUVVf�}��Y�|��W:�^�^wRϱ���G�Ν���o�>kB ����U�v鹻�����'��#F ���޽YU����c} �����$jlJM|%F�ֶ��M��δ��&M�S'�tҙ���bZQ�5���@�"��G��օ]XvY��.��۞�BMb"�}�{��3�s��=砻�}��ږ�       �PK>���[��\.�x�hjj����ؾ}{zL>Ş��,,L�����~�A��z�@�X�r����������         �����'N��Λ%�ޓ�}ǎ���;w�L��'[i�O�筍;6N?��ÓD�g�}v�v�i�V} J[]]�������ק�B;餓         �E����.H��
�Bttt��{[[[�޽��$�'�8p JQ��|�����$dOfܸq�ׇ���Ç �)�4��MaG��|>�V�W]uU         @����8w�&]]]��ٙ.�ݳgOz<�8�������><�\.�BUUU�=���5*��IB�d���'3lذ ���r�ʣz�1��˗�        �UWW�3~��#z}��P���חｽ��$��e��^��%�9�~��d���M�#G�L��$^O��#F��O��m���t�G������]c��rJ          �+�
h�: ����hii9�s�9pO��UWW�\sM           ��-[���9��=����          �f�B�+V�y��oڴ)v���ƍ           H�_�>:::����
ܓ�>��~���           $�.]zL�W��X�xq|������           ���߿?V�\yL�w����7n�.�            (o���ӹ��'�-�w           �,Yr���K�����ԧ>���          @yjll�m۶��������k�?���           �i����u~��E�	�          �TOOO����u�~ܷo�1a           ��$q{.�;�k�[��H���          �Oғ�~ܓ���o�ѣG           ��7ވ����N��i�~��W           �?��'�5pO���+q�UWEEEE           P�zzz����_���{SSS�[�.���           �m�������/����=1o�<�;          @����`��~�ހ�?���c۶mq��           �iŊ�k׮~�ހ�_|1n���           �4͟?�_�7`�����S�L��c�           ����>^��~���}}}��K/�'?��           ��̛7�߯9`�{b��O|"F�           �����X�zu�_w@�\.K�,�뮻.           (s�΍B������=��/Ƶ�^Æ           ��޽{���v@�=��{{{{�X�">��           �m�����; ���=��/�����FEEE           P����.��J���Ԕnq����          ����/FWW׀]P��̙3��.����           ��twwǂ������Ĳe�b���          @q�;wn��A����/�<����           �}���K/�4���Ҽ��-�.]��G          ����s�E.����*�9s���ɓmq          ({��W^yeP�5���ݻc���q�5�           ٖlo?p����kH֨?��q�W�	'�           dS��|ѢE�v�!	������          �lJ��<xp��7$�{��矏�|�#1r��            [v��?��O��C��ݻ7�ܧL�           dˏ~������{Y���7o^\q�q�g           ٰaÆ�����i�~��������o�=           z�|>�z�!����_�n]L�4)           Z�-����!����������          ����3g��3�777��ŋ㪫�
           ���ٳc߾}Cv�L�g�y&>��Fuuu           0�v��/����2�wuuų�>7�|s           0����+�����ߐ��=�`�����?g�uV           08֬Y��P�T�����G?�Q����m           0�����,�T��H��������K          ��5w��رcGdA����?^xa�=:           ���1gΜȊL�QSS����          ��W(������ȊL�ŋ��_]tQ           п�f{����%��������c���          @���쌚��Ț����֘={v�t�M          @�x��ǣ��;�&Ӂ{b�ܹq�e����           �U�VE]]]dQ��|>������O�Æ           �M.���{,�*�{���)�ϟ�_}           pl�~����般*��=1k֬��K�3�           �N}}},^�8��h��������aÆ           G���'}��(
�eE�'�瞋o�1           82�=�X���F�U���3gNL�4)&N�           �v+V�����(E��������_��c�ȑ          �[koo�3fD�(��=�k׮x�'��[o           ~]�PH��wwwG�(��=�t��x�{��Ї          �_6gΜ����bR��{�����'Ʃ��           �-[��g��bSԁ����ӕ�������          P�zzzb������Ŧ��ĦM���矏?��?          �r��ODKKK����gώ/�0&N�           ���W_������bU�{�:ڴiq�=�Ę1c          ���ر#f̘Ŭ$�Dggg<����/|!��J�?          �m�r�tixr,f%U�o޼9jjj�[n	          �rP(�?�Al߾=�]I�����y��'O          �R��s�E]]]����3f̈��>;�=��           (U�֭�Y�fE�(�����7���o�=�����          Pj����{��^���(%�'��~����������          �R�,��w����RR��{bժU1gΜ���          �T<���e˖(5%�'fϞ�x�;��/          �b�p��X�dI�����B|��ߍ��+�=��           (V6l���z*JU��\.=�P��?�c�;6           �MsssL�6-<��,�DGGG<���q��wǨQ�          �X�ٳ'�N����Q��&pO$�X��w�w�ygTVV          @�����q��ݻ�ԕU��X�vm̘1#����<           �,������c۶mQ�.pO,Y�$�<�̸�           ��|�����~�,�ď��3fL����^           d�/�/��r�����B<��q�i��ĉ           +V�\�.�.7e�'z{{�[��V�}��q�g          �Pۼys|���O�z���������/��t�;          �Pijj��z(]�]��>pO������ߟF�cƌ	          �����<�@twwG�����;wƽ�ޛF�'�|r           �C=sggg�3���z��������          �������tttD��������:uj|�󟏑#G          �@ٻwo��{׮]���-���������>��1bD           �����4n߾}{���`���1mڴ��;����&          ���r�4n߶m[���ۿ�������������          p�8���7���1�e��QWWӧO������aÆ          �����I�������	܏�����_�������Ç          ����S�FCCC���Gh�������w�#G�          �#�w��x��b۶m�o&p?
�� �w�}�w�wQ]]           o���3퐛����N�~������}�sq�'          �o��֖�ǭ�������[��׿�����?cƌ	          �_��Ғnnooo����m߾=����������i��           �$�q�����#8r��k׮��7��F�g�qF           lٲ%x�����
����8�޽;��~�w���          @�Z�vm<��Ñ�傣'p�����&��n�->��          P~�,Y�=�X����F��Ozzzbڴiq�-�ĵ�^          @y(
1gΜ�5kVp|��(�����عsg�|��QQQ          @�:x�`���G,[�,8~�0��hkk��n�-N8�           JOWWW|��ߎ�7�C�>@^{���7�w�qG�|��          ��]�v�ԩScǎA��������W�w�yg�?>          �������ַb�޽A����_��W�����.          �x�X�"y�������}tww�}��S�L�n�!          ��R(b�ܹ���8}����|>555�������cĈ          d_WWWL�>=֮],�� [�lY477�����~z           ٵm۶�6mZ�ڵ+x�!�lq�������[�K.	           {jkkcƌq���`p܇H.�K��q����M7�          �|>�<�L�������B���ҿ��q�m���ѣ          :��|'��'pπ5k�Ŀ������g�}v           �o�ƍ���Gggg04����_��W��o�+��2          �������矏Y�f��:����3f�ڵk�3��LTWW          0pv���<�H���CO��Auuu�y����g?_|q           �o�ʕ�ꮮ� ����=�P|���O~�QU�G          �!����O?�-
�E5�a�B!�ϟ�֭��n�-�9�           �]cccL�>=Z[[��������򗿜nr���k���"          �#���c޼y��$����l�����x��'c͚5���~6N9�           �^[[[<��#�q�� ��Ef�ڵ����q�M7ŕW^          �[+
�x��x��#���'p/B]]]1cƌx�������bܸq          �����x��G���>(�"�f͚����������xTVV          �����x��c�̙q�����܋܁���&~����g>�?~|          @9jhhH��777�I�^"6o�_�җ�뮋?��?��*?Z          �C�4z���1o޼���A�RA����^x�X�zu��}	          �l͚5���G[[[P��%(�H��~��q��W��ܫ��          JI{{{<��ӱ|��t�KT�P��_~9�-[���Ǣ�ʏ         �����,�9s�DOOOPZ�%���;jjjbɒ%q�-���_          P�V�Z?�����-(M�2���S�N�I�&ŧ>��?~|          @1غuk<��S�q�Ơ�	��̺u��K_�R\s�5����1jԨ          �,ڷo_<����K/E>�J����������c�ҥq�7��{eee          @$���'?�I�r��|��XWWW<���ӟ�4�L�_|q          �P)
�lٲ�5kV�ܹ3(?wb۶m1u�Ԙ0aB|�������          �%	�W�^�nlojj
ʗ������fL�81��O�4.���          ���nݺ�����[���5�7o�{�7���wŔ)S���~w          @J��g�y&��mڴ)����ǤI�⦛n���??          �x$˘�����>�W	�y[ɻc֯_�^zi���Q�s�9          Gc�ƍ1k֬ذaC�o"p�
�X�re:�z׻�n����}QQQ          �V�u�����s�ECCC���s�6mڔN����k��ɓ'����          ===�lٲ�7o^���)�;Ǭ��)f̘3gΌ���:>�я��ѣ         ��w��X�pa,X� ������������f�J�a��8���7n\          PZ[[��_�W^y%z{{����~���b������/�<����x�;�          ��B��ׯO��5k֤_�����������6��������率�O<��          ���ٳ'�.]�nkߵkW@�3��o�5551s����>W^ye\t�EQQQ          �C��-Z���Z����Aq���X�bE:g�yf����+���N:)          Ȧ��������F[[[�@�3�ZZZlu         Ȩ|>6lH����ե_�`�3d޼�}�رq�e��?���0a��         `
�hhhH��W_}5:;;����Lhoo����3nܸ���K��}�ĉ         @���Ew2g��݇c�SO=5.���;         @?ٲeK��֦a{GGG@��ɴ���ñ�Yg����Ɍ?>          x{ɦ����X�|y����d������ܜάY�����y�{bҤI����7F�          �BWWW�_�>֭[�W�����!p�(%��-Z�NeeeL�0!�����E]�w^TTT         @�H��oݺ�pԾaÆ����F�N�K��nڴ)���'��nwO���8jԨ          (5���KC�$h_�jU�ٳ'��	�)9����t��t�����|g\p���w�;��>bĈ          (6]]]�q�ƨ��O�۶mK7�C)�S�<��O&1lذx�;ޑ��'NL���N:)          ����-bӦMiԾ}�vA;%O�NY���͛7�s�駟�nvOb�d�9�t�;         �`��r�u��4hO���_���΀r����ܹ3��������������8�����Ϗ��ǧ����         �xuww��طlْN���� p�_��磹�9��K�~~̘1i�~�Yg>&��G�          �*	ٓ%�I��t����v�
�	��utt��nݺ��UTT���g���駟�N����N��#G         P�:;;�`=	ٓimm=|ܷo_ GG��!�(����t6l��k�5jT�;6N=���8nܸ�x�'�)��'�tR:Æ          ;8�����ݻ7=&�r������w���� �ϡ�����_VQ���QOOO�ر#�ߦ��:�ޓc��}��ч'��G��F���UUUq�	'�����Ǉ$߷1        �r�,������璖/���������/r�\�'����$�O���+ړ��4;��笇.���{�ox�{��}����* (&�w�u��        8F_��ϫ���@Q�,�l�뮻FE�*            �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��          �L�          �	w           2A�          @&�          ��;           � p           �           d��       �v�X    `���4vG   � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �  Ԯ�6 �h ���T���,Sĕu�@�'pg���8        �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��~�y�_˲� �<ϗ       ��^��x <�i�~O��~Ǿ��[>         /c۶�[> ���           $��k����    IEND�B`�PK
     �9s[��n  n  /   images/6b551873-9f16-48c5-b1b9-2fc6ab10f815.png�PNG

   IHDR   d   �   +n/�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��io[U��Wl'q�fh�6miZ(P(C�2�|x��
�*\^!U�B|������ $�2�I@�g(3�<�i�$�<��ݿm/�4��Nb;��U�:�9�׸�^۷v�Z	����as�J|*0���o��Y�FNt
��[�1m_��?(}Q>P y�2�I�2��d��0��a�$�(H�Q��< Fy@2��d��0��a�$����SOɓO>)Ӧ�1���/((���By�g�D���!x������<�hKKK�u����TWWK �/�A�_��|�/F#�x�
JKK�D�U�V�=z���s���/���<���E�Ge}��O���.�����r�9�șg�)ӧO�_�F��2�O�W��ϟ�ɕ��Ef@���� '������o�m۶�P�%<���򴵵Y ���3g��2(�P]��G���zc�� ����<>묳���[��w�{�C���t�M�b�
��@;O�!� GU=����7�xþf��E]$w�u��D�y��C��}��7KGG�lذA|xW��8��8r�<��#5��z����_����eƌqՔ�� :88h?��,..��<����ò<`䫗
�U܈�***�ꫯ����� ���#�������r��!�wsB<1<�e˖Y`���O(�Q#�{�n��?d������ky?/^,K�,��<s#@����R,@ ��_��_]�9b_}e:�mٲE>��+v�^{�}�D�xs��ak�qaǒqi�o������n��.���%ڀ�u�A��5��������k�9��ڱc������}�Q�n�:9x�\��8�r����s�=g�ǢE��s���)���q�mmm%��}��ɽ�������NXTT$?������L��>Y�`���w#F�����+	ut��y��g���ώ�/�Ђ�:��h6���>��o=Z7�D����nG<����=�!?L�%}��6�d��ZL�qګ��j���[��K/����!��������vl�駟�7Q�~����|�r����~���	I���g>��SH���x��N;�4��#�@%�p�裏�w��~�Ao
�{@
���ᤵ��V7�L����%����#�i�&�=JJJ����'*͍0�dxq�4���@PI���f����I֯_oG<��t�RkS���c^4�sҪ���u�jµ�`��/�l@E�}��V:b����Μ93> �'F���h�y<b�J�g#�l��Ih
��~+555�����7�6�-k	����u��D�H4¦&��� �JB��ro�n3�%�C��`?�s�o"��ƛ��pR� ����ܹs�n�AG{�z�68�(()�� �� ��_|1a��#%�\�*� �u�1�\`A��W�w�6���'�������/�8���� F�HU�@�͛'W]u���/�]����\S'|�y�g�ډj���ґ�(#��P1�P)�}T���'Su�o�ݺ��[���<`y4��	�0��裏�+��"�y_7"2_�j�̚5+)ҡ �t�v��dp8t^�kU�G�hpL��<���L��c�=&/���͆�#�{T�Xj<f�#�?��CV��k�ڵ블	7���f`w��ɂSQ90~�޽6�RCc#��jj�#Xm���=��q4��xnj#⻤����P�H�XUI��95̡ǳ�q+u4�{�6e���q��o�H�����Ǎm޼�zy���n���M��&���ß�)�g϶G�~s���d2��kll��L��ʄ/'�tR��Od�&\J�?� 8/�c2�����n�߄Yc��t:�q�Pka�atõ��7��T�s�ZhH���x�sq�\+��)��r�{\�x4Ƹk{�m a8*f�ƍ�@j�NrdN�<���eV���5Sf�AQkF^yY��N�F���_::�䰑��C����Ez��#��B�0#Q�ؙ�J�+L�2���E#����Q�,np��`�a���e�YK�43�j���Q������2��2��a^
T�6��J�4̑�b����a���l���wȠyn%J�͇�3~��6͚�L�I�(3��O?ّ�TM#L#�/�@�_|�̬��ζViڹU6:(�248��Q���{
�WX$e�RS7S�<�t�	�ɮ��rd`� � �R���[���Λ�)��7Jf�:$5�j��������/)/.��[7��쐞��F�cm�S��Q� ��~T:����l_(�J�>���A9�;$�<��ະae
 *ݩ���`|��W֋rf����"�,�V"��e���d���� �����{b�|pN{d�%2��H�t�38q a���V���⊈�.J �����TQH��r�,�.�B�G�6J��	�`T'���3�,/�ș�e��{P{�1��T3�H��S}�F�/��b� c4�߂�2i�*������_Zp4@C�_J|���/((OXRv��i#~���	"�Ci��۳g�5�c��)5e2Ϩ��y5*-�J��k������V�l$L�QA�r@{�׿��kk #	?É��K�'a�f��k)���Ԑ�*	��Rm�S7�\<�AUU��܊i�V�`(q]uFR��h��5�H
e�����ȓ�kQ0 �ʸ���L,5���I�p@Z��#���@�I��J H�C�y)��3#nQm�}�fn�/��{( ��p^��r$$u�A*(e�  �z���o��3��@����{^E����鳪�()q+M�����cS�"�>�̭,�h�P
��|s߰t�=AJ�:<��#�}�)%� �='f��C�7#/��@�Po�I�P([���$e���$%�0��t� =�bVyqVH��y��'e&��ZՅ=dS�P�MI�Y��Ө-��ߨ�l"X�nTW����s�X�46�0�V[)��w��|��7����H��_u�O��Bb�O�d������P�2��}�4��h�I�%��*1*�g$h]`@���E2)%6�Y��+/�I��@�K����t��H�V�$���ǩ��d�9<fl$;�VJ<�{�'����${�$��p�\$ӡ�쇉?
�Y
E�Bj�+#��v��{c�j��2ɤ�K�h-ģ��l&��A5B���2��:�P,����<����hVˈ���pd��{LE�$��۲�l�e��6��7�#���&��$���H�>���[2�QH*԰�������@ h�

}٫�
B�;��үS��kcG�gP�;lt��X��
̠
�0ނ!  #�Z�.!�w8���%������did��S�:l���= F��TBXA�n�5����������30hT�h�����(���2�c��r���=��/���2�B� �%T�3�2>�9׏P}���/��[����0e���c۱:d�ɤ�KEJ�]Qe]Ds}C#���'��*�M�.Hl��!i�鋬[�5�1+�� BA˸��eDy�>���!��+%��&�utK�qL�U��V�H�SQ4���2�|;�������]�i���,��=-!�HS������J$�h��ֶV9`�dѬ�22��6H����FB���*��XYU� =
�c*4Q:+v78,3��O��փGl�)��d؏TUç�r�~��!�k���=��"�����9u6��d"_u��K��f �,{H��[��dPJ�(�� &aޠ���o{�dn�4)-.��
�Y��Ws�d|���6�r�HJ��ѷt1`1����
i;�.w7ʕ�J���Ǿ&i��^``?h�Ò��p�x$g�q�]9 ���<�*3*�dɼY��|��E���;o�� ׍!�+C�WR�|}��H	�-R�4m��(�b�o�|���d�v��w���VK(�`���A)Dq,��=9��Lp���|�u�\m���)0:���-�lv��o�����0J�C��nA,��(~`xX>۴S�0�d���)5�j�/��ξ�H��8�A�tu�N�*\n7�!Z�
�����7�e'ϓ�s�lf%]ޗ��3�^�o�97�/'���Ő��y@Zpc,1V#���������+�Ε2��.M%,0~hĸ�����f;l!����%�\bU�xvJ��1mt��� �
3o��P�4wt��sda]�-
��J���1��O�V��0�ל.J{��A�#Q[�π�=0h��n���"g̝)sk�I����:�x���oj�-�Hc[�Mr��$H-�ߍ7�hw����@S�Hk��O�%�۠kK�FCk��������D̨��T��m�����F����#�����t��fm[���Æ["��_$��Q�>�[lLi�,n���l��Ma�.��X�f0�����(] �+ʤ��T*K�RRTh��Z'��a�g$�hO���xN8����x"�PQl9���=���N���ʋ�ԛ�h#)���lS��vx`�g[�zCK���C�CxG�0@�ZC"F�Փ�v�M�z}�c-c��'���������Pg�Ήxg	���H}�Z(4�pɄN�ŝ~�u�u�YF
�x�W�Ą��Q58 �1��nq���g+8H�o�ħ��I��������9���DS.q�޹tc���/m_D�Fps������W^iG��<�E��k��L#}�9YhI�E�m�H[h0f�Z��m�)=�^��d	o��}j��U�!�(���&��`L@`8K��>�7C� �Z0�xK�n�ak�׉�2
�#�d#F+��1H+��Vm�1p`�Y
���&� ��-a����=2o����ZF��O�g�F��Uu�7Dʈ����J���6c��p� I���РF��n2�;+��E�u���
��DM(s��%��*����o�۳U�4J��1jv얂��޲�wi5�!ZL@�L0�w�y�e
���F{��=�$������.���s�F�����B���-�!�n�Arcm)F@ ��5����21ʈ(I9Fs*����v�`����R��ڦ�-qZܺ
E�T�Am���]�=����v�A5 &�-�@訊M��@�F�RC���嶥`�]�Hc`� l���q�}N�H��%�梨 y����d��5G����s�v�7��q�]�
ށn���xQ��-���X'�8!���d&ݤˡu�F\\T���`g�`�"���m�Ǩ*�7��0��܉�Ts�TB�d�(6�$��r�U	IB�%�m�G��������%�7�R��%7U�.�x���7ri�6�|9l?ՐO��3n��� D��b 0Q"e��sIm�ц7ZH>b�>a@���B6Q@k���b̝I�k≐��O2���S;�m���?�1��⫉n)HP�vn�k�/�X�º�L%J�i���p�	�'��۫1I"D��ʕ+cnH�3��f�5u��#��X�tH,�o I6ܹ\2�c�{�~W�^-�֭�Y�x�d i'7�<�8ad�1[{���(� �(��G�D�p$�	$#��P�_�B�ސ!Fs���e�5�{2F#���c3.MiG#��a���q��y��)��6#iJ��	��0��&��0��i�h�g.}�z��bef�=�R��^�6�D&����Lx��0���A�|$ ��z������]ɗM4�I0-a��^���K/ى�B.{H�D�ԟ�4�}�v�iY�p��b+��P^�KZ����y���T�x46�L�9�ׯ��)�ݱ[�:~�Ɉ�_���m���d;��}�����=�*��۶m�h^f!��[���r���������:��ۺ�/��w�o��<���:;;�� �f�V�}�RM��K�����gÆ?c�!�K�e�He�s3y72�an@wL>�)\��͹!&������ O?���/d͚5r��ڵk��q�NJ����[�韔$�(H�Q��< Fy@2��d��0��a�$�(H�Q�#' �M��S��iR|q�g���c<*I�s'1I��;��w\e���7㳑Y��    IEND�B`�PK
     �9s[9&��ސ ސ /   images/b01488b3-8551-4b4c-b09f-2812c4acc168.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  ��IDATx��y�m�Y��=�s����n�$�I��� �1���0(. U�D�	W���T��
�+�JR�#�B�Bʩr*�+�	6�6�hh���o���{�=��o\{�s�{��H�}��^����a���^��}���p8��N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p�������8�;�ñpBw8�c���p8��	��p8�=����p8{ 't���p8� N����p��h=��?���0>"�����0<�޿T�fS���bߔC�S��)�P��� ����e�C����0x`(gu��]� �(�X�_��y�����<�����:�=B�6�n���7�k���S�#�F�����S�1-0��!$�n<���!��`(���x~��'�����'�G�iX�s�q�8����:��q)v$7���GY4��1@�a�נ��?`�3��`�G1���3�����|��(��P�����ʢ⯥�(e#�]����eXq���8�W��&��n��g�^6���"t�����fq}�4��/������;�M8ٟ�瞀����O�(��p�$���yL��&�PA���-BꊠDO
����La(Z��g<�0Ȝ������I}"ţM-�I���\�C��x1D<���ؾ�,�"���U��_����>��W�7O��'��W�c7��－�y�������� R����g�H�7B$֌���fd�I���*��@�7%t2�}��|�W&��:	"!j�X�c$~���(�#l�bn:n��kuh�$���y,g~Y�����?o��oCc�F���YBY���c��pp��5�[Bo�^��|�vs'Oު7�/��>������?�R�UH�oA*|��Ȉ��;��0G��HDM��3	'}T�v:�lRO /o�g���q"�ٕ7���Zk��'�]�z�����>�=u�*Y���(��TAQ�ş�Y��+�>9����x��py�W���~z�Əݽ����!v_��Ư��T�8��:�e�����P��'mQfDr�^��L�l��0�Kll@��,�&���Mu�1$��َ'R��ь��ND[&�k_�Ch���{=m
��a�X>���D�.�-*Mź(ʋ0;x�<{aYՇЬϡ]�C}p"���w��.^䟛faqt\��_X޹���߆��N4���؟�l��)�u����	=z���S�(�a��<�ؓ	�I=�p{�|�\�b����d�X�]#y_¦_�r��
ϵCR�c�z��MQ�]�i�Ԋ�ҡ��B�d���U������>��!��������~���~i�6_��)��;��.�K��O"W�����ߌ���)��}w#v-���]�$oB!�3� �g]�0���zg�"Z�� +*�&�_
���D�7E,���dGeO>�<{�˘�b@��|�Z�->�	���2���3h��iQ�!��$��ֳ�����_����� ycI�8�u�X�7�N���g?K����N��=��au��hѾ?��si�n�^X��"7�B�L�=��T�t�2�ĉt�
�&�υ�)�moz�G�'���}�B�Y�MS��-��;G}	�8�[\�C? Q� ��hU�P��]ࢤ+ ����:̠�j<���&4q��0o�;��{����W~����?����O���_���p�Ʊ�l�B^-�����G��}ٛ�z�����}�M���[#-���S�dN2eM��@Y��q�o�U��	�D�!LB�&����׳+s*/�GCf"/���*���ҔD/(8�4�ʲck�,��>��~����
��?E�����^���������_trl/��ާ�Y��)Q�=�������8��Cw���+=� ;&Q
��ԍy��.T7�2�q͚�LD��1�<yF7�����~6�ϳw�>Ç�cH����Bo���*{�$�t}M۲�>�WpPԜ�W��y��Zz���",XC���� �1�z��_~���������o|ӗ���_ï�*@�� ���|�����c��ɧ��}�bx��x�[/����E���4ϴ�͢�܁�d>��B���OT��s�|������T{yޡ�� I=Q��š8LeQd<��s��)M��v`�<���Y��c��kfܐ�-J1�3=Z&(�Bq���1��W���Q��A�gB���a�������������z�w�m�\܆fyN�z���n	}u�.�G7`}����3T[ᤆ�����G���}�Z�5S�ؔ���i�T�2�坑�w�'#�4e��N�d�����Q���s:�l�����A��c��(���s�G�������5�����=���-|\C�⍞�u�x�u��妄��jg�c��?���4|?.�_/����o�\U�G��ߋo���!�m�bq�&8��?./ɥ8}xx���bh\��{��~�����v}�n�7�A���j������	�4x2RzT���e���8T�Q�D�/�EٱZCs8��CR��A1G%H��rb;��l�d	[ϛL�OL���А���E���/�}�(
s�� m��#��b�F$��*�j���gc,�������^J��1�Q�'/��Q?I���g f�NN��}��Ї����'��_V�_xk�^�N��}kHm�3�'�h�B��$nN�	�svy�y;2��K[�r������F�<�t��B�� l_�&��ߨ��]��ʱ�4��;�i�Z|o�E��P���z*_KhŇ�-��H�ҕP�ڢa�K���b����g��{CQ�VY��)��o�bY-u��Q8�AY�9�@�7����ڥ� 	7�>����n6'i迹o7�o��˴z[��<�6�e�������	z^)���G�60l6h��Tw��xǖ8���F?�Y�%�n�A�$�Y��s��4|���i4L�dː7b�g�C ��Kz_�qx�z�� �TbB9E5C%�������v��墨>Z��C��̓�%~�N�i뻟���m����S��$��K����@<8^\���7�����o}s�̆�eDm�Yr�h�V��G���K�ʄ5�dYm��YcM����!�v7M�8M��ɀ/�y
�&|O��k�U�Q�je��"f&U	��r�kv�G=�.UH��hS͵�TO�%��~#�E���))Ѯ/C�>���7T��+c5��b���P����Z�Z]U/���;�=��Ւ�+�����.U�5���
{���E1G���gp�[����a�~6���0���$^�+$�5��Hͮ�'�S\����f��ް�=�h��:4С�,��Sw��s�2�
K�� �x�2����4c���ו-{���L,�P�����Q~����N�1�8����$��
�����TTo��_L}�eU}b�����8T���'O\l���3Y�A؃d���_� �,��&4��A��g!��*RW�0�Q�S�Z�du)��u�gk��S�q)M����m��+�l���
$�d�v�ZP6�'V|B�.���Z���J�8U����)X����.�"zVf�R�D"�Ԅ��ǥ�0P(fhЮGB_�tX�(V]�Gl�B[?W_�ٷB��nS�ˡ]��jV}�(��P�m.���%
�ri����r8�]�..�Cc�������e��ě�Q`<>��������ƾY>74�[�YU�6�@"�e[��_Ė��+�=Z�d t��54���{�k��}�V�F���뇒������5k(�K��U�q��'Ƥ\<&��Ul"W/F�}�O^�Tc�e7K��*s���à�����!s��9�/�e��{YY*��G�}kY�~��_[����Vy��G�7�������?�g����˟�xYΟ���c�o2u�[ 6���:��Բ�(RBG�fR��g��6��h+OB�2��Ěφ�Y��^׺�ǔ�L�di��4���L�$|Mnw*���D�F���E�"'�pգG���"��H��S7������c��E�`SA[́lzS<VE㊦|�T�SE��[U�R=�J��M���P��7�v�X����r�D�s�������X8_�`9�K��-���m����OR�^?�L�>�$�o����Ϧ�����9.�%�힓l{%�8l�:O\���wQ���m��(�sȑ��{������oт/��·��K�P����#^!�%O2��v$�6�[y����^N��CN�R�~�=���
�gCk�X;�zM�KB�C�R�}a�8��q�}E,���B�+G��_��x�O���J���߇/��y�ʬ�����	QǊ�T׮~��6-���&���)W���Q�b	���q�	��p��P]�{+ήnQA�N���dr�4UR����̭��&�WRIZQ
i#Y�r=��]at�U 瘞C���v��.���E��GQ (�G��0��.�es���^��t=��~��$�7AW�	������������hj��)��Op!�A�	����⳱�s�֗\N����1G�5�hL��m/��"\\�`6;�cjGIM9�)��NZS�Ã�r*���5
D�o��G��J.iLI2x#E���H=��Fi�"SG�rhg�'b!U��"{)�K��(�|K��<���*���Z'
}	%h��%T�+��J!�!��KK�Z�75)Ih��4]`F*$��>pl�M3���1� ��nA���ֽ�3�:��v�SCGCU�ۋ{Э.��7Mz:����ͧ���w#�7����U���,���q�yG��� �w/G��m�����^�=y�^�	�������.=�A$s�)u����~J���.�%�'�P�D��c||�7$�')Yk�7��ŉ��ҵ�U�+�x�HO\�(M��>Q�ܩ�m��B���Oԭ���j�]�Q_�_�V��b�}�ŋ�?.Nn��o���]� �W�.}y���Ot��?Em�CH�i��^<�nٔAK4̪6�[<F������;1e8�~鉻
s&{&�4#}�b�*��	lY�y��j�LT��Ob�at3��9穓`\CC�*��Nϑb�%�コM#[�ȝhus�	+ 2�;�̡���Հ¹9�*q+�������f�~>���jTZ ���{|��Me��T���^@��Xӭ>����������"�#���>��~���o�!^`���?/�"h��N��-h%�o���p�f����};��ia�p�!A7����T��,J,����8���������3��JiV�+��j(b���yR�xW���*<Ӫ$������ U�D���Vt��X�&8�(�K��	L�ہ��}4eT���� E�Aˋ��S��L�'�n
�q M>���}@8�%4�X��8�ė1Ц�������!K�8�����#�@�%#�p�b��CH�Z���[�D��Et������OǛ_���m��%8΄�������
m�F)���(���X��e;	Ք�Q�����y6Yش6HK�y��vu�2hv�Ϋ�(��?��|G��Սjv����Ko��zG��[`�<�Fǭa�c��s)J���*���"�@�5$�~#�nlq��C74���$ �+�*P=���\�K�i%lG�[P�-*���ch0�([P|���l�	�4b�Qz{�;<�2OM�mgeU]�v����L�����0Ns������
c�R49B�U7<XI�2�4��������x������/7����۟��7�^ox���hKU}p��\�5��?����C�.�A\O�ՙTlEP�S&�MD^�,���gU��L��q�#���u��|�Ŵ)ô=�	b�;%i��x(��z��'V�P����WE9M�R��9��Pc	J$�|�K0�ǊZ�ThTs�[�V*L�����S��'7`�EBm���p��[�(����CYm����(6w�P�����S�� �t���(=5?8Y��@�n�$�i�:P�O.I���@{�T����gI���+��^vE������t��~��3����|3/�^�u3���F*��0�fժ�JT_�<8���}y������Ev�HA-K��Ʃ��yE�j��!�4�5��B�d��%]���i �<��YJdr	����F�sx��-I�Q �E���j}F�ވ�2����.=��.��=N)���+���ŀ����ZS�d��P}�Cw��g��l��lx�?��Ռl�A�][�����csA��k0y���{.m���E�0L-�c�ln��uwq����@B��r�Z�7qt���i�c$��YH}U��H�MV�X��!b�M�"o��K-y۰E^�0�͆Ƥ����mN�|O�z�r�<{sHq�{N��z���<���th�]���b���J��Ē���s�˱u��EӺu�-o�O�{���4d%+�B�%�E��vgҤ�|ҿU�/V����-4qP�B"7e��!?���U��74է._�$?�fx=�5K�tcW�}HV�Yt�����8C߀��,����5�g�O #tB��'V�ul掹jLf��>���.E�>��t�M�&�������QH���ļe��r�6�
�Q[>D">��9#�flٍ�;�%�v�,j��1�GKl)8��-�9����dk��Q��l������([3�W������v=J���k���`���;*!)��)2��Z%�u�h䆢���] ��~��ۣ5CjyOk�%�p��ف����ʒCd̗����"�Ч�bٔ�.6Ų�l���k˾k��l�ȁ6d�H�&Uz��"�21�j���z��I��J�t���xYx���w��x�B�4��l���ob�?�d3�?�<4����s}����(��'ǹx��5yTe��R��s.�K(.聆9#�;[^�ǁ�5ȓӓM%͐X��yE���Ef�ܴ�<=����0Q2%:j��s�A��@�'T�-B�J~��N��ZU���J�ޢ^�Rg�70�ȑ/-g�8$�\�x�^W��ѲB�'jr�5(p�0�RoFT�bI���X�{����(�ltD�W�V�W͠���kMu�%-��#B_�E���]���g�ZVG��X�ְF�=���C�A�_�Vܧ��,}���9��H�u͊� .�S�t>��}]��NaDjޠ�49�Fu2���&��4�Iq6Y��ibq���ۖ�p��gV����s�$���-��2~�䉪>�ţ�����۟�q���o��^��~�����p���?�ͱo~.��/A���Nz�v���g0�1h�7+	��;������?u�g��>:���6�uu_7k}"6���|��C��,a/���F�Q��g�`���:	�����2Ֆ�G�u�J�2d%s8U2�q�R}z��Y��G6�uZº?��>�cΔ� @��)ǥHj����\Z�P���λ/�%�$E�=�Fu����b�V�*��`=����B�r/ǛJ"v�[�Ҭ:8�����{�Xb�s\?�h�[�鉧C�FAn�U���8�7��"eU5̩�.�nG�pX6<�7�5{�c���`R��G%1O33�A����{LЎm�E�~d������Lb�8����\B����v�g�i2�3�HF$}����1e_Ǎx���	I�<���k�y�(g8��8<"��<�y�1 �I܂v.��c"�w����KRmjua�d)����L�)�6�ԇ��ј��A�I�.����������V=��q-�R��zb�ʥ�jΉ�I���y{r���GŊ��΁C�(�ig>-y���]��;e��\�:�~p�fu�2�����i�DR���
�x�2�*y�E��bY�t�87��jr@�l��"��UPi`v5���x2�M�=~%*�ܶ�G��,�8��ʃ��u��CC(���?�w�N҇/�K8��'�����k�YB?��8{����L]��C�|'��L�"(8�&%jZ�6�Z�I	r��u��f��<�B�j�$�C��]w�|턩sm�������7����ط6�2�(�L�L.qd���:�*�P��d˛�v�GV�y'���=�2%������hL��!��(#�f)� �N�0E�6�,o�&`�{�W��G�����x�D�J]&l�d[ઔM<%��� ɉ}�*���� �h�������8�'NR�y�)o�	d� �h��o襱�0��)q�
���0��f�r��Ǆ\%�����vϓv�ں��oד�u�J�L�{g>�Jҕ#Q~�6��X����y �q�BB.`J�L�ڈ�:�u�ذZP3�R"!k��p��Ť�1�2�#��<~�bmr�&��8�e;�n�+�ΪL�ۆ�*d��*�kR�C�
�������Z�c�N�?)�9��>������	b�2M���i�6�߆L�����$I�a��A����;�CCV���%,p<o�AlDAExݒ��Ĺ�"���&��h���y�D��d�o��ɍQ�]ޯ-����0����Q�C��U&�.��Iw��-dW9I��_yi�e#��0Gq��������+��#��C��?Ã?7�y���$���6\����=�u��5t���~�+����nZ��y����!7]fi����u��!+����ֻ>l�),aG�ؙ`�<oBhT.$l]�8)IB��9�}� �������vr�L���g�8	���X�d�r����Nr��Җ�k|�vu�mZ˨J���lM���}��vT� �$&�tY`�.zV���UL�)1+@�!��Uכ�|�����|)$5��0h<�h��!������Ȥ�K̙ȹl��9�n���:��,��+A�0�2�HH��P�<�u��<)��nv2a��3ӕ�9�.�_}�x�т��)�۱F��.��Iց(�EI7�7Z��
u�KTA�6�UC�=��� �y��Y�cR���2�6��7�f��%�ާ���9.u$J؜@�
�h�$>>%0����ш�5mLĥ���L�ٚv�?��37�ƍ!���5��O��}�9{?)�z�$L1���B�A�Y�Y�4�1�5)U�;0���\o�
E��>�آDc¢��������̲mQY��@e�I�^>�y��QǮ���#������&H[�����<�V��g��D�b��0=W>Q�#~��C�����-";�Θz�UF�KF�!��ή���s�O�{p����~�f��{�����=88}^�x�:�(��w�C���ط5vm�xs��\�����Iv����4G1���mR����#׶j��aO?��8Q�h�{����p�b9���W���fVi0˗��Iɐ��%���Y�|�<N��PE�s�Rd_�T���-WH�����K�����P`��	���/ �4ٶK�H�E�{�QY�1�@Vq �HQj���+��� �|�t(m��k^֯_H�v�����
�yݣ$���:�wڵq��,IXr��ĻSq}o�jr�Ib�t�d�(<gh�6�@���*H'%,��%]c�O��qlǡ	ݬ��3��ᔼ��:���f�lW��9�M��ǆ{T:��+J$�}䡠d#$�yGLJ`�~��$v�:Eb*��(�q]s~G�]��2�{$�~]�d�n��/D�`y�doX&����׷eM���"0�$m2���a�l.�4~?���]	Ƶ�Q� ��Х�T<@��`
}��<����2��Η�}��#��u���z�U�=�K$���ƷCI��0����`���q��YwR�T	�J�I�@9�����DCi:�Lw���ԟ4Z�F���`��'�w���?��(�ā����4E�����<0F�9��e�)o �9��bhP��,����N�������S�-\�{�_�h^s�~��'䗪|��=��FR���9���K�XdWyT!i�y�u���}��'�իߝL�f������P���t�B�d�T�C~�]C~~!���S���ݎ���=�ɽ{��c�x�cB�7P�%;p��ě����k�E����s<�,����I��}�ǭ���6��|-�`�VJQU��r^B)K� ��qU�`u�I�ˋP�n�D�Z0z��0�:+�]?�}� ���]l��͠��������.��;AÀ��J�`�I�pE�>�"�{{�ٮ`�lН�����;�V��Im���y�7ޜ�i�ز�NpK�n��晓�se~eRR�@���&B�F)�� �p��F��T)����LHj����x��B��ۥ*�B8�^ݓ�D�³�A�`���{$�ް`'��f|�d�R�!�.�/�Jr*f8�G|CJ�)Q.T�F�0��q�ړ�7{�tM�ˣ���[G�*#9��ǁJjTdC#��$f�\�Z���n��%��>*	��wI#oܜ�Y� jؑ��*�EI�B�����~]!7�\m�K�-����oI��кR��G!wAE���ْ���e/�$Ĩ�y|�
�K���$1EP�sZ^�Ī.t���JGCP���Vu�����`
��+�,s0�m�\��s��c��3ߏ�NGd/N���P�)����,�_�����?�6��x��5E�ͽ�x��>׵���������Nd�Tj2��%id���T1J5~���
F�hIJ�����,[J��Z�8
L����M6�r"��%��k޲��T( 'k���#Yδ�6)]+�})*�x��+=_�Z��,x]l��IL#�r�_@�c��ڈ�����ńD@��d��b&��"lT�l5�R�/���c����T��O��d4��c�(��Y36x�{R�B=	�_1��!˞c���7�&�Q>=���f�ӸQ)$�"h�����ɅD�Q]�����Ċ!9���R��f�U�T�;���z�Y��;{��Ė�iĪ�R4�%_�xL�{=G�b4�F6��*�T�T���D�;ϱA�օPeO��X ��G�b��B٢`�)y����-TցK�&L��57[@���0�D��I>��N�Y����4��n;�q��_�,k[yT$�l����MB�1�_?M�5�a:m�&:�������R�d]!+���Fj�ˊwQ;;;��2ޣS]��^�ry�M����1��������m�u�� E���7
+u�(�h���9j�<+w,K��8?�B[�Oy�<s�^ks�5>yЕ8'cc�%������a/�:���<`	���l�S�����t��i��-����q.�7���u'��2�'_{���f�nD{�e�f��zy�7�n��}Sp�����c�w�z��MsY��MH��hxbL,��X�8fB�>'G�J�c�2�V�D��1̮��v��Ӟ�q��4u��B m���^k� �[r��SsM�E�D ��z�->�	-�ܩ|"���8�nJS���,��{N�+E�%�fn9I���P�`v���s����������I������4�Z)��M���}�������tTW/)7d��TaP-s�,sj��콒$"���(�%O�E�DN�&�����%Jee�x'�|ÄP'�G�U�{����X�%K����O���)����tUm% �͓����=�<_�$9����=�2@B)��0���m��n���B�����Q�M���$e�v��4��C��^�($a�/vyvY֮ t�lO���{�	�#�&I�N	����z��k�pDi����.�CMbp�+~����I!-�8�k;RH�H�TvF�c�a�4�|R~����@�����8�/��]�?kT.���v�H��������۬��S�zY��^��&����DS���|�܃�(&.x́���)��c���C�=7@��c�8�01�tE�Q^�g�r ��is�K�Gp��������b�����^��zp�f���o���� �͇n���l�Z�nȚr��e���(���M��Td빘X��\��DI;�6�ѻ#�sc��l>=�}����������Y��.+U�j��s�09�-�(d��(�rW<�a���@��VzB!Q��~�%5����s����V1(~�wgܣ��ϵ�!7�$���4�萳�U�N�����o0m];ř�`2�\�+{O	1G���H�G��a���$@Tb��J�8���bΨMb�Df� DRP��Vt-�?ML�R#�O��j!��-�o�����t��U1�٠36k��r�10�%�`����kdKx�8�(㼘(SI�N�:�dd��#�LÐO��f���Wa�?�4��#�QY�<�()	���ce�TE��5���d������\��!�I�l��%�I~�����X�۩I��\�@�_1Fr�!Q�>�����\S~y�����*[W'&�җ���6��#�w�����j.�a1�s��r����c���]=���Է�($�Y���mzQ�Ed<���`�J�G;��4giz,;�Ȍ�呻�}<���J���HBoAs�ݖ�)1��`�n��R�F�5�h��#�!\���ǎ�^���p�����ٷ�k�:���w��\܇/������Y�x�g(�F��ҌAk�q�s�{!�s���X� �$�]�*��t���D����^����f�I�qb�G��t�Ԯ$t���&��������[=�vۇ4�,`V�udbˍ]TI[В˽�ul�Ak��]-�k)�T�f-�,�I��� ��X�n6Ht�l�*ۻ��a��X�`��Ⓡ�'j)bN��C�R;kA� �5[#�5j�^�GU��yǥ)m��
Y�I��iY8[7<NG�^tb�S���%����(�@�f+%p5mtC�XQ��`�QJX6?�߶��D��57�LR!mϡ�0h9
S���jc!�dR`'
���S~g&�a!W�tb1S,���Cz��Ф�ˬfR[]�|��<����v�N�<!�M�I�6W���Uyͅ��!_��r�ZW��b���I=�)�Y��N�y��:c�rS�t�ɱsK�k�@��g״�W6^�A\�F�D�k$݊���Y��Q{גI�Y�q�%����!�z��BR��з=,GLt]��K<�j�\ӆ.��o6|�y�dx�뮥nN�qx����ֺ�~�I�*Iv<�����!��v^7OȘ�d�J�@T�9d���C�ׂ(�A�6�{Xv^l�g��&ޫ��w�ò�T�x�p�̛ᵀW����/����E�'o���?>��o�\��ɎBd�s�$�q7�(�7qU����Z����	 �I�:�^���0�|��ڼ�xcn�|�te-\�I��+�8�K��
"tr����ރ�8�~��2Liܖ5��!M��T5W��%���h���!�����QM*w�Ӥ;w+��3N����	mbB��]����l��h�Pn��G/~G���[-]c��>���bΖ��:\P�{����4P��>�$��Bզ�1���Y������e;�>�Y���\u'�Q)נ��8��+������ܘ$5U?mNZhŬ�Qh���Y�[����?m}l��f����x*A��!���D�Ĳ�8ւx�U��L�)�1k�@)��FY��j�
Mw3�I��3�j�y�-C5*�3�&��L����`� l��0,��d/���'�S��Q�7��}O����w�LTe��S�y�͎P�#b��K"qT47���T�V��.���	�ᙧ��'��{w���y�՚�?O{�d��B��:�i�z��3���Y���.���d|�qMoW�����7���'�P��jχIb��3��d�e��њt-��dI��/5�81�?Eq�.>�o��2~�����o�O=w��[x��w���W�Щ��ʃ�o��woo���o7({�}&�ȍĥ�V]�Qj����8��,�rm�X
�\����Jj=9d�i2�¨�e�|2�R��_�l��oyH��X�K`�m�N� mX+&s\�x=U�r�<%�����%�e�_���(��L�n�8���5��%�[6j�V�D�ԝE�QR&�1�M��#��"���P�7meK���v-��ɯ�ތ�}�ݖ�7����Ę,f&_3��������"'XQ�{ ��A�=c�-I�q�2@�޷�\I�Z�=
W*]�{��-
�
')�P�6��(�Fʯ�-
ZY1�����3Q~䦎��}�rL��5�ig�yQ�[bʅ�-��5����g/j���9�e��鐅ɒLXN�
<�Dh*��v=��(�$S����[���EU`Ұ��?l��y�Dɥ�1���b�rh�s���g����QT���є�`zOG%i*���J`r���[a�MY����P�fL�D����pr�&Z�K� 97�l��ԭ[h ��Z�=����3���{���.��p�\q%G�JYŜhG����RhF�6Y��ES���>[÷c͇��c�<
���d��=��M16��{�c*��c?���`��Q��Be�$5<l>s� y�Iߧ�L
�7D����������'O��^x-�U#tv�o������m_�5_��RO;�Q�f'�M��7�NpA��<���G��jN�R35�tڈ�Z��L[�����/�V-{\C����[�����ld���Z̠;D��s\"i�����O��UD"/�he�`1H�N���UQ�1�'�&�c�A2ԣ.�a����%Bt�lQ������aɄ^R�
7��x�k�AA���Q�(���ZT7����\qY���e�"@�ՓUGJB�V5�)&������1�3��I����T�D Q-�������J��VT��������ٔ %4od�W�jz��M��,xR��ͥ�~@W�O���x�m�C���%}'=�A�������*ق��mL�]�Ģ+����2��Z)��YK�y�=-��X�h�&��������F\�4	!XPG<�O�X�k��LjB��vO��(�<`�-�9�ӝ����)A�[����\FK��4����� '�qITUq"�Q`	�A��҂��ě�|mZfv�c5���1O����w�2�]fǯi�Q���笔�=�s�5���8V䵛�`�cՓ!T8�y������§>����wh�p��!\\&h.py)�>��q�KN�f�a��=��������~�%嫝3�D9c���O�	J3����M)��@!�v0�WY1���i����@%�*��}���j�76�O�Y�_^<��Η�=�x5�Z�;/�;������b���D���v��`z%���C��'��\���8Y�r��(�f3J�#��Qdd�2Y�-�h;NH�W��f"��=�	�+���6&�lZ4�q_!�N.p�Bk�B�po렞�$q�a����$�ʽ��I��uAP"_�;IR;���%4�x9l���P���v�@��%o�BǓ$2�(H�uM��cCj�e�m��kzKpduJ�a����L���&&�F��%J���-�M���v��ڴ�EU�L&tRU�8[���H������*o()Ǩ����#nI���\$8[Gh��̯�cu��i&�:��X�ZrBT�\��m�e�F�+3FF�ºB�cP�5E�@�Y<�kŕ�'��{v�Ǚ䮔��{����9�y9Ve�=D��7|��E/)Q8��+�y��l�'�QJ�����c���L}f�!L��S���2P'@�܃�ʥ��p-��(�SE 4AQ��wjmZ������$���������td�^�8��
��^�g��R�d�/8�������{د.���I|����x3�Z�4��,�ʻe�cA��HS���:똃���7k�����k�V�֘e�H楄3��Ys��cE�$�a?U��y6Ie����ݑykk#��p��S�Ǔ�\J�Ѐ���*�G��-��O�x�/��w���pt�Yx��zsvNN�~�� N��uH}#��P��h1r}�F���8�}�s`����Q_�w	�Ɠ�'�����p�[JȵưM#4!�b�[�����F�B�R�7� j����L��6)�2y��UKB���5��� �orC?�|-�5�)�v;�C��5[�}�HW5�4�-yG�4"9�5�lr6�kK��H_	a���&�D�a�5,����B�Z��m�v��1}�Ĺ6u<�en@$��ErCJ�m��jVHz.]��I��8��cŊj�_:kᅳ _zZ���E�q�z�t�/�UO��7����2w= 0n���jb\���|DZh��-JAR��֪d��G�G��[�!}"�.���$;���95H�L$|���������k!��S偽7Ɖ�l�p��8�2 g�ш��5��nZ����$�ܒ���~����nP�=7˱n��a>/y�ɻq�8�c��ɫ� ɯ�+���a�����{�����P�A��ީ�%XR�=��R(1fz"�
]I��Gͫ��Z��>okc+7��q]O����ŭs�[�%�Pb������W0S�Q�x���~�o����'�O��77˗�o�1� �^B盱�B�9{��.�o�7c'�9��i)����Jyw���V�FBFw�#0�~�q��ݷ^)B��M�T�Oj�(��7���T �h����Y �WJ��h}�E�Y9���
s�r�`��	��� 	.I�<m�B�z��*�|��`6�Z�Գ�w>��ۈuS��{A�|�E�F7t�^uɤ�4�
&�^]-f$����ȵ'q�f�(j�M���7!��J�B���Υ�!R5�^E'�Uڝ��������iܼ��2�^z�����}�n�"'lKD�g����2���``ۮ�G����5�$����1L��
6�7���8�M����/�t��9���lߛ��R�V�J�R�/����"����(��܈֧ݮ!f��zy��B��غ��eO\�$�Uz>�M����څI�O=OI��^&�����[��N��� JIp�g=���f�
NN��`�d^�ť�w@��е�T�6dE�&��b��_��h`�l��ym��� smnM����d�sK��9�۝���������5����W@KC9	���310���"c̰�r�Ʀ%�E���J}�U�Uku�S�|��?���~�s�j�N���]��>K5̧(x�߬�<�:[���9��d�jKCޓ{�^����7QmL,�.Fbe�MҰ�x�+o`��R��8=�� ?�g�w�W VhT�膤wS�5�$K&I�iސ���9W��.b����ӽZb�e�b˴�e�#Gv'M��K�:ơ��s)��삋��Ye���Y��uÊ��p�tL��J��y���Dr��ܥ��d-��Z�K�;�d��F��j������0�OJ]8E3Yon��q׾P�yW��(\�o��O$fg
�e�@�m��v��~5��h�
�]�`�����&!A����JMi�Z,tS��Q�n[2_C�X��e�=|��4��1����⍽z6L����#Xמɸ�\����Ҵ�_S(&��C>.�<�sV� _��� �W�=�&vlK㧍@�gcYƿ�9���1�
��LZ[k$�7�+�-o
!=��㰘��Y<�ٽ�R�f15�w�`��o>�a�Y絜� ��\P�6<B>JF~�y���^Qv��;߷�I����5z*���VVԜ�2��B,�>I�d�=��Fϱ(�]�C��R?����ֿ���\��=_�M\����߮��ˢ]/x蚿�7���mX���ZXw?b�,��d�=\nA.@�`$B$׹�G�\ՌU�]gAoY1��)��?�zVi`���e����R7��w!���F�t,g�X� �	iyS9�� �z�`�B�]�TW�}�E�������Jv"���8�t���s�%�4He|��D��yC�$�,�Y�W@ز�L��b3����
d��`�2oՆ#�/fg�{�Ƌ��8�4�D����,�l�XJb��Ś�X�i k�K�vڃ��3xжp�V��&�WD���5V�5�xW��Cf���ˎ�%@�H,�ŻA���Nj5�2�˅D-K�d:Sd�e��}[����{�P��M�A�zK�"[^V�8Q�lL���9���Zq��;M��Q1�މ1�vW}�q�5u�5�M�� ��=����=9fP�6D����w�w�	���)�Ԝ�m������'�C��%~��jV��Bߺ����{3,�h �ӎm�Iߴ�����D�Ъ�]��E�:O��t,�*�Y1�fM<��d��f/%+!��^J�r"��� &���5�ZE~S�]��șh.w�o$;���M�cE9�����W��V���?;|A	����7��+a6?��]��Y>N��ҾɺI'[�)�֨bK�BIE� 6���Y�[Hٕ9�Y�	Q�R��mvZA�א����i�^���n�3)с�C����DpqM�$i�媺��ؔ��dRW�-��I�u)[��ЙЭ_�N��]R��.uqXs�$MBt���*ĬJC�w���7�'�\�㉘b ������A�D�f1+� ���Ж���bҽ�)9���&���b�Iw��)f��'*g	��W�]�pѯڄ�v�Ǽ
땐���lܵ��<rz>z�N��e��Io��22�;z�;��=��u3
g���[�׺J�����>�"(9!e.5��q���Q�*��[�f������k���My׫�Z�6'caT&s:�T����7(��|�jS�y2�('.xs[v�g/����
��bG'��#i�~�ʣtB�F<5�[3�..a���=��S\gN��ٽy'�'N��=�,8==�^�FZA���p��1�+��	����d{�\�&��^����Vr�����+%6M����ż�ܹQ����s��8��,T�q�GjPV%{�����>�۱��Aw���܊Ο=�`��>?�A��^��'C�~>D�s1u��7,�j�LV	b�V$�/)j@�.A�����`$�m-������B���y����W������B��ꦁ||�V��GGv��Y��Fi�ܩ�O��2�M��g�'�&)����ִ�]�T�ɼ��7m�J�mM�`�voE)t���D�����nd��5O}M�U��h'�<g�j"|�u��FO��_���Kq�L����ͪ���~"̙��$�
*y����8&��"��Q2� ٤fVע0tH�\Y �O5H�ڑ���6��yr�u�ǧ�E�T��0q7�5��O:)eK]U��9>��޾�z�$.֬�ۢ��k���5��%��!RzO%瘃�:W��k�֯��A�%:$�G�'�v��C��{-+U�,���q�U���my�;��߯S��ؓ�ܾ�w�J�A� "_��>�
�ɯ�s��K �1i�
��25�s�|�V���N�H/���baW|�e�{�̏P� ��/pXpY��l��U\��� �����Pq�Uڿ��R�k���ԃ�L�������mu����2�?���J[1�Za�'��Jr8�\$�p�y���H+�,TN�ᨖy*R�\�;\Փ t�,H3�����ۼ�o�-g?�V��yo~z
_(|A�k��(@������6�ݱojj#)�C�G���	���ٹC\��9�eM%�����ė�T��4�['%��Xr����c���[��M�W�9d�`�����抓�"�Zgk4e��(`P� L�)�ߣ�1��&����d�S��
� Tiꓩ�6�����k��6*�};.$�.¤5�J6��R��JB��5*=�6��v�|�Il�ܠ���}��yF�\$�g��u�㺃YAЈ�*�</Q;k=
�V��ӆ+������Q2��h�T����-슊
)�Qq9�f���D��Z
|��엲���x�"ߚ�6S��+��0��ʓ����
��Ne/}��,Gj�K%e�Pi+YY���d��[�k/��O�[�&�?��i�YҤx���AjV@���E�	�����Ī��xt�,�q��m��.�O���#v~�]��\������"ϋo� ���k=iR�y���pl�ĭ^c!q񪬳\x��Gp��-�=u�\5��ڼ\�f.}+��G��ʧ�D2�����qP'�ڔMf���Q�޿�������k�h,#��lyu����'
jV�B���f�Dm�
�*�*5x��۝;�C<HR���x���>�+*y�0/M�p+�Q&L�~���z�7�����������i�����З�_�yw���OR��t��J����	]���i�&s���?�Ŏ]����.�	�o�g4Ɍ�����N"u���ͳ�29N>^'�Ð�n�ט�	{�)�SD��,K.���hЉ�GڧE������\��r�*y�t��C�lx����zr���U��_����bw��������ըoG���j҇5�:
L�fJ�uϊ�.֔욖x�w�;+��%g�����$q�8.�`����� �^�����>�H�?u��`���h�L.�d�G�,9�}�~[� �[�+��|)�Ňg8.sn�kQ�	����c�,?�L0W�Z�Q��H�5�G���S���G�C�Tyz�enϧ�u_��re.��}-Wb�3� 6B��c��#���� ���|~]����͛�m�۩.Jj庀�>��x�e�g��g�>����Ƃ�"Q�Z��y�PE����5m�u߄�2��M��'�}u<��e�ݞ7�Q׍�f('�'a���޺?I� ��e�
�;%ҽ�R�ް�j0�@U�+jo�BwL�
k�-�&��6�\�[,� U��{�;��o�/߇/>yp6�w����S}���خރ��[�Z�݈Ƹ9g>�eHY�-�=�7�)]�l�&�.!�4ɴ�^d[�G�u!��Ab�����Ʉy���nPS��/��c-9͍����^��kRO-�:��7ߦ�,�YE-�Ӗ�X�%u��������v�c;�)1�'n^!�ȅd��wǥB�\&l���Ucۥ+c&��B�t[���fz�-�v�ޟ1S<�X��M�t�EA�čt8Ӏ,sj&�.*�!��G{r%%���RuA-�QXPc���A?���N@���޷e�?I'�2.�>+Y��w�I=deI�ħd��)E{��Wf=p�y�����1Z���s�Q����i��@7M2덟S�ݒ�)�����~���Rj)AQs�NC�Ӷux}B�u��+�r�q��W��%� 3�ާ��{1Q�g�1�l6���S8����//6��@�s"*�(��n@�@����-$����N��E���1�y���5u>��:ٟ�6	�U����z��l��0�E>�=6~!+}��NtJ�ZJ&�V4�}ˊߞ��S�>M��i�3i�6�(�v:�0�9J����l�I	�)Q,�PH;eRBe��5�3�;�凊�����c�m._�����������4H���tެ����.�J��,b+{�Ԣm1i;2iB[��5��|��F�m?X�%�+Y��D���C��n�V��qn�kH�:�ݴg��191X&1�d
ŤDm��0j��ʠ�\��;$�%���)�Ei=��-��ص�m-So� �~�~�o9k�Hb� j
���]`B�=7[�V�&�3�a�����K|�V�uu�E&W������S����cS�<�<M�A��x�s"ur�i�R�PgŪ{К�pQ���-���a�1e5sC-Q�K� ���G���X��u�3>�p�I*�Fg2=F(]���Bھ��q��9�X?�q��ǿ(�2�ę3�r���&��6��p��v^��a!����g�'W��z��y�by]��nb�+��QK�aHJX�6�)��Vб�(�3T(G5�Pt�>*_�f�!%<v���|
���H%n�wy��3��U04�,����@�P]�}��r*T��v�����{f.E9�+s�����'d�h�)~i*���!�,�Y����c�E1GB�>�A1���o�I�5v�g�G<J�;��εC�a�7e��+����'��v����z��z�\�3?�볗�v�ڿ�oV7c��d�iQ,\݀%��>���F�����Z�$<��c�nJ���Y %\�qڍ���B)�1�ʎQ�u��j���D��:(�O��>*x�#%�¦s�꒝�QM�n`�.�I�Y�gy^��(=�Ţ�ms+�$�`�#W�}ZpB�ԄG%�"9�Js�b�m�9�{ ݞvz�����l�̇[@��:�J'��}�>l_f���y0]�����g�#�j�������}�%NJm39���#�;]].�J��
Y&d�RNӒ�"�>���:�"]���u��ļ4ꉹ����&�8�����G������,`Io����QP[�#�r�r�X�R�'���%�T��)����v��Q�񑐷�aK1���n���&�]"�
��הG҈������V�����T*q���^�Q��I��QJ�+��XN���]]Wp���a����K�Z���vg�
�K�G�5`��1oDĝ���!�~���Z9I��W�"�v݅���V�{-f�|bi�c���� �����x!}�֕ +p�x���mu.�B�&[�Vѡ�
"��̶(
5Ri����V�?���_���~�fu��x��������i87�α��h���з_ie�����s��\wXz�Ķ-W�J��Q�y����}_C�y���Z��H�8Y�6�f&���˙���da�
��s���2��S�`\�I�=��$I(��B밂U���A����3�jId��6R��>hֶ�֔`{��-� �h%��Q��'� G�"\7��)5��M:�!>J L?ÉA�|n�h�.4S�̃!���p��JmH�dT�8�90� �E�V#��ą�(���yAU�7:��I�[ɂ7 ��r�Q+>��Xm�!!��,�_�� ���[�}�C~�k�:K�s�5���CĞ
Ʉ�.M��H���Z�Ie$�[P���;,��T �"�6�&��(k�Qޝ1������:���*���6},�I��c
��\s�#n�[�V����8<>��%	�����/kr��PłyX!��ap����T� �d��|t졛�+VVc'�[�S�MFXZ���m�n�n�C&W�ǳ=/,*����#q��{���D��2U� �*�p�o����HZ��N'y:�U��$�����bQ侢����q㙏w�;/�N�y�g���B��l�8�<j���f�]�݄����n��m[zP�}��2�\����s�JY!�,�HDDL�5�
�1JIb�D_�<��� �)�A0��/�!���*����9���֚�K���k����?�Z{�S�����s����/�����F��V��t��ˋ"�A#�"���鑹,��`�̈́�[���5��������B��x�_�z�Ν���|�	�l��([�"��mܒ�5g&��1�f�S&a����_RQ�<�����l5O��؟;�vW~߇�٣�n�;�)�+� F��^`��T�h�=��Z�&Ώ_M��^�����_Rз8t�G҆*�mc$����&4/����^�eD@�h����.jW����%�	�� �ѺJ"Zsƹ�o��]�4�De��V:݀�-�?Gk�"T����6y͗�`���Gl([���\��*�B����=�����~���:~�P�=��FӨ���V�W�B���ԁCa$e%�aj'XU	��U14D1���7�o�p/���#�%l��Go^��ڝ���F�H��Q���t�TP�O�F��/�"���t���h���F#�J�� ���Wo�p�Z�23ʴ�O���s_U��P,l�$Z=��}�WD�u-���Gn�Mw2��yvs>�mn�"�}���_�_=d7�]�WFțu����ϑ?�^5�d��0_�ޡ�es��)j�3ݨ�>(��K#ǳd�D�3`m>��)$�HT�V��ΒH�-��^�"��~|������������*�]�o�B������]�@�?|�����_���ﱰ4W�� jq׼(N�E�Y���̳*`���*��m1��*:T�
dw��gIQ@����ș�ur��.�"�TK�L�g�^+Y���S�Yy�r��	�!73P��q�o�[�MY�,��N�^�*�8�ŭ�v,@X�c��>�5QAU#�U���Z��ރ���š	j�Q��
�&�tcg�:Z?8j?ۚ�O���M\P���M(4�� )>X�:R�*�ܽ�F_�����c�vV�MiOh���J�v2��q̨���#�246��L&P�����6�$B��a�9�vC��4,e����=[Ӯ�B������|��{on �J����\�2�^�h:�C���Y�綞'+"�����b=9� S�^m!8�,=��� ��ת}Đ5_1�V���L����v���LD��se����^Id��^8�Љ�\��ֺ�y�M�����tu*T�iȑ뱚�x{~�PFQ������Ⱦr�e���ʔy�/
����u��{a�D�ߊ�����f����ve�޾���\<�(G �޾�<�b8==�W/��U�z�F�W���x�z�5-���ES��!��m��|,Z�{�ϛ�����&��!J]e�+y�׈�hx�]��8w��c���
%�\�c��5��]Y���P�����iz5��O_�~�W�?����{���o��SW�K�������/��ߙ/����R���3�7�ޔ 9Zz��zG�ඉ}���?��-�[�p�G�Q�w�& Q��<Y��Xt`F7��z���b (�ZS�@3��j�m�>�/4����ۧ����ůy���A��O���=R��ٵ: ������(.2h[tC���{�gI��X����R�#O���v���?:�.�7:�:��G6zv���E����X��5mg�k�>SV8f��E�=h`x�y�2�	t����vʙldΓd?�#"���z?^�6�Q�эk?&��@�E���Mݷ���;0��~�*�J�%��T���'%
�R�m䳃��d��1M�y:t����~�Zm����O.ج���ѱ�3n�B��k���	UrC}���=J�1�}[E�-���{I�Î�	E���E�V���uAWCx�b��(�o�J���ûw����������׋vYC�1z:�z������|��ƛ���z�����M��n��V����qQ��
;��#X��6��:I�y��B�-K�o1���嫿�k�����߿���@8�SU��E�b��:������r}�̝[��܅�k�}1���ҼUe�F��& �WK��׷�z�2�|�/�����;�ë�)��ټR��x���k��My�R�!6����#ú)Ѫ
~�ho�G�A(�zz�t���$��˸�!� ��Hκ�RC�4ԑ��}Ԯ^��T^�jJ��Ew�w��+(K��kZ��L��*��պ��7�$����@���?l���[��\�^�� �Δ��Z��j�g��^"6}� %��QI��45��}?0���:�1��-�y��d����q�۵�\	���Oϕ��zG��j���uI���^ڌ��Τ���e���A��OƓ�C���Y]u�S;oto*��B��ί1XJg�d���ߎ�����Ɔ�����i�G�KΝ<�11����=r����X3x��:}�x6���u���o�%����(E��(��PN{���=P3{ʾ��Fˣ����ʚF��3ӵx��� ����_��*E�5��,��g��=�*���֢%_�O�����q'��uq���ֶ�A�Q��[�I#�̅F�*̋7p6���	F�$�D&�5���0��y���X���oǽ��:e���)���տ�L�j�>�3؞�����|���eQ�y2��W�����j�ӲP� Ǣ�K�	ia �RʂF��p|�J��3��<�R��Y?_d�슥��D�e�a�bļ��{jA�\7w0���k����s� &�Q��~-�I�C/j�x�E�>�P61�i(q�ﾐ�fDn�^B���E=Kg8�|%�v,�j���^z4�'U {�+����^��N���r?v�|��~�c���"��"�n��]{�k`��!wc/ÞܱEj��[�������g�/�t_�6a'Y1�1����ӱr%ͼ|����qS�^(f/c��hG��U��y�ݼ��a�n��h7��^��n�
��
�j�f�k0"+g�5���xM�%R����y�0��>����_��b�X���k�n��m���x�9�˽��qel�M���wX5Nξ��zd1��q@eBGE�j�B�\ �
��G��OS��4�e-fI�ā������2���y^}V���<͗`,�Z�ʆC��՚^}�u�v�.ݙ�]4��V�	���Q��6��'��%�%�������Dr0�-���4R�`�"���i�?��|��v�ǿ:��/M�~ ��?�S�����~��o�ݛo��e�������4=�}{��������
|[<0�B/
	 ��V�3������;�t�,�l�╏P臷���J�{�M&0���T�%��f���z��az��ɽn�����k-�^��I��[m�m)�ħ{J���f*J��(�L+zW��(�=x����Rf�UE���Q�'Q5 ���Q�6dw��
��>�x�;�A+�cإ���i��S~3�)�~/�#�������/��]���~���gi�`�z��+:5�)���Nb)~�F��cW� j��L��W�Z�0/s*F�j�0Pj�g�yP��y�A�j��`Е���,=�hu���nê��"�� �vh��>B�6{ġ�S�3�Ҷ��e#�:e�yVj���{�V�+�^���7A�o q��v	~B��7���=��Y��s�[���o5r��������xi߱ȴ"�v�����	��ݴ�`0�e�"'�p'<z��PB��2���^�O4���^��q�R�2���Mꮽz?Rׁx�[|�0Ѯ��~o��Z��Z�k_�� F���ϕ���VV
�WC�H�ޟ��Y��,w�X���\�����g����*O����$���)�߲B�^I�w����[����z�3����M�'�Xh/j��f����K8�}1��̛��
��-���H,�76Ў�$j�w�P{�H(�I&� >A��La�ڊ NrJWq"�`�#��/lG��!�������Cs���@�4�@M��|����=��y-�i�g"V�adi8�!4�he����r�����ʹ��Q��=�VkQ�4tƇ�ܳ�uɳ[�7��B�aý�x���Xv�~��[�@���g���ES����]�Mi{��+J' ��\C;�"?�Ctk*�=v�K��f5C~���Q���� |ٓ���5̹a7�Pn@v5�Xg���nAp���:�BGs�?�?�7�ɦ���9�sW��Z6�@:�ixI�ui�yr
Xc�����f87�҇��{x)�ѯ���|��k�z�O�Vv��9[�IG�t1DNU��6�M�GMљѢz(2�un��
�<��1�9�n�F��D%4�gww�{x[��I�����E uw,��`�P��\���R#>Fm,_Zu.rۿ�&�.�w�g~{T��H�&�� _t�m�~��"�%s���v,��]xv�b�5���Z���1�xw�����O����q! �G�|??7]/��\O�X���S`]K�g�kW�jW0�Ek�/��nu���H���T��$��g�B5����T�Ҹ3��Q�	�T���������<�Ӣ��y~g�3ⓖ��v>[*���z2��������NĚ�d��$:AMyy�>����R���R<yx�0��ё�Ex�(o�����X�v(w��G�n���RPϳ���Pc3�|�I\Y�:��g�/��7��nKy��%X��^������s�G6��yR�O�d�˂9t
_�9l�:hy������G{���<�*Dd��Wu��B��(�#�����1#/��KJ��G���*�j@p�Gq=�߶���#�#`��5�[����a����s���oU�Zֆ'W�5����
��@@%�=��iP��h���j���c���/4��X�j�����`�o7"��]�d#01�یZ_OU��� W�E�2�a���rc�^�v߮��#Ǒ���Ԩ]�GN��=����C��g���쳢�Sq¦yV�6@��"��tY�S�-�E�i�(ݛuy��y�u�Y�i�.ku�;��~zA��I-��m�]N5VMRq�6�5+;L�$�x�&�^�s߃Y�����'q\�w��������X�~���:b�����y�\�����?��O������I����r:���;����#C����^��MTDs�)�	�dJ3��-d8x��=��j�pn�gXwP�×�f6Ҳ-�lԖ���#��T@�D�d�T�gm"ϜJ�'��`�	�fq�`�nf�*���)ن�Z���� e*�)�{eIT`h}KWB7���F*��~���BN���I%E�3D���d�|����x]��ˇ��	H������Ť%q���<?E�7a�	��|k������)Ȗ>YjL8w4��l�o`��톻=|�ݩ�`4��|��m5���E��"����Ma^�߆��/4��;��e��t�Eq�ky|(c��F9[s�`����]5>_>��z�^o�|0!��V#�ټ�Z�`LF�\���EԨSwpz4WN����)�1_>���hl�s���ma�c�{�{d� *n���Y8��M1��"�d�31(����JȪ�*��.���OU���;Ԩ@Ȟ&0C�*1�qI�A�
	�X���F&���솲�_�4"G��Vͨ�=���@)�� _PE�.w���Z`��*��R<GI��eY^e��N��mr�|�^I>��V��:O]e������`_�����(6��~N�?��iT܉�0�
��� h�<��z�� QE&�=�!4�����f��ʎ�q�ȏ7�b��s���c<���K��-ʗ���)|{v*<������/?���u>������
}z���;����g�z��G���o\Ϗo��(�f�o�n_k�9�hiUT6=��u���
�M��Wa?�Cnop�Ml�:H]h�V9L�ʏ����?d�S��u��z����_/f�����)s��7��s�}�5LIDds���z󰗻�^r*�bi�y'sQ;����bя� ��:��z)C?�����ߒ���2�{��N�~$�r��nA��z%�����`JX|C�}��C��2�O���>&N���ۼ��|;ߟ>��
P������15t{��RE�&,��8"�l; �]����A��J��& ���=�Z��Z��i�Li�̅�_�?u?�z���ކ�o���Wf��n�m���TC�7�^�lS�Z�f�3Y�,��x�����$���uj���4�^/�k�j��ag�[�}��-�S���%r[bթ�hN�hk>�����f��;^A�������ϋGC�`pg$�	�H��?ʬ���P�����,?S��Md��{�Ҍ���2X��>���]�~�x޻E%t����>��e�fP����nJ�fpVo�0�Cu�܈P%O�!V:�i�#,��e�L�^�-��r�4���\�J���Ff���^.���5�a�%8���5�c)�U���$��_����Z�5�x1"��?�B�ݡ�҃���?���;����r� �j�-$kɎ\�ε,�D3��ܳ���nl�G~�؀3n�s(�k�z�5�����TA���~'�~_��P�����pS̛UG����������<�I`����ьr���-
���܅;PHI�g2����/�,S���{Z~$OO�,ro������^����=�q�N��p���b	k�k�8��7�v�K�*�AC~�4k��7k�!���y��>�����><�~�.��?d��z����ƶ�])�qP�3��M����Q�e0J�P ��΢��40��B�^��؟�[�}��
�l[�7j�'�b3g�!�[�L�<�Q����sg^����W-��Fz2�ޑ5���t�Y%S�p��Y�_7&��6����S7c���Zq%�G�|��1���H��ӏZ����^q��P�5�^�s������
!��x|(:�c����6�"J���W��g�q���g�(F�8��*熕k�
7�mܶw/�6�V�����T��!�������Hw,���
��(�=�[�*�\��4�F1Dfᑣ�eV��:?	*���, F(Y*����=���m6�=�q]��7�s�+{���F�����������G�����_����)�����Nq9?�����/ͧw��KٜW�6S�vX�Y4������>�j1�:Յ���E����6��=��� Z�����ꅺ��+h*��}��·�|��m�^ͯ�3a��Ԭ��1��6
�C�Xl���CQ��������l�}��+
�5=x��\e�'�J 2������[?/_����Y�Կ
�i<�c��S�X�.wd�4:)�0ރn�$�_��M�JáG���`	U��Xނ�^�O��S�Q��>Hj��X�K�ȣ�N]���y~92u��2L4wYv X����xO��ˇ��-�ZL��mpٓU����|�$��.���YM�er;�������]�|��#kh�b4V.��0���Մv�HYt$;�C�0�R"���HY�R�Q2��o���j�U�����ߩg��ٔ��P�^���{��cp����������K������ah�`�'�����Q��=Gy�;$�eg{���9��k�*��2CM���LK����(鬕;���U���m��aE�`.<�a%�����y�-oU����wP��+%�}i���9�7�w"���R'X��*�H�~�>�ax*â\��s�5��<rR�l�)֋���*����=%d�_�9W���(u��)ʟ\b��������w��<=�H��>������|щ<�-�g�\��t~���ǯ�Z�;ԙG(oҼNT��$��y���@��h�Xzu�&��d�.���`qԉwf��
�#ʮ����X�Y�fx��͡},gۉ�vM�b��ڭ��N��=���P�*�VEUlQU�vo�8��v��+�Rm#	l���������}W޾�L��b�;��>�I{G>V|*w��vh�`���R꽭/�=5T�B��z�~
�U�] �����龻v�����dyҒ+��C�Fs��:ۅE�wr�������E��'�;$,YS�g,�R��j���|�|������V5�7��C�*�|M�#Z*�yD��Հ�T�h��: #jpr�s�AHF�*�g�v<gO�ʛ��(�\��p%V.���#'�	��l��>k�q{�.��t<�9�܍C�>o����о({�ES�~���VC�5�Η�pxQ��f �^�7<Lf=Ǯ��p�� ����1����%ˈ�'��G�����zQ��R����ƽېf�9�_�7�S�l���`�AI�X�m�0KG뫆�6�BE։�@C��x�a���gȸ�V��HAʈzP�VR ��4F��K�� ��V�l���;��7�7=�wG@�4�A�p;�FS�
^oE�;{�a�p�2�)#�o����o��O���	w��Ǐ�����&-���r�����_�>�V�� �?+9�D�����Dn���P�ތ�J�<���}���B Q�1z�C�/�v���LD���D]FCZz82y��L�%k���Ѽ��� �k��A�u��9�F�l�+�2?r0[,g����Q�~�/9\�P4j���g����O�$���坻�����x�����>�s��r?����!f��A7��;=f��թ�r����7o���<�	�m��	�7E���j!���N�UE�^0�=�]�0ʎ�xWzp Ѷ�ݩf�+Bc�.mL1Ez�#̡յ�xnU�o�Tz�ln�^��z����.u��v��Ô�y*�w3�=��5u#�͇�0��a�����	r��X�EP�7��4�S9�U;�dݧ,�,��n�WȵwOE�T�\2Дzĝ� w��_B���+bvy�/מ�����i_�V3���9�lQ�\�/n4@bM�Ziٮ(���ӎ���l錸�ދT����C���~�B^�AK�H�؁�x��P������^���A�]O͢�9T�0We��h�H&�<�8�X޳ WCJ��u�_���P�@|_�eO<�G��X�Gp��j�]�G:�����`�y�������ȝ����.���9m��8�}nʹ����z�f*/��#e#�rT�	;��_ᡫ�D�M��~���B8��?��5���p�V~��)�ӻwEYܕ�9a�~�x�n>��篧ޯ��妴-��֯�Sd
�kiU.w�PK	�]�}�]>-�p��<DW�����db�&�ڒlK�hf���D7�O��?ف<ǟ{a�B�.�*,�1��|�<�gR<��X�Dw��jݦ�=��r�E�#<�{���@A���x�&:��C��x�k���*7���{E�iX��Q��r���G������o�#�h���hlT�-U��{� �(z�\eq�H���k>f��?��j��"���c2(N�/g�3�!0�נ[���Ƶ�&wE���p����r��������{ �s^�<g0�0�*;<�1Ve&R+7N�KG��{v��`�Y�֥�^e~����������U��e��W�a���$��^Z-�9b�A���Ú��geAiL�����4Sb6�we�3���_k�;���-�$����]�:�òq�ۯ��$���o=��R�7n<6�C�>v�-O��i�{ Os80����{��Ľ����@�j`��dW���[��As��_?��.���H�w�a�^&�,*Ӯw\ټJǭ君���)w��w�am4bi^jmuٺR�g B�)�"�"���T�����i�/:	e|�����gU=aE���}n�Ý�C�Y�tb�<��JW+m�]n�՛��c�������NW�@�fݪ�oķPw�m�9���YC��Ɯ���ǿY�\R�U���M��U�yz�R!�����ݟ-��_ZO?z��w��IO��fKN�=g״�rP�"���:�ⱆ�����Oͳ��F5�-�����&ر i"�K,���w(�Sq�)p@�;/�G>yY�������Z$uY�b��R�ŰZ��޳�n#X����+��:e�/��-���� ��+�,�c�w�5� ������;I�b�.Y���o�)�2V@ǿ>|F �~X���/ ������읟�����E�5M�	(-xS(dHKk2	X���ee)HP��i��])\���e�]O��VHF	�\P<g����Y]i���n���;֍=�t
Z�X�������#�	���W>E�G�W���2GE��/�\�2v��/㶔�>�c�OlMH�J�-Azu�l�1�F����k�^��pC��4T�J�[.��c[�c�ߣ�j�@���(�в<�j6��!W�&�����|�����W��zY�F�ʚ�F/(u��G%A}��%��ٲ��T��X�W�n3fl�A��V~]��|��\�@{�ym���|��:�v�U�r@�#��6�
v��16 ��<0������y��)G�o^_g|M8���{��@�T����^�N�^�Q2��j7ID4g���I�5�e�6�>I.���0%a�:�M�Ր���~��� �	Q�M<��!x� ���h��u��Ɖ0���i�(�U��p�J�|(J�]��ׁ�]�L]6�Dyٵ�����~��]����`z�S\�=1""�bK��QvEE��%��x�����ͯ�ӣ\���oV�6~U��y�����|�{���ry�3���'�R//`S���^�{vK����ۉ�{ܿo�Ym��|r��������jZ����P&XЁ�D��}C�Z���NoF$ӟ�<��Iw
��T��c��^�]�+s���p�Y�~����s|�#k�A0��I.E8^�<w0�t(J�(��0f��JA���;�k�KV����Px ��(��;ʮ���Kf�����|b��N�/j���roZa^�-�"5���^�OE�(X����dG:K'�(��pZ����֮��Ɯ&��|�B�y_ky�%�s�j��5����H�I�}(61\\���f��24l�7��ml�T0�_��-���kϏ�U<{O���e(�����]_B�����uL
����|�`�+���t�j���G2��	 �aQ� �0�M�#��%��������k�F3��/�H�zu���^��"��ЯG���G����J��(wϻQn�ѽ�u�������)�8����׮u�5��Th,|�M���1�t���`�Q�A��}���!��8���@�3��G���U#�u��
9U�ƣC)/u洚A� e�����@6;(sz�@�f���Q�2	�@RW�h༃�;�sU�����Λr8�Jl��/�?|G�&��J��n�����t�Gv�a�l,}9�3�Ǘ�vr���_�������7���w�vΉ4x���Q�$��տ"ǻ����r�!����|_~�w��w.~����ß��>|��H!�S����	�k�CPC�#7�e5A�7�k�xc�Nw�=��Y�l�ia}Iئvj������
EA{�@]<��K��Of��~���7 �&W�F�ҶP*6��9�����@��(�����;��ϏT�;@��%ɑ)t�Y�XD=����xG3�3�b/J=�1@ɸ��(�VTeƼ(<*�1� c[��B[�d\�
�t|Ey��cic��@�b,(*�8�T�V�<u��aC��������_�9���>m���B��(%�2(�����#�zܰ��Oh�{�k��cUVַhƗP�[��i�/��}����6�'%sx�QwH��[�u����)����Yk����W��ο�_-�bD�ƙ�%�g�_����&D�D�*��9�S��g�0�������K����_���E�0ʳ�~��fS��*W���u-�Bv�o��90!�y�V�}�����'�TY𖵁e@9	0HW#z��ޒ�#Q��ma���f^�T:Aw����Av��F9 'Hڲu@�JC�Q��L�x��]��'���e��7 ���\�SJj5��jm� Wp��,�Ψ���#��b�5
#��li� ���Q��'��7�]���d��e�$��r��xqGE���t��G����FU�Jy���LGd��pE|���~��?���ez�O����cw~�������3ǻ?F�������o,O��}�ˤ?	�������������K�:��ѿ6_>��r�����,��2��B�����(��#C�z�B����.d]�>_��Fl�΅�Y{o�;(�����`ĬV��֖�6��j�Y�͆ͧr��V_7��jt��w>z�t�|�m���P`�V����0T�r�e<�1���/x�j��ɱh���:'-J��<� ژef�|����>�G���ͥ��Aٟ��6Z��A��$�X7�_S�p�V���"S4���깣.tz����<&�����N�p`e�)��z[�|���{p6���<�����Buؙ2���T�����QO>�,h���&"��'2���	ePF5����gZ	Q 8�y�T�=���k	�	����h��B����~�`+�%i����L�ԑ�Ӵ���v����a������������o%|�=	o��^Fxxz�AF8�i�ծ'{�ޒ�S�6ɪrO��&�<qk8�X5�4w��֛����;�:��:��g�M��L
r+z*`o��ͤ����7I�v�ow����Jf�s���� #��a���SLf+�|!4�R�mQ{��U��){РZ}��*�C�s���a	�N��\k�=��(�E#?��rw�A��� 5�+Y�"�(-�bmR���̓M�{�<��k包�s����z���ȍ�����W� 	�X�n����7����������o��Q��Kx���3?.�w��zz��/������E����1�zJ���^}�����b��_^�_�L�~(i�uU�����)�\�0{2�sS�J��)i�o0�S��k������^�M�3f��2��,����]��Y��j�XRi��f�<�`���E�F�Y� f�H٨�q�� w���$��@�X�z���+n(�u_'%��%B�k���|*��*��H�v �����S`�:h-��� �b�6!p�،7D�`D'�i�]���N8�����N;�&'J�"㜨�I�h�6ʺ�TA�%�".4G�ܽ�����}U'O��(�$w���RKn�S̐c.�6Y`?tr� S�y�>�^�b&�x�	��\��\A\���U//(�M�?�� ����s���&�B���f����^W�c7��-a#�
�V�x�5����=H�'�2k�hDyІ�@�Q����[�3��B��p����hshƇ�_h��o�����'?2p>n�N�j��ޠ�#Z���j��dЎ�����o��d�\���2C�l�F��|]ƭ(��q�^aZ�*�s�>C�"�F1��tb4c5cdD
o��l����rN:��#Д����0p�*���)s���aΡ�9��K�b.z���i6�mvc�@p�ph0�|
�Z���&�e�@���J6��=�]��3���1���^��P�U�yv^<R�Z���h5��q �^�kz�'ְ~+��������Ç�����c<��7��.�Yb��e��\߭���^NOO�qH��,oW,��D��JT�U�B�8W��JD�є�hyg�vӺI\��B��J�6*xcguk�d��,��J�7҉꥛'�JK���o+ָ���Nݕ�e�m�l9x&��WE�vޠ�������M��P��=��_�sQ������l �@iڒ�J7�/. ���w)��t9��z�R'q"�@��:� �̆���\b���0��m*�QK��8�k�`"ܰ�$��? ��aEe_5E�C�჆�%���1�"F*C��{܊?C���B/F�Ս��q��s�xkY�D��╧����6H�A~��4[F�?�x� d��HE����?x��y{y�yA���h��Z�����~�=�E�Z�pg�D~D	>�8�}��lmO3�(����%�:G:f�Ww���YY9�G��Ywo��.�E2�K�����@pl�a���<e��Sj���؅��O��kn��κ�9���E��^�6����zѡ���F�2(��30

JvFU�Y�~��B���ܠ���d8�S����Ho����B������T��a�g��7��N���̢eFW�!�2�.��"Vn��R#�ڼ�;M�e��˼�^��3�k;���׌��Z횃��#�H
j�qR?�K��̈]��p��;�u�#N�Aκ*jȽ�_nijX���^�Œ粀�?����,�{w|�_��W��K����o�P&�nW��8�e~?~��0�{w�æ���7��&Xsò��Ր�W�#N�-�.�Ym��o<��+��m���t��z���!��O�X��W�UB������h���ϩ���\-��_b2/]|��í-C�n,����W��w����W�v���P��sD��&4v.4�������X�����^	9��bw��?��r+���A�T����k�"(�E�� �a���F
���cK7A�\ط��G�M�;�"���t���ר��qo���I-x�\L��@���潺���^Wh��@ܫ<u��Aq�,�X��t���Y��}Piy��x����.�]�y��6'����R �W���B�\^𸫡ZݠfH޶��7I�t���<l�zC!7Ӭy�����ׄr6�Bx��i��Iz0����#a�;3������*���*=i5�Cv���bƚg��0���;2�4(�f�u��s�Tai{С�U�(��@Xwz�96�	��p��C�l�.K8�f`k��/�_�����W��ْ�)�x'/����t���8 pV�夥���;**�ʜ�0n�FUi��}4åS U�6��
�ZD���ٕWVO��1j8z�^8�/h����ɼ��O�欶�:����c$�Jb=�����!zS�t�I�l{�y�?���� �G.�a;r�����$A<�n�C3��N�ةde��:�Hw��`�����ͿYd�����ey�_N��<}�5ٽjy�1_�O% ����b�}��_�����|�����vd�P���G��X��f��h8!�����n�m�	d�w�j�I�-#nl�B	.�sd^kf�C�D#!w�aRe�,�b�b�?�!9�a��1�6���S+��.=�nl�f�TO��C��+0I�
�<�FI�h�K}��+�B8�X��R,עG�j��J�p���V��{� ����?�.��yf��$�)�;B�#����
*ǫ�㡚���k��-q����͑-Z���"wAv�9�l�Rjq�j8 �ʜ�*^ h��fDqj�ddC�M�	��?���LP�n���Z��	x�����4���TҰ�z�D�fF��e"o��!��}�E��[w#�H&���uvZ�;���u���˕D��A�{9̛r�q|�y�;�W�7�y7q�[p��1�
�P�F}��0��憊ԥ�	���TƦ(��Pq w��5]N���Za�@����'�>�8��K	�*>�*������%kŬC��
a{&70k�q���p��,-]�m]��*���G��"Ζz0#2�yp����� *P���}"�YPB�n5��3����Q)�I;�r���)΋�����2��X�h��j�RW`[�F]Ng�=�d\��Ԩ�<:\�i4��H�Ȍ�[��`qs��	�R�m����
 ��e��F���e�,C����m|e!������fBS�`|d)�j�;k�8$u�$
��R��k��7D[&Ϟ?�LsFkHD}5:�&1�3k�K 8���g��g�����H���S3��,�拲��鼻�}�l�m����U���!��_�K�]���˸N_r�W���EeMO����d���伝γ.w�hO�pe5p�{_m+�{g��C]���6�79��Mx�ˬ��[�+��5�g�{)*1��P�@ќ�#3�.e�3��Z�֬��^T���{C���vv�\=�g�K*|�N�{-��Z�
�s�k����X^/
�28.x��lp���9��a�����bq�z�j��5�I��Z(ڽ�Uw��V9�:Ҕ��\���R58"m\k^��`�	���x�a��1Rټ�D���H ��頣���'��t��{x�QK���+S�k��=�1D���ܤo�4u�0�,{;�A�s(FJ�*�3Il�{�U�^����ж�K��c�O����F�˖��"K~�~m��:=�J����X`�i�d�� ���׳�X8Y-�X#.`B�関p���	4��K�?烬��A��3dނLF��-�P�O�u�s�;���-�"-7C񩣗o�xĔY_� �{n7/^���\���/��K��R��` d%�B�G3�c7��Xj EO���Z�b@�y1,&x�Eֳ��jT�Ҝ��2'�E��4ן�>�zյk[݇Nڢ���,��f�mx���|J+2Lm�G���cr��1jU���eF�y^x�+��"����l����]��~_�5�-%%'̘��J~�٢7�����ڵ�8}�ݘ���/��B��e�v�_,��/��t<��Ӕ����G�Я7�����ӍW�勁 ��b��Y���CUw�A�
]������f�5G�7���T!�usl�)s������7���H��,�����묗����Vt��x� >v�F��v���ϴ��ȊBNū�3s�$��!�0�arS!�[6-�o*�3-t|�aa���f�żj�!0co���	I9�~�Z�fz>l�������
�-{�o���]�E���@V�VU�/��5�l�R�.���8E�ࡺ��z�NAE�ymC������i�2Ӓ>�LG[��:��M,I��iTH4� C	��\�j��<�:c!�����n'��I��GcV���TI��](�5�T�F��-W�^T�P�R\�@�X��M0xN5��k�^)l�R�"�;�S�t� ����+J����e\��I+�ɈA�]�^ۚ/E�.\�2�|Y�I<<H��R����JP�"��t���/5�����9Ϲʯ�7M������;�=�a3HhU��0T�orHr��N�rrh�W�o�ߒ�z�����e��@��vy������Ϣ��e���AT�]Ǌ�մ)��ޒ�0e� O���҃��ү���j��L����X�f�Væ�5צ]eJ�� ����ݞ0B+`����l�25<?�F1U�N!�wa��c(�2n������*�o���&g�Ôٚcjs�Ϸꊬ�<d��p���Y�_��Af�0��N������(��?���!��5��z��@��}ݓ�_.�~x%��t���H�g�s�Y"�<#n�κj�\��j��Z}Zk�y���ÿ���s_�b����b�Hj����p:�a�[����b��l�+]�|7m�Iܣϝww n�$6���Þ1�.�_{\P]P炞j�,����}�
�j�-�= ���"~HT1cf&x�˩x�g�ۓ�,� ���_�lQ�FMT�(�������4Dsa�)�f�;f�R����U)ЋAsj����٪$�Z��Pj�ˌ9_5�5���U�5Pb�^����[�LYU���;�ژ�7ڔ�-3He((��S���|\��zb��z���j,rL��H�c�e�>�fr�{�.r��|I��5�5��r�H[�Y�����f��8��FSp����;����`G��QK�`
0m2g��!ܑ0FZ�;��OD$���`|���aZ=��dB�8�����Sj��������ӕ�2U��Y��ۜiV�R4�w�F;��hF��ٔ�a%˥v�\�eK �^KKP���)��A��r��(��#�qnTc
f�	���:q\w�}U(|�S�e^�G�
�_k��t~z���|v�]Ĕ[�*4��N��Q��$w���=4�&]5���'���9+(5ƀtƃ���(mV�/j��?Z�T����DC,Z«F�쾴[�r�h=�b���2��A�����^,ؼ<i��Ų{�|�?��b ������/RH������rxuW�O��p�6X���n0o&�J9h�`4��6ܢ�;�E�T����$7�i�z�b�s��C����d�~ּY�YoQ��;���� η ��>�ռ�zn���_��$�%�Nj�lY�`���(�q����ղ���ٰ6�8]�����_ɫ�D�k<���<�u=ɮ̻#�;�6�A]����q<)S�7�q��`�W{>�<�^_]�b���F��9.�[�S���kٻW)󟗵4���j�\�,�5���ê����Sÿxл�!Q����Q��a#v#W<��<��,ݲ�0�ؙ�z�ȓ"����F8*VܰA�f,K������ �^k�PG��j�V���Z��k�~�)��G�p��h���H/d�AO��ֻ@��Þ�º&����j�!_8	j(�t(+�)_��>�$���`�,{K��^�>-����y�����)�l�@�*n<t��k�p���w��\W4�{�;jgyoW��N��bH|��f�>(�J��#E(t'a-�{��x���c�̇2�����2�߳�C�=��_�8�\.EV\�ф(�x��[h#խ�>�A�s����^gk P��#Qcx,�O�14J��I�����:C�FK}�hA2'�S�T��,JlFͨ|�]���T�����/��Y������6*:fz��y���>�(�N����r�2;�7�C���d��Ǹ��dr��d:�dBn� ��-H?4>�
ָ�k�]�݄�{в�T,d�5�ja�P����^�:k�-�TE{��u5x{V�f�J����[E�pc@����/yX���zo!KO������wEi(���c�2(����/:_���e�����<�X>��7��}���?��˗r����H��x�[k/rL-��FmF�]x+3CX\��BL6�5��C0�}�J�j�n�[�U�Ì��E��\��z��/j�2�s�2!�˓�	6���  ��(�	�rMG��쵁�iJu� 2�({������LN�'|�!�J!�0k��܋��M]�zO���-B��^,���H*Ą���hB1�wW���~�t��=n'Dhj��H��ܯ�e�~P�c��!�ދ�P /�׈�l�j����TJ(�J�{Y���ԕ��h�l0�H	���F��8YjE�EANq^ߌ�'����?���d#Ϝ��	����u���[�n��O���uͲ���酘�x�^��T��h��S��H_15�ߧ��O_�r~'+�9�1��YRԸ�M�/�{+i�[���S�mܺ�Q���a��"Ug�v��ji����1K�{��C��T�u��'�*I;?�"�CB6��+t�1�^�@�0����Π�"�:�W*T\��%�2~Wˊ���S�6E�
�F3<E��e���;a2� �f����b�9M��ray*�x�{F��#�t�-�+��_2�u��W�fZ�8�?�2W��� �]U��Ԉ	��������A=�Z��r������O��lR���Dj�X��^6�q��u%�߫�s+�ţ��f����G#���_Ex�7�y�B�zF��F���l�f��`��V���
S�e|1��ꗴ�T�M^C.�@�`M��t�K:˵x�;z�څ	`%ҷ��l�_W�k`��0�+�D��Us5��ZUw���ɐ�bv��5̮�E�tRj3_I%\9�E�!+�y�Y�A�Ϻpԇ/:�Oҁd�m�'���%m0Z���9;Qs�S9�u���	�cC����|-�P���,ic�-#|�;`Q�����͍d�Q�5���D�N�g| �}���T�\�����%�^�E�o����S�A�US�̎a-�IM�hx���=�f
 9�.RG��|���LX��yR��e��	�Zd��9�e����<��K��)��,�B���d�Ժjz �fT����x��OGvΆ|s=Ίh
m>��I*7��܊���^$�B1��ӏ�B/��I��;&�~��>X�ԓ������si��s/��m�#�{UIg���4�<�5��q�5:��W��D7R�F�S��⍲D��B44+��:_�5������ƃ;�v�xR�ol|�ը��!�ֵ�K�(���U_��)�Ք���$�������1���[�q��:f��&^�o��e\���ڴ,6��Yǔ�K86d�7h^���YrUug��EZYWP+?c�&��'�jq���6�D-:��m���s��DVj'�mj�����m"�-M�D5�j��;@�7P}�O��n�v�7��(Fs�s�4q8�p�Ѯ��9��L��;pYhZy���4/^>�T�2��M�ZԣKy�۵Eu�1R�g֍5�Bnat��l�'"r�F����K��^�ΤOP�%=D���׉��m�l��mfX�sX6�Z��zs��9\�/��Bw4�S�s��Ra�Z�3���2(P�Q��շbp��]�EC�;4	v��Rk�1�E=v������H�k�>E=�$-�Y�Y�=t�Udu�ʗ:b;�ڣ��x�Rt9�Z����cɏ�� �O�殏�-{�@yG�R� �[�rH��2%b�kxD������qB|��U��%w{_�
�4:Ae�-:j�����U����0D�QC�.�U�j6Fd�ޡ�/�+%ș�[���H(Q?�T���1ƫM�c\�%=���jy�{� o�-G���ʉ��D������x���Te*t���*V���б��l��u�>��1����K�������+]ĕK���,5luJ]��T�k��D}3��1�!-4X�{�Zme�N����Q����~�y�P�����\qЛ:���a{S[�f�����)3x�9I�b�Cgr�#�pP��8	qG �A�%��dT3I1p	�v�Qe�=���bI�GQO&���^ƽ2�h��);Z�^��� �$����e�ު��o�+sg���i9fiHy�4�'�����Ud�1r�-�;��>�	�g��9�]k�]�)6O?�S f{�+�>�_8�4� B�)*�o͚'�.B��a�'�ZiT����kFY�P"�l^�������Z�w>�{h.�]_�sQR��v��M��`����s�G�~�U>6$�2GG-��$H*�n�O��j���rϹy��[d�om�U�W��e*[�4���#䦠0�Z�_�˜����h��O4�P�^���y���e�x���T�Us���g�u:X����n��u�y"������lF���ڢ3��{&U��KD�P���F�0��j�v��,�*�I������bYҵD�\�8��W� .����x�.2�B��K�'-=Pm~�+a�c���N�8nkIjtI�8��=��"iN��yP�i�����|4�1�M�w�W^���Tʀj\+��2��!<E�W��,�>(ۜ5�5��|��ӓuTZ�L�uVC� ��'�2!Xʴ�u}9��۷��o�][��H���t�xj�J�5�orP�����~H��y����������J[�	t���9�����T螇�]֠!��Lup�"��b���`����9K#4[�@*��`Z��Z�c��1���w�t�if�&.���ھ��4���	>[��֐OX�D9ٞh^�vÈx,.����-��{�m/��K(t ������ÑN!l'����$�K�e�����_oy�f����E���u�,�r�,�|fDdUJ&��&�8�Z~�� [nz� Թ�3�c_����{�ˇ���]�-o.��4!�~P�=�U�h�og�XH3%��Q��HqF����7c��{T:���һ7�a��а:Wm.�3�T<�� �������/J�м(��uR�
Q�{4����= �g��%3�@PT\�W��8�d��F�qԖ�=p��2��j=����d��+����[��{��ކYuL�+��
G-�A;߻�.ʚ�S�P�>� %H��A�������1��ԹGid@��9��-E�C��(��o��<�/y��(���Y+]X6������TCY��q�A2V��bڿ��]�j'5
��fP�Z{��[����Z��+����j���a��.ZX�5���an���z9�8�}�5���|p�b_��A}:�Gft�5�:Q['�)��c�Ot�MQ�x(t���5��3k�n�B�^�����4��7Mf��
dd̖re��3�U��;uF���S�7 u�4���wv jߝ=��u[7Ր��Em���X��j�:���L��i7��N�3xogL�*����, Ve�̄5U+�X>1��Ͳ	ղ�&p�y�=��ج�ؽ)�d�bo¯�-;#�sM����oW�z{!:)!wO����J�S
]ﱻyq#�3���o��S���N�u�j�QsE�����Dm4��|[���TVS�k]��pV0�\X���/ ��2�ҟ�����O�G.�����ox�����ɭ��Ɖy�®�\���B�h��y��Us��B�����љҎN"�=���l2�+�vQ�1޼��@���I�hHvd��a�SK��������nH�%;����Y�:�Y�ͨm��V�����O��u��$��/:T�\'/� pѽ��@Kւ�!^�!���ѭ��� �8_����MQiL-�I5��'�,'�����F#=&rVG���޲{��>zy[�3�O�p_{o����)�*�BS��2Ou��=�Z$�ys��>sтqT�cP�~9�.�������|6�G���{y����vd&�Z�tU�;�ᄓy�����F���(5���������{�7U9^���9>�h;R�J�D�����S�!v c����GH����W[��h���-f2�uh��K��/lݔǮ�a�����t��M��%*k�����X$:�,	Z~�����������4%��A��?qD�兼!�ߴ�+���ArM�6ewd�5o� @�e�?�k����u��n�u�&��1ED�mg����ք�ǎO��)���\��V�􎓆m��Z4����»�}�>[��� H��Fp��.Ys�:��	AX��H���9'5�ZAdN��p;���\}��u2��4�:�`�*`-nV�N�kf{�ME�k��ec���.�W-d�ls��>��\H�JO*4��Ž�' �,���;t�4(���,2b$E��dB�Ě��|ءMk��!�u-��Z�?|M4�����s�o�"*D� /C=깷X;���-KW�z����ޅ��bWe�J���3�m00	[U�.��+y���~u������b(ܽ"�BXic�F��O����@��1�8t/�M�on���C��\����h����ޜں�{��ޔ��1���UDIt���ǫ(��b�u���):�_/W9O�XT�|���������P@a���[��c����ɯS�ٍ��1k`����椦�����"�	���|�n�<p:��dS�jWx�7|q|t��'�<�փ�+MK��������p�%Ǫ�=�Ө�?&���tG.�9�b��:�t�rOM��T�����b�FPY��B��e�P�;�<����5��rR��$+uj)$�7�M���ɸ�T�5?%n��{����Yn��d�mYN���o�u-��,�q���@�k��I��j���b���d��5��i�
2 �Cq��`�,e�f#Fl��� Osy�Z�n"�.�թ������7�W��7를��`t���6���NĐ��Z�ǋ��S�P!^T@w�첵�$��)�K��t�vmv���s�C�u�:�ʎu�L�X��yV�e*m4�*����U��!�O�?�yN�7�ej�Lq��&��#����x��qhy�m(>Kjv��ﯼY�7k�ז�:N��9�u�Ϫ0�s�8��(%?�¨Mfg:5&�5�����؃g�Δ	�8h�U�+K����hS
��cq͐�0ߤ*nU�ye�BW���D�f.t웧�&�z�=B�wl�	��@������.܌�.�Շq��ȸQ��\�yY�3x��c�s��B�tr���i*��|�ӗ_J.?������#�]#{+^�ݣ*Tx��v5t�����<�͑�_|�Zt�sp�$�x�7o�U+���Q�s�fD��إ�q�'=�g�q�̽dN��E'����Lu�J��5��l��|Tm~�^$�q���t�ь��YBL��1A����o��.�r}z����s���ւzk��<n���1�������&T�Z[բ�������gC
�pb�u�s���iH��s�m�N�Я�Թ;���䣇O[�yօ���BK��?zv�hc��)[��>9�cQ�.U�^�'�f�u��:@P"o~�>3DO�T���� HaR��*>���A���Q��	���z��d�P�ZZ��^��H�bV O��k��S֒W�L��>6����`
ٵU�� �X�	.�k���T����D��@Y�H��s�S�gۯYs�@�/��uT��}�o�2[<��h��^�	��c+���E�!���-g��x���Bl{D^<����3H=O�)�A��).v&-c%���S���Y�8_AJ�P��!�>�.Zb
Q):��WOO��){K�V-QL.���SJݘl�����g.��q�ѧ�i��-#K���[:��L=E�e���v'P�Kf�K/Yˠ��9o�����F[��lNZƷNgF㰗�W��1D0�2�^)��O���"��x$�/OOdSŜX��л�]s��alo�^���؅~MuQ��}�f�\����a�x�4S�����Y�7j`[�����1���`kC/'��7'��B5���P��?��C����d\V��Z6-�#T%wZ���:��Е`6�ࣩ�c�ܢʧ	:(��$�|-F%B=g9��i��~�xSɄdp�!6!Ѽ�ҾT��/�`��!�=㩛�I^�Zۘޜ�n��p�M�&�:�F�J�dl �`�V�<yp�g��6��ã��}������n*�ȸ����V0e���	9��+����}�e_��+zI�*�Es��*�Ȗ�'6���NP��8/sA�q�.Ve���'礬M�se�^��jW/�}�.�a��:˪�W_T�F���.Q���5`sXC~m�5�csB�.G�i�K��tm-?W۰�jȬ�w���0`�T�sE) b ~�ݛ�L��6��!��fy��$)BXؕ�ꛒ�j��J5Y�k�)�X݆@�OlB�a}�ƨ��F�Q݆�v��s�Bq��wķ�r/�e�O|_NE��"�V��e4�����k���@���l\�B����YEpk>1�=g/uꗈ�닥�1�C�76��e~�QŮH��F��y����vņy-��r�F,(��XΤLV$�������|jb��"�o-���ZU�'��YB9����;�o�;��9?��L�H4��e�����\�����d�Ie=���yk��2jȇ����\/�H����q������j��>W�Q��J�}��j�;cb�r3���9�UYVI5:C��U��6�^��;��Jι!��Sg�(�Zw����ӥ?a��V���^�V�H�"�a�`����R�&\�ʈ�sq_�g�Q(��	�TF(t�8��Ud�z�]TZ�ƌd��x��F��M�ӻ��EK�Ue��=�mq���t�=����{��S��C�i����5Ёoܺk�h�Xd��8���">���٨�"c�˥�+j�͆A3�(�e�,eU�d5|��mDb�D6n��	�Us��J�C�0{NT	�1c`���A��=dޕ.�X�"��3u��Ϳ��0up+���i��l@6����k2wF*
,?J"���b���F{4쌶��ߕ�q�#��7
�f7{@�v���zdqnJ�[��������r�T_˭�OoU�**����`�&�TЈET���=m��5f�J���Ns�'�aqlJ�[��f4��k�zn}4��ހ7{��ą�&B�c���W%����hBY��A����^�t�̧"S�.�r(�X�A,DB�l�>ur�NV�J��RP��|.�j��"����͞�3�g��z!qr����k�����;��? �}��]��:�w�K����}���G����B�n4��W�i��ϛG5����S`&V��й��c��&��YGH��a3�ӎM�d3��V`�<�k+(�w���b6jZ�_HC��;zd�`�F������:�9��kx��e�\߈R�9�' �4x�B�5��ቻ��=Z�=9����s�����t���s�P}�ze�^�NG���~{�\���=�ݤy���_c�p$C��m������<��,r9'|R6$ ����n��d���m��R]-̥u�qc/������|�ڂ�\�y��m̭���Bwo��G���6v/�7���Q���T�,����H��#�U����(�~@/o�%�JAp��,����J��}��C����<�~GR�f/_�O���j%Gv����L�?��-���V���=�����/|���&�������N?����6˯�6���Ssw6�*'+u3*MOC��<�>T�J�����u7�>ro�w��Y?����.g4���)���#Zs�����._���\�/ܘ_�aKm~~{M����u(�y^h� ��B��f�@�����'t�f@!R� ���q��}�B�`Z�k J���O^2���P������J���s��Moϫ�j���jx��KV���[��,f!��}_�D<��/�/g�>q]��C��i획�0l��#Z��E6",���6�QJ쵞,�JE�2�)fӬ�ͤg<��(�l�9j�=��?>���s^ܟőϣ囌|$/��P����IjzU�a�5�7�_'����Q����0|��7��	�ȿ�������]����E���K�D�د��@♋��N �q�snJeET.F���o�Z��DJ�hD�TV��w	�AS�h�{�aC|��7�\O�m!JEs�u����e�q�yގe#q�Ǻ���戊|U�R�����.֒4g C�c�qI����1�^^Gg�W{��wk���ft�<S��~b�ޚ�'
j/I��9�����^Z��k��Y���sG���܌�d�
��IN������+�w`�u]�� ���y2�l���W3��Iޘ�U��d }�=�����V`h�E�Qۛ�J�`�t���C9_��LG�f�"OW���漸�S�,����k������ X�q
�d����E��	�LO��q5,��)����s� =�����W��I�q�ˌ~�De^�q�(l��d����V���\��mc��f��jP�h�D������T�������m�}Иs��9�}����q�Ĥ	�*��"Tj�����_��T(�*�TI�6UUTR����
A!iS�$�$`'q�q|�N��{�}��{�9Y��c̵�>�~�{Ϸ_�1�c��c�>/�1t�B�q�u�=�]x�Ơ_"X�Ew�f�g-#(Icǚ(�j�B�D��c�'��Tv���O�b�9쵵!GAc�b"���u4�����%#��Q\-�B�y����4L.ׅO7��^�
�B;��w�.��+c�M��������1�tḖ��(4����h���'-wt3���F$7��I�#�-�HL�fF�N?5]ł���7[j�T�0��#� � r��q��e���ۢQ�Y3�&�33������y1K1;����Ɣ��\6#� U�[C��T��HQ�@����\w;n��趚Y�r�ɯ���ū1�{g�I��6�u���J?8�]x�}�\ô�]�馝W��YQ��>�f��YX�<�YE�dAZ�k�:��d|�+%�{O�U>������J��,~���ٽ4�a|��>.&ĵ<*�����\��X�2�-��e��51��v�����+�na'1�?]P�H������ح ��N!���Q�s�`�I{�}�X�[�Z��t��3�b��d>�q�>_[��T�[�F��?��5�����/ҭ��ug\Q׮���
NâpW���h�Z��Y6�@I�퓺�80�lq|��\p�i�
�#J�դ�g�h\+��Y���!����mĚ�N���IK s��u��}�Ќ�%�
��ڔP?HEYj-Z�Brs��%�V�n2s��e�_����Q��h ���V�]�6�%e7���� CFٓF���iY�I*�OU�	��
j_�����"`Ò�{*1�=������]�9d|�nbT���h�p�#�i�&�x�c�X����?���0���ŝ_�ĹK����<G*8un�Q��s�}�Y�/ִF�n�axO��vX�;�փ��tӻ�7J���CȠ)Ow��ΩT�5؄08�Yc�۰:��{�A�����fD_�i��2v��U��0�6ޙE~�n�Z'Ԉ�o��7�����`��( #�=��q1Â�|��<�4�[l
{Ũ+5#�}x�X����qL���}qa4Ɓ_\֕�ĭ~rGJ��&��V'.�49���r3 ��v;y�,Ϝ�Z��޵�]ځ̜a69윀7�˝F|��4B_`"n�V�9#�tC�@�[~o���z �����i�=`^G|������\QK�P�CI�*����Q�f��]8�8����j]���^+����!u������%����V�(��r�0�E�0�i�b*��[K���63j��Z�����f�q�dj���#�)ƓX�3���������:7���R6p��G�(�NC��wT��R�u'�Q]L�3Ўj�ڔ��]�^&�ɻ���{�~��ǫ�ۈ���Ns4׉��lD��q��_"��T�j�\���#�������ALk�����Ê
,��̚�!#�2ݎ�W�\ڵhz*`�U�%d���?# ��E�kc0�⸎��ÞfC1�-�H�ܥĈ��.񹷑0��-��dk����]�/��8L�v�<f�=^�\�u}`+�hȃ V����0Q��%
�f�������X^�����܉�ee�|N���z�\d��܂i������V*e��a��|���.w�P4c��ֽ��Uq���l�g�c_m��7���:�=+7[U[\.N+���`����e��V3���͵��AƁf� �@��=��f�p)�2���iܮx���"��Ê�qL=!�X+�3�ft'L�yh*̊�Ϻܝ�G�;	}�cZ�Nk��D� `$@�q��H����q������S���h/}g�W�ݥY$�	�ȿ��Ђic�J3�5 =-�c�Y,W��3L��-������	�f	1+���
XpM���G�o2$�j�|���K%/�k�3(�|�Z�emC{�t46��2���@��׋��_���Y�pQ�ެp���"h�V#`��Ͻ�5bs������(��	�T��F�.�R��@�2<-��<H����=��ʝ y�)&_�ۆ��ݢ�v�ia�YG���o�ڣz!�+wf�e�\�ئ�][ϔ��Ev�4����{�J]P����v���FVO� ~u?$��Rv�ýy��Za��+A��"� bgA�Ҁ�"��royN�ֶE�qYd��#����GAP�JŘ�B�`!2�K���[LZ�a
>����lx�k��ժ��a�~�լ�E=��f����ƥ��L����x�gQT@����n���'� B�!qP�����4�b��� ���S;H�	��him]#.0#�Z&��юu]���ȭQ-�<X����s�>�g�5�� p��fm��0�e:mIr�	�|,���ik��f8h����s	ymqP� V�R�	eM;J��Yk}D�j�a�Ә5�3�86R��3f�=Sk:�섶혠�n"�͓.�D� �����4�B����U�g9]�ok�`/a�f�=6*^i@���Z�b$�"4%H.���NӏM��g��+��P_�9��^(��&J�T�KP%2����s�Կ�����t˛YS}L�Ե;�ۈ2���e����pÐ�t�$uD��NQ���`uŀ�[w=7482���ژ!LfZO@�"�~$Iw�}�Ih����#N�-ޠ�4`���@��bܪ���Uo�f��T-��Y �;���������y�Ǜq1����kh�Y�V
@���,�&[�J�5�Xs�6�y�LȜ�%+{ttjD��>�l�v��G
G�񩠐��|>QUP�܈�(��X�,'q�; ,(]�K	)�̤� �8�.i��pz*|����!�k����œ�j.Y����N�>,����j��1q��x6A�n�r��i�wgb�a�� ��oT�U�����z$���l��8nIﵮω�n�<��}8ϊY���Mg�����q�Mx"2�wD�Ϳ;�i���,^�.pW��NR;�$���Z����I|Cާ���#R%t�@sf��%?H�<�E$������ :u�h��n)Hޯ�н�_w�,��"ť�\��{7��4 �u3����i��d��:�g���ɭ͹Y�/n���� pz���'�o�^�ƚ�BaU�sg?�����n�h���'�6�ӳ�Q���Y�+|�X�`����_Z4Ff�m�*��7�j�#r��q ����w�`k���Q!H�,v�I�aM��f�XZ!k�c~t�Wj��e��j��
��]��ʧ��`��ڄK�O?q$��*�<zw�&V�RE��],͚eh�aA�	=��O�	�#K�k���������z-F�Z�#���|k	O ϠWy��`���k0���7��o��3���y�m�c�f"�r�q斩];�7{��UQډ30RP��������x���Y�Av��2���]Z�oRZ�@�G��rof��ks\>c�K�8=ZǏ��LU�e�µ8W�v�/[.��{��`)�"����t���ުR�����c]���������y� �u�]�:<:�4z>��R`^��p:����b��ʖ�A7��I{kI7Q!D	6^�J6��``�:� ��Wj���y�v͎��>�P*�	mC�j#�<M+_ԿT�!���\sʛ<�S�fĝ�w��%�@!=�<��.T��[Hz��Ͳn{Y;Ig�G��4�M�ϒ�dk�01�R�+� 6!���tuiz��ݏzBր��t���^�'[��1��w��`9�qVeQ�Yc
�����,���,ǿϨ-n��O��2w��dؾ�̹�0u�G��%�$��|�k�
��q�����t�HFk�R"Wz�	�*k�)�bz�����-&]�*!q�m�g5+V7*�J�iׇn�c�L�k}�z�u�F�`aL�k0�.�u�	��x6�^XZ������onT�������T~���E+\��t��b��Z.�ia�Ga�w��o��a{@S�w�]�-Js� �yŗ�����9�������{C�z����.��혩K�Izbh���b}�hq�Vw��P��5c��G��a�����hI�K��K�i��yP;m��LlYT.� @�F��kD�"�P�F�f���nv0���Q¯� !�q`��I�>�a�ȑ�it���������u���&`��_ ���b����|$H#q�o�8� �`U����|����W,]j����q�	�3S:J&:�"��֧!^�!x�y�)\.�Lg��M��߁ ?D %���D51>јM�q��G�F�)����Z����L1O6��0�p�\�+��axI���'��(R	����r����{�wt<�Zh1�	���e���e���h��<�3y�����.���>-��ӻ0b{��0�!�#s{DFg�>0fʖ	��{\��yuL�(,��Θ�2h�S��Z��+�s� ����!ɞ��Ip"�7q��"f\�7P_�iq3���Gm�;K�׳�׻�9rt{o�]v#�����·�Y֒ �-|�/�~���g�^-��[3�O%���F�"�cA '�<�_W�Bꑠ�w8���S#d��vtް»b����� ɿKᙖ�>�];��&���pԤ����E`,��TJu�är�S~��
�6��ถ�ň}au�Ƒ:���hv]|lf<�VR����sN�0��u�Ř���+y�9���L�a����I�R���>"�X�G@f��ū�T7~+A���̠��~��h�04�q6kAIa�֜� ������+ENnù�
���v:gÑ��k��9�l�*.w���H��j;�uS*��^��=����J��	��Q��̆�Q�Y��xp������1u)w*f�es!��Z ���ݵ�)�W�� ���4ֿJms�"����-�k&"�C�R��� ���x�C��z�A`i-}��	�U3�u�y�J8.�u�7��7�(|'q�2u��EF� \�,��Ѫm~Y;�tn����e ��I�ﬡ��j��t��>�ܵ�R1	Z�%@��^�w����J�����f���^�a��nx�E��^��k@�*8�=M�'���}^] �Qg�g+f+�������'wV��TLY����,+�
�P��ӣ.hlV��O��'��"��F��%�yF�D�畡��Q��`\S)D0Fri)�I�=j#�Ј���x�Z���!,�v�;~���	3����Z�&zGzF��:ޖw��i�������R�ŊDHY^�0����
"��1��br?_��!,����Ee��Z�}�x�J�Ɠߒ��.�K�/6{�����A�^JK�+����su;T�����c$��w1����X��� }X�np���� ���~q��D@_}���\lN;� ���I�E��(��{�;Msbߟ�&��-F�9�j!��&��Պ%�>f 9qWᔉ�X�s���M�#bB@G�a1J�]�(����>�� ���8hό8�n��Ҕ��x�6�$;�\��
=�CҴ�b��n����1�gߏ'�ة�w�Ҝ%�� ��2��@Ү�2��i�+ h*��xD�M�NG	��gk޵���PW�q.(��x�.�U;�us�ٳ�k)�E���\4��!����4o���YBd�����2����Z�@��Ҭ�s�֖�m�s��z03
f��в<��6&�Ŵ�6���-j�Z|�u��S(6�1anҶ�I�Ō�C���������t"�됬1/u3��bE�P������ыC��L
�EϚ�k��Na��w�3�� f%!tz��5a��qJiJ�>�&?�Z����`J� ���B��q�K!�u��'�>N�,2��[o�4���L�G�9���m�g���(�16>C��0�?s�0W��ҋ��G�?*KI�uIT&S	e-�,O�7��%
��\w��-�J�`V�G7?�!
��ӄ�C��E�!�=�> �n&r��b4�}"�k����n��V@�}�XP5N���vI�*yOK����������H�ͼۓV�b��^�3x���Ü*x�H���|!O�=�M��s�Ҟ���A��k�^T���,%���d#��W�t���~wRYF���Ýu�d뇔��b>fF?��լ>5���̋E�a}�^�Ҏ���������ʨ��ʄ3>��@�8�\K�����z�|?h�X��N��H?GaJ(l48�:6d^=��s=��	��5h$����e&^sC*�
n�Q"�7K�#W���ERM#���*�g���_����;.����U�pZ�D�X���ղ��,�P�?hZ��|B���@|����	��b�Η�d�	�#���<3w*�+��DM���\Da��m���f��V@��'H�(����3�AtqN��5�~50 �13���c\��Z3h���@q3z�T	�vճD���9,7;�`�V^�1Jܴ���!���hKb����=`N����º:|-"7���[��I'Ɂ֍WA̻�C�;Tfd�M
(ml�h�w�Vl�#����FC{)�o����y�V�o<^K׎b��z,��hu抙��|�6 �[w�h���Pn�e�����Ѿz������b���颦|���O]�*Iv���JѓD�:N����srC>�>_Y�2m�� �8�y�ZA��i�u2�ܕ����$��u��w���&s�Oi��m��6���&�n�_��:�������i�KVә�T�T���~�Q����Y[T֌�ř^C!�0
K�Z��z�R�dVU�X��r'V#$�1���LXXP�X���p.iA�ϲ�;&tu����˖�5h�*IGl��b�{HH���H�ڱ�y����9�:����i;��.U¸j?�j T�Y�b� ƌ��l��7M�C�"'��	Q��ɢh>�dD�9K�f��6	��KB��B�p���+�2s�<p��O�H��!Ee	��^n�KBɈ�ù[�j$d��(R �Z4�j/@�ԗ��V�fl"f>Y�Xh��n�w� !��̓���9�l�g!rZ����tuA�~;]�k��輐k3�ti�5*�ŉ^�]�g�C���tMɓ�SP�M�ݘ����h�L�JD�7AG��t�W!iw�U�%��fL*��H�݆j����a��'F�y��g���r9�k��D]w�YQ�+��gۣ%�1gMٙ��M�rww���z��U8i-�؊a�:e�L����G�kDN� �\�B��  �V�%���t�,�^�"P��O�����:U��r1�s:SU�����[g��')v�4eB��,������k��/�����Q��2�둾�{蹊W��4 �R�"�~X�v�=df�6Բ#��X��j�f8�h��AV�<<Vƅp�����m��A� N�C6u��ꎙ#	����sc�Y�:k�ZjR�gQ���-�h�[�m.���QD�$ؤ�YM�z�d�NXL��WH����_�K�3�̀��ʚ��ֻ�t�f��C�M�mhX�Q�&�s�S�k5�"��\�0�hzE͘RX��gr�*�8J��������C�:���-��!���^'�MՀ_����<��@D�?6/�S�-�6��u�{B����#[m��ќ*�[`�3�Q�^�GlS(�!����,̼r+C�?�_��n3�f����}��8:�AV��<֌��o�9�[+��|�v���Q�+�k��ǯ�d��m&�{�E7�-�;,Iqm�j��M\C�JE�Q08�#��bKp�`(���$�ǵ�ٓ2�������\�Pa��Rm^"����,����#j͢��j�2Ƨ�e��?��6�*,p��q�* 0��~�̼j�k($:�0������:@�-�}	f~���"���P�����g�h���Z�;��"�u�E܌�����ޭ
'Lc�VJ�M��E�L�h��p1���&�`��My�h������-89e���	a�E����_T���T4���1�N)��4����&�����'�m5���+��Ȉ+�8&(C*	�J7[�{���|���K��I(�oG����!���D�v���}SF�+�8BjR����JT̏H�'\L ����[@*6���Q���}M���=��}�N(��T��QNY�`�I^�2a�D�)$��k��]�m- ͥB``�ؙ�s�"�����'?٫H�u��7�{Z6����/q\g�����>�z���n�:�d���U
�2`������l�5�k���g��f
�� �s�5��k���8���/�"%i�<�=2�{����q���p2_�Tw;�/\̭�Ћ���|�#�ό����f��n�`�)�������q��9�a/L�S3c���R���G�S�>,ِ��>?�z�_��[�kz���S��5S;�F$}[$"�%�W�;W	�ě�Q��<��ݢ�	U(}ߛ%H�W���R�J����3&���˝��5yA"z��$^0a��BUԷ<+aBp��ު�#*�vc�
�t�QzFE�,z/�ܣdkhU�|i��S�6}��&��s7��x��c���=��@LH��>�1�FT[It�q�$/	�`��;Lm����Qp~0�<Y���K��B��f�����Ho��7O���tѨ��o���	�1��QJ>t�f�N��:aF��݂3Y�ٱUj&�IX4��L��W�G�:�Uql���R��jz���㾪�D�,i]Y�F��2ФjE)�$�:r��t�u|yǥ�k5Z���\�0���m��\� �w�2"�q_�����9<$n�9�1��И���˵Ҝ2���эg�B�!���
8�&��|U�&{�����̍V�)��R"��4w�=�>��F�K:�^���ٞ�q�uf��-qK�:!e2�q/�u�9�5J���-�ס�"�C{i�
Xo(�����	��
���k����Vz�ݼ!���T����0X��h�J�|���*n�|�\Wdn�=,�U��"��ϳ��U���>�Z)>�%d�i)y�������Z��?b^FܻJ2����ɢK[�&�H�Y^$4�&�K'�W�?ؐ�z�X���\k9=]A!�\c�xZ}]�@�|D4���&o��g�ʈdU)Z
ZkE�h��إ�Xҙ���o��ʠ�Ήq�wS7�i/�R�P�N��0�|��%L.#�����MP�/5�l� 2���&b�Q׈1����@��5"*V3���C���aL�w��7�ڜ�g���]�Hf�����Q����jy��̐�- U��vg�:��P{Ȳ�eI����C%��dyٶ��^D*	� �_D�*��@P�$m��������]C�K"�9�b�u��H\td���+�}4�$б"�(�?�4�:HNO�>WÇ���I�]d���T-�c�,�������L�����T���ր��V��d����/��J��v�@X��?ܪ[w�D�Qud��$�O���"@g�Ʈ4��XL�@|K�)~?�BKf��Ǽ:,��\��C�q��@e�´2_���D&�5�I���Y��Ц������$��|*�|���*kb��/�|��8�N�"~�N�sJ�Hx��>@�l�w�  �h���M�S.��Ϻ0�̠�:�C����K�`�
ģ�c�鉑��t*�K�ț��a��Jeϲ���D�K�j�M_r�t޹��h��l0��{��ӲSŌn]����M�B���bV�I���d�rJ���/֨�ӯ�t���'�m�� M��h͌��7��0��o�ف!D×�8:0�1�٩��#���a�����w3�kXnba����}Y�b�ikSib!E5(��˒���иH�&���H:�Da�,jB�$(m�TP���2�����
h1Z��h��F�����Y1�6��t�ݙz�O���s���F� ����#�`ܢ��B(���W2�l0t����뗙 �oc�N���*�\)i�0�e��tA�ga��Hf
iM���}��X����-�rI�MG��)�-���h�b��dunrҢ){� �>���v�E^O˴)�J<�8LPsz���2����ή���b�K�{�%���t"v��$h����=�D4^��ɜ�W%d.(K��-M�g,����r���Ͼ%i/�N�2��ė�&�;�����J�Ĳ���{�-���>sn����;����vz�����/ݵ�����.���)��&�	A
����a�w�b��^���3��]����L�p�-�)����� #�iy�����*_���	�hc�}O&&dR!P=�&r���x�})�Mэ��D�[�L��Y�Z��YM8*#A
V�R�cWW�#�=ʚ����u��x��U����)�ަ�.T��`��K��	� t��Q��k�����ha����!����L���ʄ�W�QXva�!��jc誙Ë!�6�	Ü��ʺ4�ϖ���n��.� �֙��ސ�V�s�*���r��a����`)`���<���k�$+��������m�1b���N�i��N�9_�-�L��꥜"W�.��ԉ�6k�'��
|6��n0��9,��{���R�z�΢J__�K��#�3S+۬�Ě�*�R�-(��GC=aj��f阭�+c��&X���ʟ�+]wSU�n"�j��&�� �(pc�ĉ�� [��Ť�`��J�.��H!\��7���QX)|�u�Y���h����Uk����(�B��V���Kd�J,�{i3��hw��f8Sc�H��l��r�;қ��#������f������2~z���dy���´������?���|����C�_y韨������������DL�j�Sm�Y䞘�d�^Y�@I��KD6uT*s-�S�S��#���� @k���=d�5#́+�F��muO
�J"F���a1�/Cc~�ya���47��EI=��9�Fq����c�@s��UC��j�z�\> ���3(��S^�C�ZE7N�1b�ܡϢ��&�*8�,)�G�E$��ZĻr�h��T�&ΚGŖ"�BR�K�H��Ղ){;�bk��eܾ�r�L���9�^�1�e�M�6K75[�
E3��Y��*
J����� �r��}�t7.[ʭB5k�/t�]���&���׉}G���w���[����%"��Я�TmJ�y��.V a�d����T�=YM��'��BS�$x��K�kJ�b��Y^U��f�^��̈́VߓE|������}�� �Eq���'o��ƒ�]���AB�v8��Z�_W^)�d��X�i���w��}kɐ��kx��߸)��W��ˎk<����5�9���G����^�����_�ly�����߲,z�/|�SG:�>���o�����/|�7����8>~������~z�l��e��pJ�LC-��ՈnW�P|����)r�K�|F�J��QN3�&Gi7�g͡�(�h�Sr,�6 ����!��|��Y/EMWa- �� �v�ficC��L]o�,�C˯��`�IB�dV��B�o���F�(�Z�M��(6�b5���M���7F���mi3��)�Ѽ^ete��޵��yf�0�>�l|�JᑠЌd�?W��3��Z�ϊ��w���`r�kJ���++"����8����׎5#�����=�z��@d�4�&�w�L��@@�Y/2��g`��,���2��1���Ю��l,G��ަ��\��dX�FBk�pt�+t���c�u5wnZiOc��1�����X����o}~�V��T\�������`�������F��Z�� �.�::
5Ñ�jJ�+��� \�rc���]�]���E�Y�,�b�WǮ���Z����P��f���|w����m-� ,��g�(r�܉}Y�����s�Z�����^��=���u��|������ }����;��a,��ȯГ����ϧ�������ku����������O~O�,�i6K��e<�G=c9��SMkU����I�TS���:yw�D-o�Qt�k�P!#�x}_�O"���,�^&Q�o4� �����'�@�=.
�=$D0v�3L���)-�+p�(#G�v�pDc�9ԯ�F$���1	�I�9��c�c�}����>[(��Օ��&�p��%��!I=kf荎3�	w֮5fuꦝXl�ᰴ\�`�J�|���g�'2�NG���|���Í.���#k}< ��K�^��+]E�mfkG�'f.\5���8Rb')|��pL\��vݹR"��2'L���V����nF�c�}صG`,#��m���k��+���x�� ��8�L�����b�cƠ�������;�����x�ީ�F~<�S{r���XV���Y�9:5b/�����|�`
|��F��5}�v��K���)��w�a�=JzM`���$�o�����4醦k�#_�:��{���\�S�b�m�n�e��7�G/�n���ۻG����O~����������>�iǝ����������K�ŗ��w��{~�/����ѿs��{>>��O��ߋTί� �`'��
z()aM)f�S�lf_  �IDAT��g5�Iw�"����.����~B�����n:Of,NhJD�n�ɣ���y��m ��Q�QW~���VL��]�&� Ƴ���OV����X
����ؤ�ƈ@�hJ�q7X�ð{�`�1�>;�D���[�_|��HCp(	�ڒY����i.��ťЊ�&�-�\<��|���GP�������?��-WU��zT�Kn�5!�f�Yg�0{ ��ī��Xc�4s#'.�J�hoO��u��UgzN+1^ujfAW�iǶ\��U7G�tG8��=�K��3�5C��ٖ�p��|4{�O�Uva�];�����:s�Z�m�:��������ߏ�t~�x�f~������vh�8��ą0�n�h};:Ȩ����
���~��]J��kCBĕ�| m��vzp}ש#��:9Cww�Bj�h���5s6�/R7�f�N�{U+z5Y��y��Go��������������G?���;�&�e�_W��<z����w��^����������O�W~�<����/��G�_)��Tc�d�������v��J�~�Z�������,�O͂!� ���ݸ$.lZ{`H}��k����M�7~��S�p5]E$~�R��q^$>lTj�4t��},&�M/���cg�� ��Γd�y�MC3��:�[E���ta	X\�'�׸n}Ctd�-��	�1o��d��lo��0'%��2�tJB�cq&$���:Y�.��g�w�=�R�\��+!q�.Dmb�y?z��P�����$�(���T�O��}�$�l�1x�~2��rP�����V�-d�1��KORT�4��9R0T��s��-k��#�&)�Y	���kF�2�ofNb��<��Z�V8,V�K|f�H;�ȳ�Z��v�T���۬�<�\�?��~@݉��hF���B�{8	5�1V$���d���z�ƴ����x!̇tm��I-����$�Y,����S�0t���z8#������KQ�Eh�����s�pw�܏������/���Gw��k������6���_��w����g��G�^����Ͽ�ߛizy��Ov�ףE�.��� K*&�����:�y,:�W�ڣ9����k����ڡs �a^s+��n;�"�)ļtiM3��q.&R.��*l���l:k��C4����~�JP�Y�L�lC%AgRdҪ\E��j���;5'��-�ᬱ�m�u�k�(]�H{%sN���W��X�������r��u����z�Q�g���.D5E6���d��VO�W��e���s<�vN������F��v��;��1�� ��,L�̂��*u���ي�4�;L�\ϟ�>�XA+]�~~M3�e�]�JL��#��A��G��I�f~~J�t/=�%���'��{�}��$fQ�M1�OE�7	���!Q�����"-p�Si�Ji��\Z�i��.���6�� ȣ��;�]���#pB1h�U�Bݬ��*H�i�R��@%W&�s���Ȓ�uGf.L@��HV���R�f.M	,��Q�?BQ��|/����	��ۡ��^�YJ��U&""0))5�vW>����m�}��1��d�X3�u������
���*t��7��<S�4M�,%R9P���Vn�L�^�Ӈ��?��w������"��]�NO9��p����_(����z��s��>|x�~���n�����ҝj�&Nt�sa���"���Q7T4�X#- C�'��{����с�\�8�!R۱����5�^F�f��:@��IkMSǇ�RH����?xM��I|�IC3Sd1IQk�G�#��� j�.&eڒ"J�dݐR-%��k���ՋWA܈Q�����2��klנEj����:�b�b.k��Q#�81u]ߢ��o�ϵ���U3?��%Bh�ᒶ0_qk����u� A���5�ɖ��=闿�4[[Q��Fi����S� �	e���
|�<N�1@�C͊�.p�!� ~G�V0#~Քͱe|��q��5�$�q6�\1�㌏�Z�@�F�?�nF�g��@�K)xZbipuh3�֭5%���ZӘ��9��-_yjxl�� !H`��?�րhE�f����ᭉPJ���1�6�С�5&5ܪv�����VN{Rf4X,I�0�i�0	=6��iz��I�)ڡ�����	!�@����x���Zlr�/��a�Ь�_>	]%�+�����&z[D
E��R���l�H�W71<T'LVYꈣ������+�ԥ-���i���Q43F��X���=���OM�y��:�g>�~���O��k�鹷��:d�8��>�������~��5���O�1=m�y~\����ߞ�ﺩߐ	��w��,��� �p��$,5�2@׊^\f֢e����g}�������J�h�*�m�}ۯf��6j\+���`�������@=6�1�QZ�)o@����J���gG餡�1i3QHڄe�� x�!�����e }��^��;��H�Ecl-��w���D,J���FkM*[a4ʝ��{/r�N��H�2H��O�T������k0(onIa� #1�Q��o��a�;������CѾ���y�̤��ᴚ�UH���E�F�iRw��� +
d- B��t-䦾ah�b�# �Ǘb��R�`�Ó�Ǝ�\���X�X�fB�Č{��/�ܩ��*f����q���|Uw�y>/�dc̋y:6m���T(n�ڒ Fi��Y����]�зaC��[×L�#��b����XX���Xp����0�W��Fs�?��x�b������%��'kv�BQBê�@-jYU3��F7���g���^����C�����ߩ���7җ:^C���oz}���ɀ�������ٟ��O�/�щ��H�R���=�������"�nT-i�IT�匉���V̵����+��4f�Nk9�+9��>�i�d�#/4 �h�C�ޑ� ��mL���;(X��77fiOp�}��E�V�
���I��T�Ĥ1��,n�vf�@�B����2UY��'ن�I\Q�z59�7�5���T�l�#��0.3���b<���ML�,�8�U�9��E�@Y��ςQ��^���\0���p����=^C�~6�{q!�}�E�we\�;7�IE!Ŧ�J��s�2؉f3Uc��kK�����cMW4����s|u>�W���]���9hQN���ؕ~����i�Nu�I���`6٣v����,Z$��F`�lX�S|�M��s�ék~t�����V�`����@�]s�X��8.�R:�]	0�Ep�(�Q���횬�ӊ��ȍ�!Q��DN�Oy�N"�Ռ>�^�ʟ$�د�o\lf�;����<�>��˳?�v�oz������:�[g�>��?~��k��2л��}>���i-�f1��TC�z�F��Pr�~SSx��Q'�_�xH0����7,�M��%�/�x���e8Gir�IA��\gу�/�<l��5�Y`���fj	��W1̩��,37I��A�Z���cs�S�V�ӱ'7��6@�Da�S�����
���Ip(��-a��,�:fs7��P�I�'����i>_�n�Z�L硦I�g�+�,&!�#�%����D���,*>rBк�׀Y���d���@(�N�q������dt�
�}�n���P����z�I�'�ps��ijB�z㳭���IM��OZ�L��zeܰ�oY�΁o[���täj���CCW�>�WL�M��<� �{@�a��%��!��0�4�\�FPW`�'�f���Y���݅���?`JҽѮ���)�?�o�U��l�v��-[���
��nM!��@���4"+N�Ч1IM�L��f���;�\�OЭ|/G�=���n���=�=�C���g��7�����_6C�C����I���?�������֟_&����ā2��e�`>LA�c��:pJ�%��޴i@�8Q����&�-d�i����9u�C'����m�C��(�o�.��R��8��c6���U��{�,����TB�NV���"r�t[��O0td����Է��o�2���<L�SM�8J�@*����m��a���!
��1l�f�~:�ܕ�ZE-k˫���7����"<3WL��\K!2֪�q�*�P�>������,2���MƑ�#������`¶���j���4JKYq&�;ES���v�Zz1f%��
@���&"�;?w��`Cv��``��6'�vu��Cp8����o^�^�ԇ1��Y7˷�׮9Z���C8h"�O��B�ե��MJ�	ꬁ�]�i���X��d�v���ԍ��{Pm����?��xu
�`>���'���[Ҟ&M�U7��a��ٝW�ػk�!u�Q����bj�IT{�b2e����VUek2��9�O�~u����������������=�A_��1t��L�����������G�y�"]/W���il�1��räѱ�-_�,
�{���j�U���Q3$\1���Ř�^��h�� 08|>p�6"u&!\2t%�-��͂�ҹn�p���DCԠ�b�E2ӽ0r[t5B1������D�+C`�L�&P��0�*��60A�������10�����h�n��y��LxXKb��Q�g���D��mg��ee��jD��n^76��6Ĉ1@M�]5Jd;���f�ւ j��o�1�J����t�c
�'��/�|��{�#�@��f�p�n�-�F��z'ʹ\��]Ts��ߌ�Iz���&�Ɔ0bxk>�f�o1�/q��;��ۥС�6���P��oԎA�v�����|Q�K�A��Q�z��s��+Vt�3����oi5���m��K1���K�Ef��qF�Gky6���P3����ڄ��j�mX" �r��Y��	�Xm#���;oy-�tH#�Hb���k>�NR����3��^x��V�[���1}��W��_��o��~�7���������ߟ��N���6k�/J���mJ���MӰ �K�D7r��Wgէ�J��ɺ6f��ߊ���p�s>J�w��-��"��<�a�q�2I�H+#/�����̌��hT`�v%2�XȋuSmb&"��l̤�6�k�(I���+��L?�a��&cj���͎��V�
ps��������p4����[)&��)���=������Ka��*��l�V��No��VB%4��"�=�����C�}ݛ��U��a[~?꠩�F6���v�g�B�
Ke0'�ܲIX��Y*��խ�\�F]��^;pM��M���m2ʎ`Ä¼2�����^�������;�ay�!�3q�KL�Y��� Df
�2��|G|�>!�Ä��}S{7��q�a5C(1q��	h,;�oґ˃2܆���"l)�`I*ˑ1�*Q�2�Ɉ`�6�X_��h;�$(/F�{�)��U!��4���YXҒP�ߓ��_��~!4��h����[Bk7���%hV��$���>�^������Sf��,�
#7�����x���o�����=����ߚ���羚���:o\���?�K���_�7���~�����>�C�\�ʽ\��iX�{�\R�J�#m8 ��@tf�B��`� �Vw�bC,�%�m�����6�(��Tb�3V�}��A:/�.k)w�
Y���jK��<Ka'<�jlk���]b��k)Iz��w�7n�`�_�ّ���ݘ:L�	��6���Q(�*��Ã1� ٭!A�y]�y<݈��~_�z��}��r�''��6�G4[`u��fF�0W��veR�l0h�>�����9T��1$s�H���mV<�HB ��f�S#B��`f�IV�5�
x((���� k��V%w*�����Z�ō����JW5#����_,E�TP1��1<k��.�by]z��]�x���g�}dV�i��{�!)��3�'�V׀h�f�h���;�.������{�l��*X��[:O&�j��J!Dv�N��MZ[�|��i�'��M�G�8U+��!*5Ł39����=�6U�90ԒR0��S��Ҧ}&8%��
y<��L�"(�`�Y���U�
�M�?4�u�⸞�	Ӹ�&r�y@��(z�Vt��x��έ����H�;��ŏ:���ED96L�nZ���w����������5o������5�����_C�����z��O�'?�y�腿���]���G���܎sq�KL�yqgʦ�)�}U�wVBքZe"�.`b�ǖ_l������}�#��ĭ����3�0.-ia.����@��'���(��*�B`�Ʋ?/����H�5k����K�t�K�)^��v2f��Q�`�Ed}(�i�6�kƗX����9>��^e�nY<�8��Y��M�x��)SŰ�#j5`�I����h��c\v�m����ʅt������p-(�^3tנ$�:>y'01�ca�����\(�7��/�Z��y��b9SS�\��jvlpE���.�>�	����/�X���t��������!0[�c>>U�K�4�Ӡ,�;���Ǒa��ʐb�S�s	����7�^E��o��c'q�Χ#u�~��[4�t�e�����g��3"��qpl�)�-h ,��t{3�^��w4�بiaӅ���5C�
wF^�/�C�>F�_��%>a']��X�ئ�ۻ)��n~����_�����"����M�����_5CǄ?��.s|��ͣg���6��ϧ�_��!<�)� ��ԏ���R��TȂ�	ȩCW�cD�w�,J��60^��͕���\j3����B����A��#u3V�A\g�cH��ƶ�t&�e�Y�0�cR5� �u���cU)����ѻ܆�������S�J��:��!��]�O07b< D�M�[�Q�fŵ="�R�$w��~��̟��:4+�Z5�Rc	!I��vhx�
M�,�Y�w�.��J �0��)��B�pu����3��iU%(�W&��Uh"+��1Ɋ�_+n�"�ۙ[�.�4�IN5�Ά03�q��H f�k��
<�1	6��s���-=	������ɴ�&U��QH�)�����v� ]�����J� ��kB~�:��O��.����"�h�)M�L�0�A�����݂˧e��'�������H���Ee�is�=�t'R �僀���lЙ1�9;�1?T��C����T/�Ǻ\��99~-$�Sq+���_+<;K��b.��j謼�ɓ�c�l�s������?�����ߥ��7�����:���������2��������M��{��������H�'���f��,_��^"��s�	�(�֦Qded�@��ȍ8ۙF�bѲ��D�m���AW��m�m;'"���#i��@��PQ+���6NaV��b�(��m�֛����΁7��L�	�/$\̳��:%�6��.];hB_���'��}����T�x>��k���C?r�5#�n�%/L���I���Oi3a��A��I��T�;�VZ������f~J�	�ȵV�閒��	m�Y*2�5�f{J��Z����z�����9�Y<�;���i-v���8��R���(Ym�|�ҸV]/eǈ��G�@�3�����k�,�W�>u�̓�lM<�u����
M\�jc��9Z����1���ʭ[#aM�X]9Z�%aZV����<����Z�t�óM_q���"��#N8�����Y����'����4[@"��Ѹǻ�Ňj��� 5k���A�����2�c-d\3ů�E e���{C��of~#���'<M��q\�^��u�dw��ov��S����
�������1t>�������L��l�(��"�}S�@D̈� Dbt9�t׵��g)g>�ɧ��D����?��f��g����>Pd���+���F��pO��5nb;ɾBP� ��Kmq��L�a���b=0^����k���}���ǤxEW�>��H�3�Ey��`͑�tiMd]֓��¶��6�гb�P�<��qٜ�g�{z�����ip� ��a~_��Z���.\'��%|�� !�U����Y�2�Ԅ!�\�"�j�L��@dR���B�+��"��#{j�v�&����R�=N;��D�b��G���GS��0g�a�}�����SR錉�B��]��UK�S�S�紕i��c'½D]��I��nF�+x����I6C����\1��[�E��2�XO�A8u����Si�hV�ЧJ�����V^Եҥ��N�m�O��|�zsG����r�|�s�f!��ZD�!�S��,|f����.��b6K~?���|)��n�Y���|X���[�â��q�kDγ�<��Ks���A���s�ɝ(.ӧÂއ�����{;�r��oz}���)C����>-ƾ����8�;���TΏ4��[k�F0pt 1�����Q�ś-W������8��f�&M�j�(�����ơL��f�	���2	�~͐2qE|��DZ6Q�t�Q��%�EY{00�����inBk�o����0+�� ��1mŉ��W����6�J�q'��䫣d�YC}|���N�'Ҟ�0�v0�Ƒ�������K��2t-�%�a*$g�U�J�-��X�و��{H�pa�L�O�s�u#TEK�� -_�������5a��j����S�9��M+V�����p'V��D��|gBC��T�Uf��:Y�o�&�U0�V#��:N��s*lI�!ÿJ�ݰO3�L@�@`�"�S2�,:}�}���(��([C�a��1���0�mY���Ь@�f;0��c8o��>�f�^��*��.�}���Oď���t���p�Q���+�8&��
du��1
ݛ���	�C��G|�y�=�9մV���3Y�x�k+怏k���A��g13��i����m�BE[�rN:��-L�c���ͧ���=��.�}}|���}����?�n���v�?Q{��K9�!�3�Y4@m�v�ཆ��{�Qw[��Q�U�-��w�`<H��8�(�"R"��R��������e��d6%x�>C�
�o����f�V[�ig.��k}����^}i��x�7R�T��D�:�r� ;2eQ��T�m���4�I���v{���檀I0(���*�����XCkp��nH���i�
Y%�CXh�5Ba��Q�0�G[�3��w�CۣRCohn�RI�<I�O&���H�p��	PY���	�ac�L�`�HeC%:���P	8��M�#zc��N�p�'�q��`�VŃ��3��q�b��pd�EYΘf�{0�UaN4=��������If�]�Me����@`][���f=�S��H����w��%��%ѭ=�JZ�@�%~�n7E��?
0i��u�%lK���gV����)֏�٘��d'��
�0�ݣg��V�==y�%:��[�ᶉ5�YbEK�J���\�
��!�A����%�3��y�����9bs�L��Εv��z����[�9�i��i�)���3���Ci3wQc�p[��R�k��s�Wf��/N��?t��}���\��ks|�:�}�{���W�m�;_�Ŀ�����w,0�6��=�I�ڮRK桐�.q����t#O�r��T�j�#u#��:��I��%��,��&���m =f���0\#@��^C�2�3n��K����kE� ��tO�*V�cWn����R;�?�ӱ�,fR6�I��pMflf�-���+o�Ό��m3��0�4>�{:������r�tKu���l���TV��:��U9Y�C0q.}7�RNU|�'6AΓ�z'��_�8�g��*�˳�
d�S��'*�)�l$��������S�#H�Qr�F|%N�g�
 '֬8#_i�|ޝ�)��	a���5�n���k��
8�΍=8��,=���Ls!d�R);��rLիL�p4ۺϊ��!P��=�2������q��v��CA-DbL��#�{�GE�o�_��.����uy3W�=f��Y�UF^�Q�0��*=\���~6�U�R��|RZ����0ef ��TA0f�x�v�qz9��nXC\��x�1~A���,��%ca������ځfX�-+��|�`�#��d?8#݄�ȯ��͚�?�x�����P.K]��+���iv*�V�OlO���R�2AT�a)g�����5��.�S��p�C��sLVN��v�s�wg��_�}�����6��-��ua�||�'~����t���������~�·g�� _�j`@�fJ��ZE*�4m6 >�3���&��oVŝ��~Bp��^��]@4��/fu��� ����m������m:Q�r6Q�"��?⮠��Y���gL��F���Y�0�Q��I�Ed����H��[�WG 3��0� ��i��/����FR�%D�<V�Of�QF��n������y5�����pAȨ3sumn:����d�n�>����||�Z�M��)�, Z�����E!Pj��)e����j(�,G�PX3:/�5�{�b:H�Ct0t(m=�'�����T-�\��F�Z[b�0_g���Ws|5G��P�	f�Kn�����,�Y=��$�3�G\�~-�u^5O�7y��\��=�A^�I}��0�P��=�Wr�f���๾��4G�x�px ^���+���$Ѡ\�,��X��v��J�����Z=�MȪ�0�\�}��R1g�@3�7����"@����E[��G��?�����{/}=��C����P}�S�8�����X��?N���ʵ�HL�����b�J��˻���$9��Y]�ޡ]���/�	�R�ȓ�Z��k]�Nc͓u�Z ��M\�Gjc�ƈ� ͚�G�	�`�\þ�s����̆ȳG��eW��-����d�r�t\�3�fib?��0���%y.�Z�j钺�5�y���6���*���Q*�b�B�y˒�
b~Nu��eGb�֔���*���<\�}���2�����9
#����}�%��|�<m\��Si�e��oi�hD\3f�p	Z:=pd�G��%����A���T�ӓ�z��&���"�Y��n��#�Q�fe�K�:��[D�2z3�'���Xm)�]�G�Q�"����֝2Xg`����ڱ��f-]_�kꭅ@�`7��>h�aɪF3�b
c��`������Hy[q˙/voע��J?�������o���3�d&��!����W��0��v߸�g[�֣]��D35R�4ձ\��]@��!/}>2S^j������Z���]��ښ ��/��b��[�����eg&�I�y�y\��4�o~�q��~�;�z_7�����E^{�����ӟ|�����g�N�������X�}���v̱v�<�V@�f����"9��];.��f�`�=cK1G`���c����_�z'��[I�d�.��4�ۂ�-�(�gT`�t{�;r6%��h4�B�OR�+n݊)O
�q��YL��y4�F��3CKU��'G�;hu���Cw�;�]���5�D%m4א,������M����س�|^���Y[��.��*~x^㳚yĬ6�J�V�ִg�'8�v8k���U��1�;_�Å@�a��$GF�K�{�w�4\�6�93��L"���)���M�i�s���2�Oiw<��]:$�`c����nX�҆E�>W�f�K�W�X�D�yM �$�$��-.8f�{u�|�̔��	-\!&�Z�jw�x64ʊ)��SZ1��"p�E�Ͼ `����87F�,"|5�:��,{�M�z�h�����(��̻X�͒k��0
O(T�4ǣtZ���JWi��f%�3�kʶ���
r��.J�y`�9�Iig��l���F8p����O��}.���ϫ2re��7'�s����8M����Ox_��}_]񘇎�C������::<��/�O|��,���/0y�DS�E󛔉��=�c�EtJ*�1����̻#4��Gf�L�LIׂy㛮G%�&Q4����iP.�i��3Af.K���׌�ivS1%D�	I�H���,�Nz!릉b#͢��_��!�Z�����"��Ԛ��k/�L��][��v7�4B�Eb�=�w��/w��)��ر�&�[��=�o�ŧ}y�c�&!�g���|߽N���Fʭ(%9@l�bG��F�Y��c.Zꘉ��@�o���5G*C��`d��B�^J䑩)�
`(д
�,�)��՗Xw�f��"k3oO�.r�I;���j!�����%B�n�\<�a����v�ϼ���_�9m}�͵%�'�B�3_=3�:�U&�P�T�G׽�﹒P�q�_�ԃD��^ph�M�5����pĻ2k)�k�iU<��������N,��}��$�a.<s�Jr|kf斁$�M�1�K�}V�h.��n�..]�b{�\];ZB[�52z-��5�"]�!v�D=����ۚ�#xSt|/��$o�q���}е"���w���[��_�}��g���������3�R��>����t��}�//J�?�H��R�6�3i�M+�RA��Q�����s�F��fk�SB��؄>�G)]��`� vg�N��!���\Ւ4�˝��s���o@���cD��,&�&���>Z\��L>�S�N�����izM���%Z��N��E���~9!�
�D9k�V�����bN:��&K%�5���y�:�����8C�p�NF؏`h%�L�5i���qa�e�ιj�^��5�Zj�Ko��_34�/��n���ay���[xҠ$>9Yh'n�"��E3R*�<��!�s�.0�R��dx�H�L�"f�L�ʑ	�:��O�[E5��{*˟��L0�*��L�j�T_g��Qj�]C�u�9�k�m!�^|���-���|�}LAM8�0������&v���I>��*��}��ձ��5@��OӀ˩@���\I�2k�糬A� (-�Z �)�"]�drT�'�vՒp�]q��5 C�V�����
N���"\#:6�)Z�~3����I�j��H��\4t,U��,�gv�pB�dM��#��@�jQ����V���1H�-���N�/.~��ܻ�����}|4t��������ş{qz���D���$��-�XU.� GD�FeMY4SmɝSM�J��ҧ��C���������MߏRY�D��s:5�_CWd��&6Yw%��tj�5T�`��BFLͤ�L�DÔF#]��{��'VN�d�U��$�4���H1I��G"��W�)Ҍ��_K��:�=�o黑�g�/����ߙ/ lMza����r�+�N_�h�Yk�kᜪp,��Hk�kmr��n&z�k���Z�������))?w�㒯���_���:h���'ZI�Mx�hc����7v�:`����nfo��	ڟa�Yk��\[*x*^�d��3��K׸��߰劥B�࡙vW��/[��p�I&B���f��%r��j�����Aq�!�zt嬸`Z ����w��$�Dd"��A+��O��#������-V�C -b=��鄈�"��8'����}�-��S��K�d��R"������22��� H��pݰ���/.�qf��ƥA�a����O��M+�V����1;������gir�z�X.�����H�����u`�nu���d
*ǁд��e#��/�އ���g�������7�����}��׿�)��*��o,���K;�-��0Aʓz�E����),i��Q�U[*�O{������� ��9�y��2�g�G�jM�0�5jRDF!F=�$8�g�5�,��u�!;I��c;�=K�b{�!i�2�RLL���;2��Y��$�$T�V#vB�w��Y>8p�� �SW��ޡ�[�Xl���<X�����a��U�p� x���g!/%*_������ŭ �U�[̘�ҹ�~��+mO/�G���'^N�-4��h��nγfV����wt{7��e� z�	��y��L��L7�I
�D�8��d3�a�B������T��ا��}�@D��N�ST��.m��%H�8��H{�K����r����'Rⶋ�{'- ���t��]?�᧍K�!����@�
��ʙ#�#荿�&8�>�8$m���_�yˉ�մ�N.0�P^,�ք
��kB_��4b#T�fݭX�#��'��1Ip��N��c}�R=��l�d�"���3gr!����e,su!D��X���Ҡ�.A�Uc-��BK��-VDr���p��8W2�Z�L"R^�ޭ%\w�B�e��5�\Cg`t��[
�eAA!P!sf�������<Оb�#1#��ig�G�'�������4E�8}�n�u����������}��7����7����o����/3�N��ۿ���=�����0	2GB�?�(��E" �����������]�V���t���F:�(��V�{W6���U�Q���5k�y��M���r��|����>N�G	�	]h����NBT�@¡^�E'���^�}�������*��q�C�M�B����&�}��@v]�u��'^$S��s�W�@B�+
�d�t'1\N� ����<=��i!
;�/���O�C?�u�_g@I	�Bjs�� [���c�UP�&������ih��Z��* ��@:�z����K��X`B�^���F�k��ɛ�(���V Ø�"���ڔ룖^���S��C�)����������Z���~/׼U��4�5?{��1��'�́������*�t�+�؃��1�$9���.Y�d��X.gv�
�LښS`׺��Z/<b\��ي�0=�ׂP���r �K�,2#�fP9�ߔ�����0�{%���Y�nD1Edx>Y��B��y�
�Z�����iO�u�D!�s�mvߦ���Z�)]p#I5��h�<W�[�w����ǥ���ݳo�������K�:�a��o���/�������O�6�w!i�נ��Y|�-Ȍ=��b�^���AcQ��ms��I���ދRw�����Tb3wՒ:�lML*�eb����M�JLE��lr?qj�4�>��礔_%jKC��jJ\�gl��{��/����)�Q��l׶��[�����ݴJ9jh�q���}��oK�}��z�dF��ˁ�!̳ᓦ��F~����j�F'��!���7R��1ccT|镧�7ӳ��1͂˞jP�k����,n�Yq�~�� �~v�^)��'X�6���s���^"^K�B��E�;׺ꤘÂ�q�̟<a�F�ŒYe�ZDLr��2a�#z�](�&���|����M��YK�1
�B��;k͌�%���ZDB�X;�
:�w��}T��k�ɘ���'�I�U��?[$H-�p���l�?��Q�~�<��$�q�<Dk4�D�Jv�-B��p��� �{+�{М���͸�T=��-{�,{j�Bռ�Lڮjt`�5פGk&�=UXơN��w,)n�Z���bL�:��8U��T_oj�f��A��&�ql��N7���~wf�������u|C:ǧO�4�~��{�������L*��*�`�~�چn�j@���_��i}��FV�k;%dv�L)�M1���-`fi�7H��Y��\I)�j(I`DQTD�I��J�fM�$�eA���⤂�"�l�p�L��$3�j�j1�r)p��km�#��!$�c�5q?i6QTS9�E��1c�n�K�%u�;��[:;�BO8��o��bm����yY�����NZ�hR)R��J م�"���H����/}�C
��>81P��c-ڠ(�N'H��I[I�ڮʖDR2EʒxI�rxn{���c���9�>�v�P�����������6p���{䁅*�%v*-K-�8]/����i��yj}a��8��|o]�S
�H����oJGٺ.�
�̊���@����8Ѿ�F:	�?�?��fQ�$��⮒�EU�7��U.u�$��\���
��[���bN�������>{7�tyy��q&׬�r��2�I[�g�}$ga�I�5��X�ܽ��z���z�e･+�I{#���lU+�L���I��N�dn1�ų�	t�䦊�x
nM��}O�N���@����r����V�͓b�,2��d�9�H���t�7)/���m�ˈn�n�]�D�F�A��)!���Px������h��"��+�~�?�4� �'��y����������n�O�A~,&s[��w��dBD+���4�Wn&�MB�}6�-�{�h��]���C�L5C�u��z���Z�ZNb�Y��X�z��+O�ɜnЄ0����4Z�����U�@��H�ĭ����._Q�	@�y�:��O�����d'($Fb����u�

H�J"X���&&v�21K��>Z��%,i��h�4deG�5��"��X��j����U����8^w!;i�u� ��Sb�Wtʲ�\精JHaz?�'��(��,V�Q8j8��u�\/�e��B���}�FoA�{/)M���uy|i"e[G�vV���1�:�˾�7Eb�<���)E)�����v#��_���ngF�SI�i�{w�%���c�9�3���8ȥ������ᾍYdB�> V����F�S�dI�%i�z��}(�^��ۼt\�Nי5��Uw�<�{�MV�F���Q���LY�<��k6�����)M����\�8^���Q+rg���B��F�$#��JkΣ(��P�B��wx���.V_�����ӊ�?pB'�'��7^�*�ůB��O��?�~�N:�ѠxH��LN���d�0�۠��Sk�֛��	фɁ_�m��[�w\�a
�/�5�sL	��U]�l��?|ә�y�=5�� =tlY}y������U��8Ȫd���7����RӜ'ʲb�m����� ���N[J���3N�q��e{\(�
�����-��.�� ��I��J��A�}�)���Q���[�Î��1QԣA-dxn	)A5��IEI3W�t�)M�+
����-kz�:�ߧ��TASr�͕9�9ۃA��%��S�K�����\Z<nO*�Q���qF�VS�q<K;h����'���0.!�>�s%��� �D������a� 푄�a
yk�"H:@�*d?�"��9Y�B���lѰ��>"���z�N�ٜ��JsOeM4o>���9g��8�@c:�%�n��_S�̔
j(�ݍ�N{�ŵ�?X�w_�L�����}ʫh���?��Q	�9�I��4'ɔ1��ߧv��Gg`Xf�D$�ͳ
lO��{��a����lK��(Qc��$5)_��n ��kxS�e��5���!t�=�~������o)�X��?�J�>Є�*k7*s�)���%i���YJ���þ}:�>J�B�Ek�czH���Ff)���cL泿��!�q+wV!�	���ロq1q��q3f�؅b`��$�`��K�,����Q�T��تC�Iq��T� M�&�ȣ����,�AW��W���e���1g�`ݷT9PT�c�O�)�4
�A�7oѲ��ER�+q��v��o��e��Ls�q��������Ш�ԉ�@ٳ�F=)6x�wܪXr,F�~�0��g6.���I�A	ko]�>��kLi�YQ0���Sᚵ$J�u�@����2��N�D��(��Q�%��8��t�����v��<���1������|�5{<k�C)c��Dnc�#�ȱ4�Ŕ�[�Ρܿ��i�HѫM��`-`����W(���u�"7H\�ŷ�7ރpR�K�\*�g}�S&����	ux[4H�wm`��]���םt/�̙�����X<02.��4�V_�Mv�c6�/����b�n�>���$��ae��b�P��U���^'�%�P�Q���<�`
k1� FS~4�F]Z��MAcE�ǟ��=r��4M
��܀f��������P�a���:'|`�~��	�q!�'�v_�+�[��<Aٳ)QRW�]�@kա���/�u�}����&�A���Xx�A+\&����ݪЊ���$�4`������ؠ*�#���s�=�O)���4!Y�H�If�/���8$�5Ťdnnv!�D��aP���:�>���2@��\S��4� ��,���0�Ʃ��3i���X	u��+���2�J�/�qԬ�՚����6lx�\"�J�4��u��{�D=>u��D�
[}�<��b�(;�^'��$�\�]�Xi�ѩ�P�>�����\l2O'c5iς�z�t���Z�I� O҃Q�X]�U��'�)
Z)#���R�i��|j@҉�d~y!(C:��.�j��Z�J���4�k��g����^"#á$4�^�2$��M}[#��"��Z�����T1���!�+٧�{'N?�Q�$J��ΥRB�����/�_ϼ��M����%���� 7'j�C����.M�Y.����d��d釪!��	���9Ú:�I�Pi=�`���n���z����r��PԖəȼ��M�|jSP����5-.�\�r^��FOTQpJ�zZA�����`�H��h�(fc�Sԁi��/7m�]�7q՛BcW7��P>��	�.b%��y�7�uiHC$O#S��]�z��[��?��6��p>(|`�~��'��?xN�����������/������%��k4��4;�R��u���ZtP�w�ԥ9�V�HW�m��-�؉Uez�޳�
T�2�%����B�Xד�K�Πپ ��]�6��"�k�l�$_T�G,/��`u�r��j��B�+�N��_"�Mq��e��k$�1�:j��
�zu�3]%:B�q?�@E��i��hh��R��,����C9�z�ht��w���,�ɿ��������ٚ�T�#!M�&b�k��GF#�?��y��zL��V�j�\_>+5�(n>�m��b���5��<zk&�s������j��zZ�8Ϙ�o�o�G`e1��wPWi��K��a}MQ*��Qq.��}KeX�m?*@�Xt���\��F�^�7�C�_�ە�\qF/�;9S���g{�ɮ�R�D%>kώ�[�|��Ǟ��'/*�{���L�V�Q��i(H]-�\��p	&y���:$�n'�+)�-Z�4G=������=y�
_�2s��G����ۓ��X���:��B�1��:�q��"<�7f�O=�0��<vz��&���ͮ���π�4��1.}��j/m_�p������k��%�L�>0B'<��S��+�.][�]S�]�����OQ:T}��]cMa����Y�(Y�Z��-y1�����"��ķ�<#��L��L�I���I��_�t���?�U~���X�t��˛�}�1W���u�l�V�е)��I�8&9e0�I�JcYY��4�����[�θNa,	+Bu�Շ�n-C-��� ��Ne�Z| ��B�6IR�n�� �}��5��8��	�C�~�n���>W�]��7�_A?�(Z�`��O�^��FnLS&ƾ�c�q�%Y\�j=��յ4��:����~�[(��V��H|��%��8���N�^�pe$ZM�0�� {
ְC���cix"�iw��̪_�{
�<e�:N��e�d+O��x&��a�TT�P� ���YH=���|-���SZ�Nd�(�V�9QԸ�疆I2��n#��	�.ԥ2�n����h`��9ю�� ���h��dD*]�Z�T:Fqx�����ܰ���u�Öd�'�/�C�S"���d� X��B?�0��U�I��yN�a�ӊ�d�T&��;�%kIn�!������ڻj�9�8�i'7;��?�����o���k�>�C�(G��J�߽ ���l�� ,��nH����D�Ik�w�ĸy�T ��-ɤ��tr-����Wj��q�2��r7��D>jז�P�B��L�畿퐗����f�J6��mD�k����)�
����&=�눦�Q�g:���K,�T�;W��Zƒu�*y"����(j�Y�d���;l��al�i���3+;�X�b��SB���fT렄��+D�[\�MGd�-c��zM�)4DN=�:�µkW����^�訞�]���BCB�
={�����2٫\��J�C���
�btn�Vl�5��k&d2Z���R��t��Iv�F�dL�Y�$o6uA�61W����qtM���K`&}>.��z�4�����$�Irc�׮�#7����o�K	VerkĲ�B�EY,���k�\��O�"�k*k������?v����:��+��8i���p�>�d�B�N��"�i��PO	e�kG6.{�D�+X,� �`�9�A.t�v��kR:j9������6Eɱ���魨���s�s�'�������],͵8�d�q�i�&���5���(��7��=.n�^�Z_��N1u"r�2����_=��~�������'�4|���	�ޏ^����B�^���m�����z�C!e A�8C�Aݕ*�6S�+����%n��'i�g�v�o�)Li���4� 
Q���=����UL�n���O(�>	O��R�M!(.�L�$�I6y�E�f�m`m�e�V��A]��]�J cR{����ikI��$ܭ�`��o$�\˙�� T�ݲe��V`�FژG%�j*�ز>o��EA���%t!Z�⑩$<n�Zq�ry]��%{�����{޹���1���1^�c����Z��b
�2OJ�(D��k�L����I,2�u#-����nl5=�P��"_�z��
��F��M��#���-N��սU��w��n�Jf1��K��[J�/���$��]�:�͖���uI�q�q��Ե%����I	��:�P\���Öm}�^��0	w�]��:%�5H����9M�
��V�e{ۄA�(PRIc2$g�+ٗ6���I�;�f���
�mu���� �$���s\C�O<{c*#\�48y'��;�Pb��佯_\ir��<�������JO������"�����c��(*��W7}��y�ik��ҵP��\/�;�LLCY��5W�<&�@�=��-Z��j���a�[5�p��>4>pB'<�ħ���/|.^x�~���zI�P%�[�LbKNj�ԅ��Z�dnVw|����Wvg����<����w�b�������a�&�=mz����h��cuS�W&tv�Ic��6�r���ꁐזNh|�A�.���V�-]�E
���dN������ř�
��o(Zn�Ĕ�Kָ|�X-ԥg�:%{������h�Z��������RU�f$Ƕ��$��VE!�Z��ΰ��޺��[W��`	yQ�+�ť�9�.�ҬC�#g�q�9UE��r�F��e�7�"5[Hc^ۣi|��w�w�o�dHw�J�.�����b�U��>���zdm�)��Lt�6I���w��MI\�r�)�����EnL�I�~t]��KhI��]���e���=mߕ.7����qE��5�/��A,�M�c#!�����+��1db�Y��}oϙ$�ir%-���ȺF�g�R�d�^�X��4��%��j��[�2��J'��E� �ܔ3= hY��y��~Sh�v�D{496���e6�^�vN8�������d����R��-yF�{o!ç��ͪ��+P��ȍ�̓*�ҵ�*8�r:��.�N��H�i��6�'c�������h���gӪY��>l?��Ϫ�i���\�Ąb��b[/�<
Mj,������<����3w�~�����a�o�2峏6���F尫D���SM9�� ���q���zCɌ�E�#���t��r�*�q�6h�t��l.t��;V���h�L,���Ժ���
eC�3VHS�2�e�A�K7Y�l�z�'�$▭:\�t8C�$��"�r��YZ��O������vKB�*'Ȓok�|���j���a��i�ꦂ&�˔��C�ʁb!�l�,�(<CIpl�I��m�`�ض�H��v�q|��K��d��}�\�J�7:ɫ��B&���}D���S�4�;���ico9K:�V��J�l���<'�*X�ps�ۚ���w�I��&ɘ4;��Awj9�b:=���uP�>s�3���Q�;��d	�Akι�� #Q9+�:��\�g���T@B��F�ޓ*��B�_	+�*W��h�R̝���w,h�"�9,�q�e��gQ�s	C��v�AP~�m�?/疔���e��NVr��2[�{2B >�l�wFA� �7��e/Fk ��|�z9[�q����������:���Q�]p[�]�?�{����U\�_�}/j�U�6r���q��R�f�Rc�,�#��S��'�`ԺWM ���qSw��Q#ڸ�ޔ���12G�0nA�,���1�F��t#�c,�O�Af`%���d�Z�a��*h��J���?N����(2�%���C`"��ǂ��A�(d�1-�k�o��*Q��@<RJ�5����2c�E��aD~h. U)��U��N�
��.���O����f1�%]��C��=Z�в[��v�I��$Yk�4��n����bm�w:�U�B��f1�������a�8��xC�ߏ�	V��ٖ��9�bR��7��ra�1��0�kѪY�屧,[�+7���J�ܼ9�v�ބJb�9�װr�a�Z�,q݁�A�YQ�4' J�'ae�K!�J˱����K��(��#4�Xs�A`K��^U[�vtTN'�9�i��`����,��M�=@�[2[��)%�(M�,�n�*T���AW��ؔ� qd���hb]R�@�pJR۱�T/��хp��H���Cc�����a&e��"��5OĿ�mВ_�K�*]$�x�h.: ���:c�)6�K��PuU��?W;O���n�M\Vc�xI4�ڋ"bJ��f�Tʂ��U�^�0Q�V�|F|N*9?�9Y�0&}N���^7-W�C���R�Zr�/�/��������gg�����n'�V�N���O�+_�2����E��e\��qH���&+I��<��~�Lw*��Q���x).ҏ*��FLP�#�6^�i��1w���ܻ�@��1��ݫ�d����S����-�iK��4�^�OU���*l�w�=���/{��Cę
Ӓ���j���3��� j[�<Y��a��Y#u��뜅r@YHTz� Y{��G,�K^���J֨�-��ф�]	CHc�n?�۞(y�zt,�m�h�JYS�������.��H�5I��+}��_�x���f�cܲ\��W�/��W��QQ��V�3�7�2߯�,�uȏ�˙�"�}�ʥ�\�0�"?W�N%��*8�R���{��@�R'�����V1�<��mɸ@�.��h�K|��ǵF=kV�i}�y/�v�:s�N�b�oUMΩab��Ɇ�\�.Ӑ�=g�'#d�ܕ'��S�똊G)�(:�ne�]=���ȑc�n�{j�+�,��%�R���v.�o��C �qD-YJ@��u��I�Mq�y;;"UR�kQش�,X� ���^3X��}(l_���i
�����PY\�����N5�ԐJ����E��CX�u���r��zE��F���b4q�y�\��$�X�պ�śh���P}�'?����9���x�O�k���������/�*��&}]$Mo�DX�轕j�4ԥب���:l�K��]Ǐ�#~��|����	#�}��V+dn� �{%i�aZgb6W�4+���|��.1zq�rIP]+!NZ�ir-٫�h���l��R����Cd8}d�DՒ��?2�E�!��?k԰X���͠*B�.�����{� ���$$��������u&���z�ԉ�a�Ꮊ�i�A"mZ�^����J�-m"���Xيl�|R���C(��+3w�`8���J��-�
�uގ8��T �+�_�n�.1�~�h��3�T���+��}>]�qK�YJ�wb}$�2��Eʍ�%{���:tM��9u�WAz�GU�J�@I�,T��^A^�P]��-�J�L�+�QsRc�2fA��ɳ��9�|�f��s�dM�������HF)i�:mV�� S#�r���G�^.�dܩt$�FB� ���i$�Ž6�3B���Tz�_�Z�S�j��щ)򽤿���Q��T��<LZ< ���-%���0����Z�(be�q��i/�s9�(��Xʨ�u�S3 ���&cG%֪��}n��` �EP	2���%���Y�W<�3�g�Z=Wt[C9 �+P/1����m��w�=x�����ے�	=����<��|�կ��O!�ZF����u)�I|7K�G�SѲ!�x���N�y��jY�`��;R�7�]1M*�Uʁ5IPE(�N��2����^�o��H].��$F-/r�U�.B(e@��TTg�6f)z�@b+��`]�Q"���*.�����u�ЊF\�M���x�D�CF���R��PVm�l��*4G�{Ɏ�����<=�M�ǣ�@n��uL�f;��;J*X�nzq-���C�1�'j�E��w�v�����x��䚫�L��o�H�b����� w�+XU��ϟ�2{M�-F�FTմ=�����|+�^�q�&�g(Jb�t�Dʺ7�
�J.�rԎx��3�lu��5V�2���U�)�D�٢\,�}�'�,'h��C�3�!��3�f��B"���Rڎjx�n�l/�qWX�%Tu��ƽ6�[���ɂ\����i����F,��5�?d�
��~M��fz�,��(�;��K�,"2�����J���-���RA�����o �A��	��9潑-X�5�H�Ѧ������_&�Q�&���(�%"�=9v�NUVQ�ίT�؃�=���.(�AcI����N�µ�=S�ሢ�{I;r�4���+(6N�-syZ��j��cH�7��_�����6�W�=�p;�%�z���ϯ@����C�?�/���?��gC�|��ǆ�� 
����$@�����֮d�W6�>N4e���ׁQ��Xڧ��m�wy����$��..A;�j�f�`����ԗ�,�`��3D�����*����|
��$ӂ�_�7��SR����͚`WpP��Z��%V�3�CT�!m�-��@�XIR�t��И5k��HV�l�CqMN�IcW� ���hIqRQ]��%#�ѦCa��~p0��t(ܨ��%�d����IHl��Jb��t��Ԍs��E�2�{��PB�^�����\��Z�J�eܧ��L��]g�k
�7���0�F�������ⵃZ6����H#y-�$�8��Ϣ�d��K=4� Ւ�փ�e�t'7gn��� �0�9��K��5%&�Ui֒�~�	���19|ڗ������)ד�,�O��19�^u$����T����j�������^嘵v�:�6���E��	�=,���ZR�j�O�f�	�LT�C���Ʌ��a
o���> "��I�8�4KnJ�� ,��D@���|ǩ�3UO��q�G��fYy�dY����?��-���\���@5�6h��<�|%��cbŻ�F1m�7��vI|[��ڠ���ј��a���7ˇd �m�ۖ�Y|�y8^�w�}.����I�^jQ��HO���C�Ƣ>��?&�$ǉrE��=�荹���d��n7���D����`�.��h��t4�¶�*JҊ�b)�RwwaWq�	���I	'$��͏�Y��5g��T�����,�54H�Q{�S�N�U^_�c^�Ѭ�&�����3Z%<a��W2�tDx�;�噄N��TŁ��� C񺌖7e���V���	.�3��I�Ww�( D���d0Tx�U��� �*B��Ư��O-�0;|��]�d��m5%0�2w���q�P��!�g{���d�۾�mkC�w�ޞԘs�Lً�uk��F��6I;��Z���{b͉�����L9-e�"�n��HP�ӾZ���Ui��@�A�#���A88#V9�zck-�Ӊb�`��i�&͸&�ǀV�M���U�v6o�H줎X��������D�Ǜ��!-0/Tֽ��}���G	��-�m���j�35�$\RI�'
/� �6�l��x 7��v�B�9�aG���r�q�*J�8U�?a��3 xhL��@��A	m���P}`J�����X�)7�ph��qw�����XVc�>�J��_�\��e��be^�M޳h�ǦfoFl�ȑ�c���j��c��w(�^�f�����O}nWܶ�N�z����P���֟�ׯ���M�#A����EU7 Iz��%���Y�>ђ/�]i2�%�A� L0䱄l�v��k�6uф-b��64 ST�byۈ�8r��q&�;+Y�pbA�d.1�ʬi����c�f���$�O I���$�
����3H�-�zm������ɪR�z���3�*Q]��#��e�o��hw4�ɯDC.J"t"\��G��A��*����RAM%y�mwx.����h-�C��H�ڎ���p�~ 3_$�ɵ�h���j��!�۝�}��ys48�u�y�<>�|��3�D,,��NvKj9������
E�!�CY3]Iι�V=�<�i	�*REԵ�h�!Y�e-J���F��B�Z,`���A۱��B\f�myźi����Tޟ�J�z��2�%�H����� ���b�ɉ�3iX��QL�a3��\�O��'e��7({/G\^OϬY�Q=2Y�P����
!�\ͻ3�sȹ�p��DJ-�zɌ�G���˝�}j"e��j��=��{�ۭ��P2�%a���R=�$����/�+X"m�Ŵ[�I�9��b	�lR���;}w�+0z�FQV�h��M������cA����>�0>є$�Už����TR02W��p�H�5��|�z4W��r�B�.�D��oլ�/:$�\U˟�Cz�r��nw�քn���O3�߸�\���g��������!4?��Ie�S��#$Gc�<���9�b� �U�U�2m�-��!Z�n�ʈz���Y7����J2vp�;&Vݧ�c��ц"p��������~G�+'j�]1���A\���k�߭UI	�5Qc�Ԓ�s4��F-
���!n�v��V�����غbwk�b��+{���'P��.^��=�q],ީ�0��ȵ�+ֳ�ܐ�̍I�\7H�[��\Ԇ�h��.�0Z-Y�H.�Z=��s���`��jA�׀\�76'���X-8Y�d�w��U���%T��ג��sE@b����"-��Y�GgP9�a�e?�d�h@I���n�0�=6Z5�	�L<�5���ֹ���s�xr� ��:ƽ�
�j��O-�$|?���Ru2��C��FؤDp�ZK��
�J��l������ZA<<i}��׮f���^k8E�kU�wH��a�~�C�!/�hF�Bk�#�2ds��W�ְ�Gr����V��\�����Ӽ%S��D�y���I�,I���
g�:Vd���Ǧ��G�RP�]σAHq��O�q��'�-�V�m@{8�~$��C�A��-�r"p��̳0���kv�x�H~�"4��EA�KaHN��*S����*�n�TH>����LHk\=�&+��
���aYD�?�"?�'�j�0�2��]Q<���V��Gqm��\w(�i�������	<��!�	�#�@���g�����z���C�Z]���B��'��-����J&�����"n�G$��PmZ�.��`�m�\�<��S����jYVy.����r7�:���TTy;ZU\sJ�6j�H�s�� �vF�>)�UK�k �:r������l���H���G2'�Fk�}���9���X��Ζ��Zk�Ce�N�����oL�Wm���X;�B�AR�
��E��p������.��Ξ�g�(�q]47�b�~␥��NvN�oT���5s�k�ъ	h=-�^���.q$�6���E�B䤣�	$vj��F�v|�Z>xz]���^Q$��T�E��zy?z8��q�,��Q���e[�1����p�)F�R��Qq��~��ِ�k_�U>��t_�}�d������<��T�f���M���O
MF�A�"�E�t�%O��uK��-��r-�w^�>[�k�Q�q�k�G \��Xq���Zs��4����j��p�����S�9��%��W�R�{1w�ZH�hl'��&q7�hw�bFY�I��d��6n��^,4�Uh�u�%�tpB���Ǘý����!i�y;�%�����Xն/���|Ơ�"Q�[i����r>J��
�j[��Y�:��CDJ����l�C�|4����=U�%ᶳ|v��	W:i�f�QbŀY�0�H�玨S�Ԭ�gMA�Q�{Z%��C�a=b{!��G/ʤ�B��0sJ�kv:{���5؜��j���nu�9Y!RWr���]��l˟�o\���{o�'��?w
�B'<��O�+��[p��5��ۻ���_T!��!�3�.rS��I�[�Q�vu۳�*k��ˤ��n\M"�Q���z��c�C��E""-�,�m�V��e�ns���� h�%)U�M�� G��I��c��JL�W	�H��Įa�~Fb���fyJ�9r�#*�X2�7p� ��~�]���#�5J�.����]6�Y��D���c5�HDQ;�|wH�<�hN�(Ԯ�G���jl7��k��*�u�8���u8IC7p"`�y�(uӲʋ%~�~�3�U��9��<Z�QP���w&��A&�H�Y����Q��E4�A�Ȃ�e��(�"�����mW�t��G����l�Ӿ�4��%�dE�p^���t�0����7���AY}=�(�.D]�&�Fk0AVV��aZU0L	[���1�(�$��p�uv�C�l��5D�Vl״��PO��!-I��Z-�;�pDb�j�"*��rW���B�ˣ���2�Y��� ������#!$`�d&P�~5H.^'Zbʽ����Q�V����U]m�.Ħ���#�-���)��7��v��+۴��Ks_]�����JH��Lu�vx�jT�������TNH��j���zsX�sV���Ð�R�V��W�\.q?��=4�q1�:=�\�Kwy#����Q41q������ቅ�����9���k�.�-d��iv$��<��*fu�P�zr4���H٠�<��5^a�B%��h��F\*��(x�{�ʆ����Xvb��.�ZF)�g"���J�ь.{��g�Wb�V���Q��Q�X�bY�I|�+�BI|!^�f���,����1}�������ٳx�"t�C��,o�7��ē�_��O��V�O�e�yLÉė��Q��q��D+Oba|��Lgس�'km��PJ
��Z�Z-��>Z�&2o]�&��nQ�p�8$��e��]� vF+}�b��#�wx���-#J<�i��sſsc��<b�H� q/���%�Y����Z� '�v��AK����+�~R�e�[�����n�����W�p�����5\���/���2.�U$�׸G���]�X��B}[/:�h@7�Ӵn� R�p�\��U�w�C��v((��t�׳�;��.���>���������^v��� �n\l�M�����nׅaP7"+����!^c��~��u��w��Y��M����e�J��A'�U�S�H�BR[��s���a���FJ$h�C���z?Fϥ��xS��ɾ<���$Dݖ��&�
��޴=�yy�=�+.q��?A�B;$t��}�V�uw��D#��<`�/Ń�b�-l�lmqQ��X]8�;T���0��AJ���G]\v��h[�K$�x�kz��^�k��P�����2��w�ڽ�_߾�� �u�&$X�qs�r��'
���?h=�m���u^>�_H�[|�v���&S|��^��>8�͡AM�;�Dhq��M�Vx-*�^ց�N�~�q��H�UN;���5\�}� �����ݏ��}H�w�НG�=���p��Н41w�#��q)���%en�zt�ā�Ns��Z�T���z����:����{��w�No�c�Q�5I�,T�F	u}�D4�@�X�6�z���0� ��!�� �s������h�{R��n
�O妍O����js'��Z�|ܰ��(H���Ԩ��2��k�ѧ�iE��2G����-����x�?���7��y�ﵗ`��rG�9�#t-�~�wP��p�Ƶ�;8�s(L��������5�!"Yǎ����L�x&$Q_�@B9J�hr�es�I���d�����Zp��y�S3�\H���r\��[��	ʞl��O�to�X܊�FΐM%Q�c�<@�e�)���>�Qk���J�
��@?j�pnyG�#~7���Us�(��j9���oT�����[H�#���/���U<@["�����W]up�{�׿ԟ�A�Qfi�K�_3��?uir��iK�5�U�<X�Yۜl�dr+c��%���������ݠ �"4i�^���~l�K��\���~�#$�����n��l6��n 5���z�����1?�-���q�h":_��Q������M@	����|�1�
:����n��Dj���Mlɶ�f���py� .��.Ƹ���N��,[p���~�|�;�] �P����:U�m���&��v7(�#�B��琻���b�"j4����6������q�9Uזg�_Y\�pyu�~'��o�@}3ԋ�B�ڰ�ߣx�f�}Ŗy�4^�!���R1b;��_L�K�Hx�,]r'�����Ac�T�-c�Xi�m8����w�F�;��&�L�{AO.���UؑK`��:���Dq�ł׏�B��h�{Y����vp������\�w��߷�ۑQ�ˇ�Ck���=y��:�wᛞ�ϵ"�?���,��!Y���q�d̮ǟ��S�n��c����F���e`�@��<}���ND��a�{�q����[.��n��Jz���u��$<�Zb�[��l^'%s+k�����v������}WNy��W��/+�r;��V��Wi����Y�F��پ�󲺊���������=���O��w��HB'|�G���߅���~m;�����PX�d����Ń�ڡX޲�=R�&��(]��еW���K6�KLJL�=nM�y��ꂆPb�c��>b"l��*��)��ޟ:`��6�a���
�#�A@�l�d���[�*J)	�&�Y�4U�������A��H�0J�_��K�a�d~����g�:����VF��hӄ�JU-�@�~ַQqx5ٯ���Z���^����������HG���hli�~��m/]z��o�	��ٿ�����ݖ��+W�c?�ɗ�{�꿼z�$�a�D�ۊ\���=���:,ֹ:��!�� ���dǡ�Y�f��F	�A¡(o=�+5K�0>�+[��*�'��"IV��K0���4b�>����R��R�BIh�i�D�I��`$T�2��p�Bi�X��}�2O��b�\���d��B�H���ˉ�(u�'i$V4Gc�3�EB�#����;���v�:i�o��^Ajg�8�:���7^�]?��uj����Q
�uj���9o���~t,m9!Z�v/g넚�7p�#gҺ����vB�r��W�n���.�;6*���oO���z���owpR�~�a������Ο��G�k}/��9o���_Ev�P�n!+�t���aN�woK��q�\�DbC'������͐�7fb/�8
U2���w�d�G4j�G�J֕�E���Yy���%�4��/�p~���I�h��_F%j�ʰ�%)׭J'�`�K��?N>b2�ѧ�6��L�d��߬���@��+�t�R�g`s�;��	w,�z�3��W�
���`5|#�.~%\\���
��>4�^�?��8�Q����<�O$��Y�͙���'���2�lOg[Z��ru��%U����"�ٲҿ�	���F�����gPK�̽Ρ'���.o9�k�VC�5�T�E�	:��)�V�~�R# �Q(!d�u�H�+����� �����M�x}h���������U��.�on��-
��,W��/����?��
\{�X<|�¦�s�>?h�s�={_E�z����ۗ�f�u<g|�RF��e{��1��������֕����Cv�$��H!��Ą#I��=>A��k�xf�'j%�T�eXw`�&�Hڿ2T�I��Gz����m��%>ߴq�*�K��5͠�1��F-5�*�!*�\8�2��@zcw�M�7�|J�+�DCjC�6�ɐ6'h~o�t�z�h7�]}m�߻֋���$}���,shW�w#�k{p.��:}�����/����+��e��[�%��
�~x	"��;���������;o���Ґ�7��sz�܍js�2Z��'�6��u����G��?��~�nG�P����r��2��8ԱC��lJRd]��N|��4�r�* �I�t�����6��dH\���k��l*��ȵ�垄F�)_V��:���b����J+dU.UG�=��O���!X�t����K$��ߝ�KnO���m_&$�o���l뿎g�J�!Oȣ?�����;��	?��q�~#���W��r�8�%H7�L��O��~.��n�f-���dِ�HIEÄ�7�5�3��57�F$�U6�&Lc?'*�;&⹲֖�
%�!@Bo�^�c�t���I?�	l8Q�`����T�R���)n[hK�,R?�0�S��-�s�sp��\::8��^���ֿ�@|�^���f����=���܃�!/�5,P8����gΜ�����>��0�k�������j�.s~)��K���%�N�ڲW���TJ�n\`h�M*��U�'�Q�"HV6?��9.��a��!<�÷m��?��Ko|�k)�T���1�_�����.n��a�1<���~�$�\��uX,Z)���$���8�N|����u�Է�ݓ"JCZ:ɭ��J�c��IR@���Gi����q��km����3H�<�+E('�-e�e�����H>�(P^�^GfPJ���_+�#��i$Q�t�fGTy�8�8���"��b�:�T.7������t��>Ń~���쳴U�ͻ�����ڍ���t��:}	�"n�� id\�H��Y��u�41���btO">Y|����ӕ���!
��՗��jާZodͷ��fj�X7�ȷ${9�PʤB�2��ي:�5�*����w�"m{�!�Ԗ�X���$-O���s�5�Ggw���}$�g�����h��[��~��k/�CIM���
.�}8>Xܩ.@ǿ:�}���{~��Ǐ^����w��/��������'и�h���3�$�����Z-������D1$�b�b�Z?*\TRB@y,�X�r�k���ٚ���+�d��/�v)�L^+�8���<bd��h�`��`Wy��r��1h5J�<k�]F���,L|Z8�]z��?�FJ��f��|9�����Z��̣�l��yl\�;�"t�O=���<�?��|��+9�r����ٕ����>R��'q��萺�����4,�Щ�$��H	]\�b���&�b�2�hY�v�K�����3ژړ�T��5ר���j�r��~♭�ƭ�7{��ó8�x�")d������$C�tc�8��ษ��98���s~���K��w��/��ڷ��wp�O���1�;w��ӟ���������1ʧgК|��}����z���Ç�j�4��g}�m/V�_"�י�Y�Չf$SZ����X���)oП�2�M4`'�(\6f8LYf2����ÛF�s),E͠�w����DI��F9Zd����
���r���Bo�3וe���;d�kh��j����WQ���ܝ\�t�)��k�|
�Y:ᡇ�m,m��~�����{��p?�,����a{W�ǐ�?�W��H��"��C�z�O\DH�B�9Qt�i����Y�Kq2}|��5sR3�?��Y�U�mm=ZWK<;8�jNT�4�Hڌ�,t�~�עl�m7�*�s�,Z���耖,�1�%F��`}p��ѽ/�q���_;sp�6�o�&��;����p8���������y�m��}���s��j��'oý��O�����w�ǡ���L�|h�Ȣ��{�d-o�zhTlHy!֜u������B�y�|#�2�����[ו���9��N�0-����9j��t�Ci1�ڕc�A��$�)ɓ�Q�	ߏ2\���'U����_����0��LP����;ys�{N�zl~�l	�0uURS���z��2R�ej,������_�{C�°[��{���Cx���^܄тG�χ1!o���?�c������\*rB�9k���E)��[[�ɐ�=�h;�4��l����i_iz��[TR��N�� ����j��q��qLK�:����"�`��{��їV���}᥯\=\���K?��t�; ��'�����|�$��}�8��<t/T����rN'G9ԗ���c�2<����!�=(��#C@�-�|[�����]�=2��c	&��A�zγu��ReI��)�|�&"�[Ge��X�6�Mr�Ř 
06�	eh��:�UT��>�K&����->�?�5�
�ĺz�m|��R׿c�^W�Js��;��g�Mf�>�0�����Ԕ���K�C��}}��.�[H�oqV�嫰~���C�o��S���U��R�8��de�zu��zf��7�7�7��q�-mkf[���1�1p���)Y���#nY�֋o�bt}r'�m��]�!"�䦪B��h���n����i�r������4�����/_���g�y�_<��'O?���}�U���08�;��G��dI_y�۰���&��d�7��_|��?�{��Vi�[P#�&��������Q�܅�~�:,�a8LCZ#!���u��9СT�ID�Ȃ�
r�'9^8�$,iD�!C��F5�q%{��Y�Xq����ax�o��ȚjJ)��O��N��ŚH�*�N}
�B��F�����Fc�*�G�]l���K''�|��q_ ��ݯ�Ï���o��?�y�3��"�)��'���{��p8�=��V�M�"8f�m	��p8�9�	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8��	��p8���o��<"�*}    IEND�B`�PK
     �9s[d��   �   /   images/d3b73945-fe79-451b-b309-b64aab767520.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     �9s[��Н�� �� /   images/0657d52a-d145-430e-bb7e-5d1be0618b5b.png�PNG

   IHDR  �  $U   �:�P   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���y���}�����=��13<��!�")Q�$R�D��,q�X�ۢ���bi��.��n�E6�i�x�,�6i⦎%Yr,K�NR�(R�I��y�������?H9�E�:�|��y���C�������~�O28sV           ��B�            ��          ��0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\(�:   �h(|�kQ���Y�    �1)=x0�oۚu   0p  Ɖ���b1�    06UTd�    ""��u            �0p           '�          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\0p           �          �w           r��          �\(�:   �D��~%��=� \F�icD��u�K�����Y� ��ͷD��e����/�l�����!��6�   �k�   W�ȿ�w�>�T�1 ����]MMYǸ�t߾��ײ�0���Q]�u�KJ_{�� Ƹ�'��dɒ�c   @��            �           䄁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�          ��           䂁;           �`�          @.�g    �zk����&�j���"�/\�U1PS��1XUI�IC��&Iz��(�D�p)""��CQ�ʾ����������ʾ��=���=Q{�/
�RF�b������i�����Kv�Pe1Ҥ���_62eC����Q�7��Q�{��u>@�z�*�gRmt7�D_MEVUDM��ί����u~MW_�w�F]g��   ���  �e��<:�M�s͓���!�ꢫ�:�jc�|4W�Hߝ�i�t�G]gO�w�F�ٮ�r�#��>�����`��(����q��!ڧM��ƺ�x#SV�_�����Q���g�b�鎘r�|��|�Od�X�S룽�!ڧ5D���8�F���Q�>F��D}GO�w�DÙ�1�􅫦�o�    �w�   ���������:-ζ4F{��j��H�N��$����詯�����ZU�`L>�SNuF��s�|�l��@\�p�,�̘m���ٖ�8���5�&�)�4I���:z뫣�u�{~�:�|4;-�κ�	���ř�qj��8�29ε��몢���}�_�?SN���m��|�\�=�F'   �q��   ���89�)�fM�S��ƹ�IQ*��	��诮�s��Ĝ�x}݅��u�D˱c�G�D�ٮlCdd��"NΝm��ũ�)q��1J��?��v������c��ع�~�L4�9�qJ�lT/��o��fN���'��������ŉ��⍸�������:�t4��:   `�3p  �	(M�8����N�����1=t�0�k���6���Ə����??3�E��p�	���i�qx�������P�_���q�T��B���D�����8�P�_x�SuO�<x�B�:C'   �2p  �	�T(ı��qh�8:�%�k*������ػ�6���e#�h9z&��=s�>սY��DJ�B�w��-h��	���u����ؿrvJ�h9z6���=�Y��DJ�$��k�C�̊�Z���*�H�ꫭ���O/���D�}�h�t{�   0�  �8��85sJ�fVX�:�G�d����6��ͱ����|�\��{,�y��3t��S*�Ĝ�81�)��q�/:�[�����˝pY넿�郔
�/:���W�|   �1��   ơ��I�w��8�|vTUdgLI�$�fM��YScǭ+c��S�dϡh���R)�x ���4)޾�B��W����}��t,�s0Z���B)�:��tL�������������U:�Ճ1��:    g�  `�)/đ�3b�yq|ns�qƅR�GN�#�GM�@,z�p,y�`�w�d�����s�#���}�B!�,h�#Zt>�+:���$�.h�����(�u,����O��:    a�   c^Wcm�~âؿ|vV��3n��Uƞ�����b�S�|�h=x*�a��U��Xo\�8�����޽R���=���çb��}1�`�������x���:���+f��{�̋���Ō#�cŎ��z�d$��   ȊO@   `�:;}r�~��8��5҂c��4I����86�%&�wǲ]b��CQ><�u4`{��.��B!�8Gq|ns���=����:��ζ4���/��W[qbNS������ʡ(��    W��;   �%I���3b��%qz攬�Lx�'��[��W7,�e;���]�b`(�X�x�D^4#^[�8�fM�:̈́��X{���_K_��^���Y�Ƌ$�Ȃ��E��:-�4޻����kb��b�������|   ����   ƈ�s��-�����YG�W��V���+���c����������'r|ns�ܲ"�Lo�:
����2^޼<^�qq,�u(Vm{���D��m���Wę:?o�j*cצe���E:�^��   �w   ȹ�s���-��a{�TUĮ�����Ɗߎ�/�򡑬ccH[��xy��89��y7TQ�=���΍e/�;�Gq�����Z�Ʈ[�ǉ�:?������纡   �*0p  ��:3�1^ܺ*�Z^ƚ��عee�q�����7c�?�$M����ٖ�x�U��cP������^k�{�B�t>���57ċ[Wŉ9MYG�#z��ַ�.�5Ͼ��9��   � w   ș�ڪؽqY�}��HI�q����{��[k���'���#g���LuE�r��xs��?���U�sw����-�O�YOe	��?~��Tƶ����/��O��ڲ�   0��  @N�
�x���k��,f�Qt��1}`s��2n||O�u�d	�X���[�-���P�����7���'c��D}Go֑�����7-��
͍'�S��t�����^�   �
�  @���߽6�k���td��81�)V?�f�ܱ?
�R֑���=-��gm��\�u��#���ͱ���bՋoG��f	����S����F����pY8=��k�k��k���u>   �'d�   �,�K[V����"���p5����-+���9���;cډ��#W�`Ey�ey�y݂H�?���������������t�=�H�U2XY�]����	d���6-�C�̊��+����:   ��e�   9�pF<��譫�:
ho�?��X��`\��Q�:pY8#��ku��Wg��O�?�ږX���㆟���a�;�`zl�{M���	��iR<��-q�+�↟�����#   �9�   p��WWĶ��ġ%���B�J�B�q��8�pzlyh��}a�*ƶ������YG!ci���5���������hv�/�;���q`�Ο𒈽k�ű�M��G;���٬   �)��   �DrbNS��[[��y����x䫛c�ƥ���� ����)��7���]�5��W6��-+���a�8=sJ<�����GwCm<��-����F��cY   ��	�   p�
I���}��Hc6ޯT(Į���������KQ�ѓu$�c*
��%��&7�pii!�=ǉ��b˃;t>�a:��I�$޸~a��95�<�#&�wg	    �    W���u��7n�]��sY��y����X��Xm��7t�2NO�~�8�lv�Q�����6��|Hgf4ƃ߼-����    �c�   WБ��������2XQO~v}<��(K��qtAK<�qv�䬣0�V���]�|o��Xqb��x��[���#�(�����    �S�u    ���=��˛W8���m�y�1�.n}�Ũ��:�At>��B��ǭ?|1jz���|�w;��Nm�cۻf^���[�=ߛu   ��q4    ����b<���c疕��|bm��⡯��gN�:
p	�����oܤ�m�S��o�m��f����b<��:߸�O����x�k�F[봬�    䎁;   ���ƚ��W���-YGa魯�G�%,��u��t7���_�GN�:
�H_]U���M��·<魫�G�%/��uƑ޺���7����   �+�Y   �����)��o�}5�YGa)+�S����kc�soe&���'��_�1�j����8T*��O�����X��[i։`b;���}�譯�:
�P�P���^��c��F�*}    w   ?�ff<}ߺ./�:
�Y�k��T7���(��_ ��̈��!��:�+�b�w5����B��u"���.h��}f}U���8������*6��(��   ��f�   ��k��K[VD�$YGa�xg��譫��~�#��CYǁ	��uc�m�t>W;�s�gRul��Q1���jzs�x��k#-�|��C�̊��ʸ��u>   0��    cٞ�cǭ+���o�yS�WWd&�=ǋ[���\u'�4�|���lX��\m��Uwrδ�_S�u   ���  �ǑD��uU�ܲ2�$L`g�7ƣ���UYG��-��q�J�O�ζ4�#_�}u:�����|2u��1y�����   �e�   U���k��u��N�1mR���M�[_�u���n�6^[�8�$�S���l���ڬ���t�&�]�e��sj}�諛�K�   ��;   |i!���]o^�0�(��S��6GOCM�Q`\I�$���xc��'?�k���d��-�xnb%W�j��n1r   &w   ����mw���+fg�ާ��&��M�WW�u���w��wV��:	�OOCM<��Mnl�Q��U���yYǀ�驯�G�%���  ����   >�����k�e>PWcm<��M�Wk���K[V�[k�g>PϤ���6Fo]e�Q`�۹yE���vr���:~�����|   `�0p  �a���������9�>~�śc���u�vݲ,^]�$�pY�'��O��)�*��c�ƞu>���X?~�ͬ   ��`�   ��ʍ��0��kn��~�.�eƜW7,��7-�:|h��&�c_�9�*ʳ�c���ŮM˲�Z��x�7�`��Y  ����   ~��f�˷,�:|d�fM��}v}��$�(0f\�/m^�u��NO�?���(��֡kfŎ�Vf>��:   � ��   ������E�3FY0=^�uU�1`Lhk���w��g�:��%�ݹ:�0&�����{}���gl:6�9�ݥ�  ����   .�sj}<���b�̏Όmo�[o\�0��k]�������|Ƽ�Wϋ�nX�uȵ�ƚ��n��bY�Q�y��y���%Y�    �"|b   ����2~�n���b�Q`T�x۪8�xF�1 ��k*�￴1�k*����[W�ϯ��uȥ����7F��g��yˊ8��5�    ���   ~I����>�>�j���&-$��}�cZ}�Q WJ�B<����ը�?��B�mi�:
�JZH��O��'�eFO�̽���铳N   0��  ���x����:-�0�*�������YG��x�֕qr��g�./�'>�>��+����s��86�9�0�F���gu>   0��D`|H#�#�h�4:"�#I�#M���Rw�WH��H��4��HJ�i�tEDJIW$����iIRJK��$I�w�KR(T��imDD�&����[QJ��$
�i]Ic����Dc�{. ��:�|v��vA�1��9?�.�������/���e�����Yǀ+���6������l�$U�Ll�όWoX�u�bzj���w}��HJ:  �z���4Ҏ��#��H"�(t�Q�.�Ig$�p�:����eIғ�J���}��kʓ$��.��")�'i�!��L"jJ��&5Ic���i�Ic$��H��ph. �3pȷSq4�8��q"M��$J��$9Y(��JIr����dr�PG�A?�t��i��Rs!ʛJ�Ҍ$
�i�6%I2#��%���1%� ����4)��{m�1��;�hF�ٰ$���v�Q 3��&ų��|ƿ#��+7]k�+�(���)��̽�E$Y'�+����ؽqi�}�ͬ�  L�$�dq8I�h��Ǔ$9���RĩB��I��U������1Nχ4"��������P6�\J�IMi!mNҘ�F2+�h�H�FDm�y��2�Fz2��;��$��i��$��H��,/?�:ԟu�і?~&"�\��ҙ3k�tn!IZӈ�4
s�(-�HFĢ��y `�V�����Ų���;Ł�RM�`oq`��|h��0Rj/+���ᑡ4���~_!-U��k"��Ჲ��Ų�����ʚ���b�X$���7-����1��鬣�U7TQ��d    IDATO|~C�5:�*�K�}}��C=�C���FF:
��y_�GZ5R^V{����e�F���j*k�t��۽qi4�h�Y۲�W�p�<����,fe�)��.���Hi8��|�����4��Hy��b٤�bY�@uEm_ue1-��Ѵ�ƥ1�ع�}@� ��4�8���/�d��q����iz�j����ΝCY�mIDmm�������M�̙<X*�����RDk�&
QZ�F�(.�:��Ff �'�� \y=雑&o$I�F)�}I!�Wܟ�>ݝu��J�7/^�Λ�840�0M�E�$Y���2"�FĲ����Q�q`�����&�cZmw�`mg_[U�������#Qz���l�o���~�?�o��튩�^[W6��`Uq�@U����Yݍ5���'�~i!��?�.>��Ge����#/�~m��\�u�1�����|頻�����������ݕ�F���r})�q�X�8X]\�W_5�|C]]����H�$������_<U�Yǁ����VE����c�i���Cu]�mU��oWm+o�o�����W�=��r��O����m�%##7V7TW�꭫j���_�ܽ��g�≨�w��  \)ݑě���I�o�"ގ��}�t��=y�ĉ�1��Ç�#�="^�ԯ����*Ǣ�PZ�F�HҕI�"bnx� ��Μ�f`���7"bw��I�����ЛUmm��]{��e���RiE!M��I�*"]K"� �X�ߌ����Y��@�_�j�O=�u.�������벎1�L:��]���jU��c�e߻�?|�������ņ©ޯUW��S_u�����R���G1w��������+�ݻ"����qI�]1�����1�Z2+�����c�9�==�=�V��4)O�wǟ������I��ů�?�;�zݹi�ZF����Q��w"��۳�1&��Q��C��g���/?�u�1������o�:Ƙ3�������������J���?{譫����3�_�,�LϤ�ڛ'5�Y������O&r���'"Y�$���:�7e ����p�ޮ$�גR���~���ɟ�t\]iSS�PYղ(+�H�dYD�I"]�|c�L8���鉈=�+"��Ȯbm�kɾ}���X1G���D�߽�����v����4bM��ڈ�u��p�; Lh=5���Y��FJ锓�k��TL��������Yg�������O���kLϏ�����/�mnX�_[e�x?�ff�}�X��P�Q��뭯���Y�u�1�l��Nm�<Rs��G�������}ɧ�]M�~����.^�ȿ����������K�W��V���8�hF��f~,�}0�(p���V�s�\�u�1�0R��mG���=R*+|�?��׳���?�+"�{������G���U�f{��սu�>߼�#Z������ ���xwӑ&�"F^��ȏ�����q����Y�Zi��,bmDamza�>7�� d�@ �W�HފH_�4^�Bl/;�Z1�u0>����'"�]�"""]��b��sM�bCDiCD�!"e ���BO߻.+�YGɭB�S�:��w�����)���幬3�:����uD��E�����X6���?묮��ggNY5PUt��xq몘~�LLj��:
\1i����]UYGɭ����S�:{��������ÿ:�u�_������������[w��O�&U���3����l�m�bƑ3�p�+�(p�$��{]�W����Ҙ��q����o�$�����Ne��׹8x������o6���������̩k�+t�xi˪�q�LL>}>�(  WZoG/D��ۋǏ�I"���GSs��ш8������e��|C�$�4n��uQ�UF ��dp�,�Xx���؞D�tDl+��z19p�3�P\���M#eeF"nJ���#§a c@�ߌ����Y��@�_�j�O=�u~�k�Ŏ�����KU�CSN���ߺ��*�?�'���J}���h���3-��F�u��i:~.���OG�z���{WDS>�����ß�?�c��/�n�ĎK���r��g�I�����ￚu�O���9ߔ~�����i�<M�_�����<II���w"����qI�3����:F���f~l��;.��w`h��O���o��~%�<��K��_�3%��;���Ӷ�M3҂��USNu�����(��\)�H�,�:�%�����MY� ���H_L#y��&ϗ/$��g��#�(lm]��čQHo�4�DĜ�s0������H�+D���g<�j�JN�<_�"��������&I��H7%�l�H'e� ���jc��eY�ȝ�s]��:�����߾�����yb�m��������O}�S[�����ZV���e-7NϜo���v�:
���I5��-˳��;�v��k��7�����D�u=�����WsJ����:=}r�q݂X�������뫫��[Vd#w�����Ϳ��?�롬󌖋����O�S[�O��ö9M���Y�_t��!^_�8V��v�Q  >�ވؕF�l!���&��g�l$#q���jD|7"�g�����$�H�M��
�Xf�LD�|��OӴ�X�䑗��q3�at%;wE�΋��+VT����w$I��Sr K����^C~$~״�G�ۻ~�?{������|��'"b����S˻k����o./�FwD�ܲ<��;�]}YG�Q��51TQ�:FnL;�~��l׿�����_��l]A����5�������=9o�ơ�Ώ�x���1���Q�ٓuU�߹&+u�����8>�\׿��g?�ˬ�\i����S�n��>�����'�6m*u~D�޸4�},�;t> 0f�DĎ4�BZz�|���?��K�=r�xD|����f�����;#��#�9Ӏ |,>�&�W#���䱲t�餭�;�|,��F�S��M�̙<8TښDzg$�]���# ��o��86�{�S�:O6���_���C�u��m�_<�FDܼ���-ko�����6�)/d+SC��vך��o�eF́��Ȃ��c�´�ζIg��֝`���n��z+"ny��.97��{�浬��'��c۝k��������}��Y����y�����lz'		�"E�����+`A��9^_�=���z<�
R�J��&A��FZB	)��y��^�}����9v��ٽ�~���|��~�\ܙ����N��y�<iY>G;�$4��w4t������w�v�T;�^���𴥻k�n
��<��ot�z�S�S�xJ�j�   �E�E�ak�#~"��in����'�֫���� %"׋��V�d��}�YkŬ�cD$�[ �,���QyJ�y g�wW�a�v�ɴ��ȝ�����Z�O,�?K�=SD��� ���T'���PW�742'��?k���r�mG߼�ey�����ƾ�����5--���.�-;WΗ%���S���V��˓��PW�?42;��������-ڎ����"r��qXOS����7-+癟�g�l_�@�ni�N
6����|���t���k���v���7�h���~�g�{Z���M+�y懋f�k,��/��N  ����yΊ<`l�~?�ޤ�h2"V��YyVD�b�ϯ����YF�۬�<�F ��ǂ;�Ȱ"i#v�y����vhH�����E�r;~�x>���Y"v��4(� P�~s�~2���3�xc�����w�f\��k�㕮������,{�}�_ܶ`���k����<s⁲`{��3Y�� ����V����ع;�n�=+vщ��7��SJ��q�&Y�ąg|�m�����ꪵ�����e�km�s,�۞[���T��|�x��kf�k�����{�|w�f��O��m��o�5��h7i���d��P�1f>  P�'b~d%��=dR�� ��J��ȣ"��xf���m̞iĞ)"�*� ~� \�"b�1"�{a�ш��������."�[���ܹG[�s��s��K `�uϪ��\����)ݛj�>m�w�ެ�Rʎ����?���O��yŜ�d���q�&)/�\y�e�`���je�A�;�g�{�u݃�N���[J��7n���'�pcӲ��w����W�3?!/�B{����?�V^9d�v�f��9���tǹ�޺���]+�;�ye7�G�����Ɵ���  �K�ِ�v}���!�ed�d+m���_���G��]Xacoc���E$�[ �w .�j��i��;yM\aDr�O��SV䟳��k��s��sx�  S�k�n�A�㹹�:�x�UwQ��k6n��r���<��pɬ�{fN��n�j�߸\�}a�T�k� ��|��~J�f��[ڿ|����v�+�lܘ��r�O߹���ų��U_��4ն�T�}~����2D��'$�X9��3�9��q�w���v�+�[�>'"�?�3��\P���F��ҡ�ȊgwJ]�v
  �0#X1w���O��4"9	C�2௫��\D.Z�`��˝#b���D�B� �O����U�V�W���0X��ϲ�W���Jm����0X`l�8�JD���  ����m�t�)���߶0ݻ����Y}��?Y��KM+^l~0��k�L�l�B�9� �`BZ��#�3�3�\S{���m��>1����o�vKӾ�w=Pn3?W�gN8P;��֥�%X2S;c��n��>1�߲�goK�:c�K��T��k��c1y�Df>  �=b�jcc���`��>�R�g�pLukk���08��f托���/�� ��p�;�R�#V���O�>eD��f�#b%�~RD�����\[�)yk�%b�,"��}  DA.�_�J;cJ�rV�oOߺ��w�o�X���iSF6�O^p��w-�w�Pm�l�Ki^1O��7ɬT�v
����[ԍ��`{��S�u�;���1�%'r�YO����w��󽡺ʲ���{0dNK�v
���1#�ZS^�1��\*y�{������uٜ���<����!�d��v�  �a�//��DC�Cf˖q� `2���v�BD�]�`iE>�Nk�]"��r D7�(5���]y�g{�s�t�a/��S��Q̦M�xl����^.;�Z�yT�� � ��a�N+�����%���v�]�a�x���G�[�y�Aw�v˔1"���_��+[^,�e4��2�E[�����og�����y�o�/���ݡ�2�~}�"F��s�\$����S��?9���G?�����٭]m�-Si�q�3� �DY��Q�\�e�g�a��d��r;�E��u�_��`{��\D�% &� J�b�^>7���� �;��>�H�n��`m���1b?/Fvhw ���W!/�B;c�4t��[��y��W��]�(:��m]��E���h�L��y�%X2S;�#�xL�?�|f����K��r�w�Z�%��gc�[�/���\�H�f�K�>��3�=����s�|���u�%7���2�g�K��9�  �-���/�s��t����Lg�v���g� ���P?�Z�6+�d��  *Xp��W�|Kl�p?���7L[�A�He:���/zA����1r���hw ���Y*�5	�)1#�i���\t��w���e��o_w�]G�x���X�<�_~s�*nw�^y��IjgL��aO�����_s��-Qv��M�uW���/��^,_/W{�����p�փ�P]�vƔ`�O��֯ϝz�]'����oVd�c��f��bC  �Uc"�6#v��$����-\���e�x"��+gy^|��yU� \ǂ;��g�W"�����~����No�N\`D��Jm��/^1O�|BD^�� �Te��l>r�vƔ�������]z�7�[��\�p��|��s^&�-��o��vG���W!/��vƔ�������}�^��_��\�p���i�g��l�g~��zٵ|�v�We�e�Ǝ��?�j�%���s�M>�ߋ�K�E���;�N�W���   �i����w:�w{a��)�� ��]��^~��������z�hw���� �ƨ�_�^����1��LKK��|CD�1>g�a�}H�\ "�q]!  {�Ö�h���1���~`ݷ�<���H1���y×��Ӄ����x�Շ��R�H�D~��z���2R�-����Ӿ�����%�g��}�iY�v�ƒQ�������b,C���7,��2xcǢm���֝�kw���7>x�O�sz�c��;�*�H_��ꕲxk �L�N  �����������HN;p��?��ؙ3ge��{����b�4 pF���P����y��l/��B�ہb���M~\�e�%�ȿZ��v  �r�|�>��ˊ,ږ����vh9�o�����K�E���Y��Z2K;��r1y�K�3&ݼ�w������Q�V���[���s*��=�{��$�t�v�g�cF��1�oi�"���?`�]�q�<x�gw�U54�Ů��Ҳ��5 P�:��/ecf�kA���v��LGG��.��`Y^�E�1�& p� &�cy�g{a��SW�;x�*0�Lgs�_��[k����n @˶U�"����}��wkw@����p�]oK��E����/��Y;�_(���^��������w<vϊ�Z�NG{�}33%j���e��R;cR-|-�uݕw�C�"���ȃK6���e� �(zQ�^����D:�תT*��Έ�ax�'ۘ9H�|WDF�� �T��������6f����d�o^��)d�lO�S��a�F������"��� `��-�G�&�E[������;𿎼��{�m�����xd���E3�{V�v�����7.Ӯ�T������z�v�ב�ڰ�]oO�Fw�-�.�s�3�?���h/�.��v�iW�����cn��}6������Ms�}�t�  05�"��o/+<����f�k�T�E?L]������"Ҫ� ��w ��m�|����ApA"�zA;���tz����"��"2�� �dk]:G���jgL��;�]w�o����:�և������D��Q_$�{RKfI_S�g��s����S�����?����xt�'�|83�%\4SzfN�Θ4�w�?~ڷ~�f���co��˷�^�e2�}��[� ��1{m>fV�a����F�l��47�����^C�21�>yY�	 J� &̊m�b��%Ka�󦭭S�	��W�����G=����/�H�v  ���#���53�y���ן�݁�l��_�����|4j^9O�ꪴ3������.c�l����U'jw�/[����]�e�c�h^�k߹2P_����(��Y���_��$��e�o��-K7��[Tg~��ّ~P �26 b��Y�ᇒ��k�A �<�e˸7xa�*/�l��v hc��Dlk>����D�����ѯ`Ϙ0�J��K�\v�o_sբ� @1�̜&��3&����Y͙C��f�Rw�-]�lK��ɐ���Ճkg ""��T'�3�3&ECGoUG�A�^zi4��"���e�[���6f��7,�� DDdwC��gjgL���������9痾�o|�K��ܬ�1�1���K�3  @�tX1_����0�XU��� �#b�ax����c��� �)���5o��`_?���47�j���>�S�{sf/11;��  (��]����1�7�_?�݂=s�w�?s���Hވ��A�$�+%��z�b�IQ98��vz��i�`Ϭ����ߖ~E�c2l;���Ұ��E"F����F���a��k�`������a����3� p�	D�G=�[�S����^�& ��S�08K�f��#,�(3|K`O�(F.����D:u���D�ٴ)㇩�9�V��E$�KX ��WȎ�hg]E.og��8o�uwqˎc�6�k����(��ꤤ����@��U�d�����X6/��߽�7k�`�,mi;bz{o�f�HUBZ����@���b��E�E��eގ�w���~ް蘪��GMo�ܛmG+}ٵ|�v  ��v#�x�,���7���?����[m.v��YDx�#����;���7V�[��    IDAT�08���$ �̦M?n���^%b�/"۵�  �[�+��X���(�����^{���jw`ﭼ�遹���K��E�!ᨾ-�صb��V��E���o�pÆ���{+�{z`������X�?�zp��ᖖ�sd�*��Qt_����~�݁��f������C��|  ��U���WU��S��T�7��ho���b�Pc�.�R ǂ;�?üd�9���ax/7�������0X)b>hD�) ���oX��PtsZ�^>��{�E�w�]�<����3j��J-�%CuU�(c[^��Pt3���\}�?iw`⎺k�/�oi�R�f~�x��Wkg��E���9���O���Ohw`⎼��oi������3dwC�v  ��:D�Ǽ���~^i�m�0u� x�����C��� �,,��}�b��^�:(�N��b;P��H�S��ꗊ5�H�v  Mc��ϛ��QT5#�U���hw�po����.����vG1Yc�U�3P��%=�I;���G3��Ǝ��@��t�C�_�-ܢ�QTFd��|��V%��EU50����o���-|�m�vGQ���w  Jؠ{�7:��SW���7?�K���b�hy\� ��w ""�"�^C�2?��ƈ䴃 ��e˸�N]㍎�k�|AD��  �sv����PT�Z����'_w�E��W��j��2�����ܱs�<�]Q<�Z�����]sWZ�ű(L_�;8��QLQ;k�;W�k�3�2oW�E�󣣾��i���Ŵs��H��  ��+�k��ŉ0������P:� ��'�b�yN� ��w�����2���0�M�eK�~xP<��gw"L]��sKE�7E$R�Y  �Em�jNs�/�^w�M�(���Yǲ�Z>ilt^��;�N��j�3P�v�@;���tn:�{���@��w�3݋_	?n�љ�����3s�v�Ў����5w��D���rԭ?ڽx[��X>��R4�U�5�^;  �./"�gcfy"L}�A�v��O����0+�]"�K� 
ł;P��b�fϋ/������sP;�L[[���9����� @D���N���3��jp4S32z�v��;�b���W�;�i����	(3����;#:3�rh,[��8C��w��j����bb�c��WI��팢��T����݁�;��GnY��}�vG11� (	?���a���T*Ў�#�O���^C��b��E�_�	 &�w��X1ۘ9��̮]����$�`�發9A�D�� �{�#v���]�]s��]���[��U�F�zǝ+���C��;Z;.=���۵;09�{�UFh�G��ҷs�|�]Q<��mfg�i��Y�bٹb^�>  �ż3r�'�a��v 7�-[��t�r/�[."W�Hd���|�����D�:5�J��] ���^�:B�\`D�9  �"J�VMm�����5�L�C��ؼ������?=Z�i��5G衊��}k�s;0y�kcj���F�b�����ѹM�/J3F�'�m���s���U��24�J:�4jg  Pn����{a��xlЎ������b�V������;}CV���i�x�ԏ�c D�������}��/�Șv �|�7�Jc�vFQ��y���{�v&_��m�޹{X��Xv-����21X_�*L�Jc[���|ǎ<����}���Ҳl�v��pm�tϪ��(�X�J]��{�;0��ܰ�c�����;��e��  �E^����s��A��-� &A"_I��3�ص"�v �	܁�b�&/�-K��K͖-��A �̈́�p"L]�7r�5�#� @yH�3S;�h�t���|D����M�2s��]��Q,A�>�(m�Kfi'֮͜�O�~�C��|f���mO�_�bI-a�S�uitf�ܖ�_��������3"vNk�'�j�Gj��| (aO���� ����uj� �>/�|�Pc�s"2�� �@4=g�秃Mgs�v����� 8=/�l1�C� mAD�cټ$GF������uf�ӫ�Q�se,�kg�Yv��奦w���:G������n�b�=MF��(����㹜��d8痑շ<t��;���̘&#5I�  "Ɋ��ȅ^��s�= ʋin����٘Y!Fn��c� ��w R�n�Q/���)� �-��{��ʊ����	 @�e�Ҿ�I;�(���|���}I�Sk�Ύ����m�Hz��D\�"&m�1�g��|f���u������H�|c$��7w`r�cF�E��lvs�S�_y7�~/3M����oD���x� ���W��#+� �ɰT
@QU*�Ap�{��l���?Ƃ;��3f??L}ӈ�{ @��'a�o��� b�� ������Whg,��ٺ���;0��X��U����bh݇�L���3$�ǵ3
��2�=_�S����}wNkW$^7���dk��$����l�Vr�/C����g���b`� PT�;�Ï�����1 �;^>���A�ʗ�������Z�6/�[��j� ���H�_���1r��D�} ��pI4nu���y���mء�M����n(�p	�/�\aD�0;�~��o߽U�:f�v��vC1��g��
DY���Hu?��7kw@GC���j7Cz���� @����K�08�O��Z; ��J�$����1s��<�� ",�.�Z1_���7�Nݥ ��~���s�����=  ��-h�N(��V������?;�G�;
5\����j�DX��,�[���3���������?��Q�Ѫ��7�jg ��L�N(��V���>��=������}���:���o:3 ��2"�eŮ���eF$�� K2�z���"�"���P�Xp\dd���щ0�i���(�����N?.���F$�� pS�����N;�`M���)W���v�;���V�bh���2JS֫��YӴ3
��ޛ>��{����;3�u�vG1��k�N@D�*b�=�A;�`3֓���g��5���;���9 �	�b�����°U; ���~~7S;��ܧ��|���%k�^�UVΫ� �.�J=Y%F��� pK���1�_�^�;p�v�-�����Ș���y,�`rt�n�|f~]�෵�o��ݟ��kw�eGL��������Um��7��/�:��ʡQ�oj��� �^�"d*b'��m�- P������7[#�H�v������@�xQl��D^b�mӎ�b0==�� �����"�M� ����Z98���c�"~��٭�[�;
���%JS����c����W�;�o��O�Ju���Q�(|.Q�:"��D��X�b���зf��љA�3���  �1ra"Ϊnm�c �XA���eW���- ��@����zsf�ӛ�c `2x���^f����6w �����3�z[s�ƬvJCc{���n(T��:K����������'λt��vJCS��E��廻�FF�������	�vs��������3��ZFj��  �4#�������[ `2���/���m���= ��@i{El�M^~�lڔю��d:;�t��F�:#h�  J����{|<�%���7������~[��S�]�����u�!�a�>qwC��펂��9�/"��tE�����]�����?����@��PQ8� 0I�Ś��08τa�v L�D����UF�~� �ǂ;P�����e�ӭ�֎�����q�;@�ު� (M�u�2��3
R�38�������@i����s�B��`��5\���J��P�74|���<�݁�2����s@��i�	��Ѫ�W�}Kt}���I���3���Ʈ�Οzf�i'  P�ˊ=�O�����d::ڽ08[�\("��= ��w��X�m��9���M{��v h0��}~�緯���� �����>�{�'�(=�}_�]Q��&�?�(-QX�m����vJOc������P��g����G�Pzj3_0y��~�Lf>  �gԈ���S�°U; ��ApS.�=H�<�� �XpJ����O���R���9���" �����KE.������{rôށq�B���b��m������(=�ܳqcC���vG!���!JKf~,o��݀�s�m>W�=����Qx  �"y����^��̈�c @[e{�N/L�h�^*"9� �;PFĚ��a�v��ܧ ��2[�0�ƈ�DD2�=  }�/SU�����=�;P�;��h7���V�1�nB��:�LU94�Y�kw�4�w����P�ݍ5��3�Q<�?(W502~�w�zZ����{`�vC!�%�ŵ3  �e�fO�����) PJ�H��/H̬1;�{ D�>��K6f���)n������0u�9� \_p��=��3&Wm������b�?�F;�;�����ݯ#V����g��B�c1����������v��݀�U58|�vC!�1���9 P������Ap�	�a� (U~*�K/�""?�n,��̷=?~X"��o �~���F�=�-  6fd���ի�F��n@��<pU<��[<w7��E	1"����{�y@���>�:>���ʘ�(�ݮ��G���n@�J��ucb,��Co����	  L=#Od���P��bv�����"�EdT���Xpt�[k����?��f�c {��R=^�z������k�  ��pm��cF;c�H6oo��@�Z���4thwb`Z�v"b�:)���__�<����h��O4v�kwb`Z�v"b�*!?��1qV$f>���7m�L����(�| @��[1_�प Hi� �k�0���̑"�U������p�s��9<�Nq� �S����٩� �:���^��=����o�����W�
1Ȳ#�d��KTU#�~�N�?Ϙ|���[�
1X����c��s~�S���U���z��s���V��  �T��͙�0�y#���@Q"�z�;\Dx�	a��R滞��L��i� @���&��7Z�?�n L�!�gk��Yn��T�?��vC!_JF�r|���ox�vJ_��ч�
1X������s~M����������� (�̉=4ޖ��v D������b�"����܁�1*�|�S���Q� ��~�n�\"ܢ  ����������(}�ãh7b���d���o�N�;}K+�F]��{�
1����c�����k��>/g��]1q��i ����5^C�q�aآ� QbD���!��ji���܁ɷ��̑~:u�v D��^��̈=MD��{  �g�����O�P��p�OQ92�����j�]�(t|ٱ"�yZ��o�G~�|��X^�c��U�5}��Y����ێ��G���Ѭv�D�UJ>�O� �H�b����f˖q� �*���W^>w��<���|L&#Ox��щT�� (^>�{��٤� �#�	턂�T�N�̍�aD�=����*d���3#5n�|�{�k'��[�?ԯ�1Q�XL�*}�D����|+���ޠ�7��r�r�|,&��| @�������k� @90mm�^��b/�nP�Xp&��5/N2mm��- PN�°��e�7"�[  ���鉑��Y��>����#�vC!XvD1�&��;��2����s�vܐq�|��G1��wT9<�=���۵;����x�vC!\�� �g��{��n��v �#�K��%b�"2���t��ߨyo"L}ʈ�c �����x�݈�D�� )�����X986�� w$F�wi7��QP:F�ܝ�U��C�pGb,Ӭ�Pf>���s~rh��7�`�Ud2N? �� D��k�9�י0��N�r���"�M"���! &�@q���կ� �ɈX/L]���E��׽ ��X��?�'��y��X"�}U��./��t�|Chrt�[��H�����P�1f>��噟�p����m�n(3 cb�~\l6m�h� @����Y/�%"Ok� (=,��b�/���o�S  �+�J=h�7��oG ��*b�����e���{^��./��4�c1�=�	��2�v��d��n(���`Fd<������V��Ì��Z���� ��4bO��B (-���ͫ�<I�ܢ��������C��5���M� �mm/y"G��'�[  ����\�eG�xF������+�%=�]1q�L>�� wxC#�h7���B�%<������d8�c�y�8�֎Q�ߪ ({���!7@	2۶��Ap�X�q�k� (�~c�{E<�݄�v	 �/3A��UV�*Vn�n LL��|ED$cYv���޹M�v��e|w߶�Ґ�+�
�	3{l�kۍuw�g=�?����[�DD�9˂;����5�wwW���+ �l=���� ت ���t�rk��"� ܁����0����1 p�ٶm�O��/ �)s�*_�I6�n�;f�rs�?��Θ0[�����n/̚\�eG��;�cg7�]��B_��ퟪ*�6�� ��#g���s� ���5ޜ�g���>� ��I���j#¿��2������^cc��A�-� � ?��܊9_DƵ[  {.w{y�X�m��cF$�:���s|Q�\��ۦ� �0�Q�\_p�Z�Ԅ��gs�>��� 8$o�|���ͦM��� ʕ�em�yY���� ��	��/��S� ��%��m��:��n ��H�V����x޺��s�����ݞ��|~H�n�����|n�E�\?�W�<�|���9;��� n�b���࿴C  W�N����E,;z@�r�[C`�ٜ{��k�  
���6_�ZDZ�[  [���|��a����rV�a��/'C��I+�|�
��]�}�r1���Ɠ��|�X�ݙ��C� ��0`Ğ�S�i�  
gZZz���SD��- ��B {�q/�8�*Y��I��l�TĎ^���������fG�X��&���X����Y�`�c���+�>�A���UX���^1�f�&�s> ��Y��9�Ç�[  �c�m����V�W�[ L-�� ����k�_gv���. _ukk��+ֈ�'�[  ѕ7�_M�)����"�z=P(s��#��`���*,3e�0� %˼�{��i�  �ψ�D���s��mP6�q�[�|�S�1[��k�  &�믶J�5b��n �y����Y��H>���n�[l�8{%nE��Q�X��ˬ_7���N�[l���*�n�Ѡ/�u{�g�1f>��5&��0Q1�� ��d6y��	Uaت] �\^��L��WD�}3�=����T�b/������a ��m�X<���[  �"���6^��;����p�6P�ՠ���Yk������pw���R��"��ߐ?:���^ɻ�P�| @�1�7:|�ik��N L?n�b�NDF�[ L.g�@&�5F>��K�C  Sˈd�0���\�� �C�/O�s���%3�~o��r2���<�q�/�N��w�ځB�~�ϙ�|��pv��8� J�s��y�LO�n� ��J�����""C�- &��_� �('�\��i�  t���`�� ��X��ҭ���p��e����۸��}1���ab2G�nOx���G�\���<��e܏{��� �{k|άsMs3��@��ҭI>�FD��[ Lg(&I�y��N]� �煩�Xr����������pǮc�����f�����~�)�`�c����!�pw��y�>��%c�c��K%6�;� ��o� D�U^�o6m�h�  t�m��#'�H�v��s�`�[kޑ�;�C  ��S����� @�?����X�l�����v�vC!��v獻�0k���� w��Y��5F;c���?�����!_��c���<?_��̯p��j ���/��� �� xΊ=ֈ��- ��w�ucy��H��� �?���, U�ȸvBAr^|�v�1��Wh7"9:�� �%F��Xw��y�eG��@�G�    IDAT��J�B$��>�A�?��X��[���
���c#���
�� �c�|�O�r; ��%��ؓXr��w�����ax�v �t�a�m�!q�W p\E./�÷����y�pG&Yq�vC!,;�@&o�sw����cc��vC!XvD��H��Y3^|�vܑ�+�n(5 �X1_I��Oiw  JW"_��ǈ���- ��w��a#��dާ (}~��N�|@Dx/ (qy�e,�7i7��~���YvD�<��+���pG�����g��忣�Jo�vܑ�ܾ�=�9 ����b"L}F� P�*��w�s��Ed�v�±��r6jľ��G�C  ����1r�p�; �H��{��hM�F��Kz�
�p���ґtx�q�:Y�� w�'����H���YE�p��_���n�;2	o�vC!��~V n�"��S���  �#�޲#�ˮ�V� �a��j<f�\�� ��"��; L9�ovM��|�\���1uF���
��g��忣�D<��ߺ�v�0\����P��0���p��3�:����7�T%k7"9��g � +_O���ig  �S�޾33'�P��ı��r�ɋ=7h�  ����Ě���n�rR94��P�����(}V�b�����㙜�����U�j'�����(}V�4TM��\��|QU���k�����#��*�k7LT,o�~  �#�����hg  ܕL��匬�"i� Â;�MΊ=?��i�  ��S׊5��� �rR����K֫8N���7��Ѥo�;&���G Q5���
���c�P�^<�CG��������b,C�s�����݀���w��h���B�c��w�H,�- S�~��֮  �/[��5Vl�v��ǂ;�I�yW"� �?��܈�D� �EmߐvBAƪo�n@��N:}��n�?�(�}n/��Uyi7��Ψ=[�����P:\�[K��j7��zr�8�H�H�| �T�r��3\�  (�d�j�Y'"=�- ��(V�|8wh�  ��S�Y#��� �f��eǁ��%�(}�uU'k7���5��op�o�Y�݀�7T㟢�P��~�?�(5n����n@��L�� +�| ����y��Xn ��K̜&"��- ��(F�g�0u�v  �A�Y1r�v D����V&��m˵;P��Vh7��D;���#�I���@��������
���((5Ο�]t����<X��՜� �����}F$� �&?�z�y���j� �3,�#�/{a�U� @�yA��"�}� ������ݾ�'f3�k7�t�v�!3���j�;
Q���R2JG��ĳ9팂Č�[��k�ɇM�Q[��Q�>D�H���7��Θ8#Rab���m9w��7�v�vG!�8� &���3o6[��k�  ����Xk�-"n��	�uW%���#  ����9�/�"�[  �L�J]πvFAF�+��n@��7���
팂L���(+R����Pu��(]]3�>���������eZ��˳#5ɷh7�t�T-~���Bp� L��x�-&��U! �)�H��+��o�� �0s���] (/fӦ�/�<yJ� ���s�vBAz�j��n@�h�>G������(-n�����֊��l�<�uU�j7"��˴n�Q<�}�	�^�J��k�2��[]L�ʴ.��e �����eך��^� @y�����ȧ�; �u,�#����׈�C  �Ǆ��8[ļ�� Q��ٯ�P������<I���wƴ��
1�{@by�)��i�r|�W������(M�Muh7��gH*r�|O����T��|�-'hw�4�M�9L��u}���3  bŶ�r�u���C� P�� �/��u� �#�=��;�e˸v
 �|����lLN�V� ��op�'�n@����ǝ������(Dc����(=�?�$"���?�݀ҳ�'��^���(3���[;DDr�Oh7��<��uo�o����(D>� ��2`DΨloߩ (o^:���Y���ǂ;"ň��֞n���~�)  �R���b���]�"r�fG��uk�Pzzf5~R��PQx �%
�T=3��n@��^�)1��ip�(=Qx���iډ�(=�Չ�Y���� (����s�0��v  F�z���ȣ�- ��|̜^�ܔ (����&f�*"c�- ջ�%1���(�@}u��:�%w���9ӎ�n(TC�/(���QI�}��V�����8U���{V�j�BE����ȸT�jg�����ы�|�vJK��|h�& @qX{��n}H; ��1[��{�#o��[ �!�����J�R/j�  �ǼTj���"��- M�^턂e|��(�:����k}�Bk�)ݣ�����?ZS��P:�}���ΨMhwĊ�hs����3#t��*��N���g�X{RoS]�vG�8� ���7?���  ������Y�g�@���b�Q`�5���'�C  �K��-V��;  *f��	��x�㗞��@i�3��B�w8�v��H����<����^hF�t̞���봞�߮��4+
3v㉜��;���_�]Q�ھ!�d� 
d�&/��� �_R��V�Y"2���u,��yV̿'ҩ[�;  �[�0�{�v D�����/#Չx>5�����Y�5�-���vG���Di��r�����DEb�s�An�1�4�-l:P��PQXBFi����HM"nS5���O8!�9����� (�����iG  ��a�l���E$���w��~��T; �=aD�����ϵ[ �uMm���3
�?��#���6}������:��Y|������X����ײ��?G+����W;5��O*����k?�� }fq�G����� (�vO�[Ͷm� ��xl0b��v ��4���~#b�K  �S��y�{��l�n �y�Yi����(X��ƹ_����;�Ǌ����x�vG1D�m��x6'����3
�5�a֣<�L��"�m^����0+ե������������s��y�]t։���9������9 0qf����b@  ���W����@�c��j�2�3Mk�  ��Lv�\�-"f�v �lv~d7"�U��kg@���qʿ�6�%�;
U58*5}C����Y����L�z�yש��9�R��P�C�R�7������ۢ��pm%��2��g|�gf]�vG��#�2�{@; ব���%�[7k�  0���+�;�rƂ;\4,b�b:�۴C  ��D{����#"�w �̍�?	��M?��|����1�����0og4>�(]swvh'EǼ����g�����Oi7�ܝ��S�jns�vBQt̟~��m�vttϨ�T���6���} �D�����
  &�lڔ�b�w"f�vP�Xp�s�؋�0|V� �B%��~c�R� p��n�gr���c2�n�������O�x���z�b��=��(]�[���jg,��pM%3����k/j�;}�vG1����c���A����ي
3��1��Г�=���y��hw3 0!Fn����  �A���[D�W�
Xp�S���$��v�  �%_�;�; �E�lNf�vkgE����?���;0�R���;��������T��]�t�;�=�=�� q�} 7@Ddqt�.��uf�q�]Y�MP��=@���=�����}߫�����Ȗ��?U���s�'O�鼽}��~���nH�pT��f;.�I$T�莟���)�W�r�i�;0�"Ӌ�%c����Q�A^j���$*�w��Y���\�g�����f�׹�� 0������v  ���;�����!0�XpG�p�<폄�l� �d2��Eo��]�[  U�5�NH��ף��=�;0~�����QV�g�#�#�
Gmg L�q�	�	�G�99��݁���/�|kya��d��ܭ���� Sk]2��g�L���Kol�(,�ݑ�-���� H#����\nB�!�-  $S�)��#�[�;�LÂ;҄��K�i�v	  �f���G��$��n�t3��';JRS�E����R�{�_h�U���RQ�4���u.��ӧ���+�o�c�j�b_Ü���vG�T�d��oj]�k�Ek�Vt�.��vƞs�<MS�k�#Y*�� �����P0
� `,�#�/;����dܑ��0�K  ��in��$��$%l� @:���פ�^�I�x���~e�c/\깧�(/�vG�L;��/) �M�Pak�팤p�Q[q��mw`���X��������x	�iJK�팤p<F]%�8�=�i����E���J�$U2� GĹ��Ը�v  c�H	�/�Z���n2�H}F�B��3  k���r��7mw @���/b;!i�K&�<s��j�cg�eg�=8�|��d��ޫ�6w�d��0c�{��,ʟ���+]s�7^o�g�h�W�Q�ɒ�կ�.Y8Fz���=3����d��W|�v��9��qv�;�eb���43� ����?���
  ƚih�3�LҰ� ������g�p��  �S����
� �Nf�	�NH����V~�#%�;06�g�,�	��2�E�gH��4�NH���)_~���*lw`l4WNyj(7�5���vͅ�7kO��خH���⯭���\�T��IO�fg��H��{C��� S�|Ѩk^� �����6�ѝ�;�L����p��}Y泶#  OFJ�Gc��� 8L��}*hw�	�C��I<n����G.��3Kf��H��.:M�ab���N�fg��>a���Ͽ�qV�q�;��M_P@z��RQs�팤�x�'f3�]h�G/�xxV�B��4s/�& ���I�^e���l�  0��M�I��v�v,�#Uu%F��2�А�  ƛiii��K��n�t1c���"ӧ���Ko�݁��}ՅeuǕC�9�]*h�U~�/1�f�l�*2��5���6�H��/xWq��S������>���B��.�r@dZ��go\�I�H����ˏ�-�?�㞙��կ��� �4�ȹ9�ܼ�v  6�F��h����XpG*rr>���Pk;  [|��Fc�E� �.f����1j�Q��n���v���b⺾I�^��4kO��d�Y{#���2RÌ����USm� 9�s���M����H�Y.[2F���/,�g�;�(2��'\�Gk`�Ꞃ	ٶ;��� 8L?	D"�ێ  ���2�p�H����H=F?̎D�� �m�p�{F���0�u��4�a;#�'d�:&������p���k�]:�vG2y	���`;jBπ��lg$�Є���0{�����\���9e���H&�8����;�}C��s���:�=�]ɗg�.�ݑT�4��| ��1������  ���Hd������H5[}99_� @*0��M�~�H�- ��m����t��g��������{�s�w������H�������@��r�턤k-/���������M���ꓦY�vIrUԵ*�g�v2�[�������[w텧�W�u����M��� Hm�N"�A
�  ���et����XpG*p�|�80b; �Ta��۔0�4j� R݌}a���3���ܒ�W}�����۷t�ʟ	�]��"���b����#�t�-����7�����lw��m���Ig�>5�����b����
��ź�9�����������yi�eZ��`�u�Y�|�v  �9�hj�c� �T�Fo���v�6���4ftG �k; �T�k�u���v ���xB�w5��H��ף���V���[p��TϜ�bWQ~��d�����v2�'�М]�3�.�e�<��׫o�|���p唗��&mw$[�DS4��@��$���}34ˣМ�{���Y�[pd��:���lw$[����h�� Hm�#�_َ   ՘��~9�k%��$.�"ܑ*�ÿ� @���_���� Hu�\z����l_[yі՟:{���U����𬒙�;�¼��$�3 ��~PrlW$�Є���tR�37/˷݂ó�ƥ��g���9��I��/�μ�������پ���*����37_���ғlw���;�� ��F���f; �T�oj�2r��v�&,�#��d; �Tf���h�ZI}�[  �������vƘ�*�/��m�뮻�]>ŭ����,�<�v�X�$��Vo;�$�w�����vƘ�,�������O}���[L��v�X�$:~[��@�4�{@�u���@WQ~Awn����Է��|�������&���mu�3  �k����	�:m�  �ʼ���HZi�pn����񘏛��^�!  �����:ɹ�v ��/��0fZ�N�}z׮ն;���ȅwV�2�ӎ1�S�Ĭ=������jAU��1�R1e��={�����{�o߻p��8w��������������g�޵{������\z}͂i_Mx��hu���&v��  �(Gη}��F�  �:#9q�$u�n���wa�N����؎   ]�#�_G�� ����Y����mhf�YO~z�c�;�z/}����/��ݸ7�vʘY�{ː�*�ZT��c;c̄���ۯZa����G/�f���4�s��?����HOem*j1fB3�߽�����݁�[s��K�N������7�$��R�� @���/(���  �E092��� ܀w�c����}�v  �ƛ��.��v �,GZP���%K���������l����v-�y�H��ڥ�/#}�}��[~��ۯz�v�f�G.�r�I��	�];���4�����z�|�7�)��������͆k/9���������jiC������ ���8�1�kW�v  �$	�^���ȵ7c��bJxn0��öC  H7���5!�&� ��f�jTp�ݿn�S��'�iٟlw@�pͅݳp�#��]t�8��k��F����Ss�?���z�v�M8g���=2�p����|��f�(�g�vƘ:8��O~�O����]Z{B��`���S9� �f�ѿB��;  HG>��VI��;�t��2H]��]���*�  ���H�1���v ���ф�W���s�Y%W<��e�mwd���\���Sf�7��w�=�)�ݪ8�d��<	'#^��(:���,[i�#�m����>����lW����Uֵ�� ސ'��I0�g�^��?-��&��^{�5�g?6���e�e,������v  %9����lW  ��L}}�q<7Irl� ���7⑪�*oS�[�+  Hw�l���� ��-��q�)��]r�_>��M��:�k�%Ӭ���سp��F�>W��+I�6��,R�q�������Yr�_>���?��f��L��c}u��?	�柺a3)m��u��r�$�f�����~�������K?_{�{G�}���� �����s���C  Hg��Ƨ%������3H9Q������C  Hw���Grn�� �ycq��)3>��^|F����u7,+�ݒ)�|����.��Q�������Z�I�Hm���Nya��q�^t�ƕ����vK�Xu��ݻp�]1����'7w����v�F:�}�3�Ed��ŝ���o}��L���W�d��3��	/�Nn�Ҵ� �T�/g�B��l  ��7<�9I��;�tĂ;ƕ1�z �a�  ��E"+%�c� RU���+I��J��kV}�Sl���s˖�,���m���p�Um�c;8,�^�Sn��q�^ZP�^^p`��KO���f��	,����S�]��~�Q�t*_�@����^�lg���҂���f�ت�y�o��Wo��?��DVf��E�� xc}M�َ  �-Lgg���6�@:ʌ'�H/{KK��v  n��|�Ha� ����Q��|f��(Iݓ'N<8�b�37-���7����7���e�K%��l����фNy!sf~O��	���_Z}�埱��F�>t�'�i8�l���r������K    IDAT3���I8Z�A���������8Xp|�anٻm����H�*�J ��F����FJ� �M���r8�8R,�c��d�q�ys�v  ncjk{r�� �j��zM̐�%)���ԝ0��o���w�u��'Ɇk/�cω�w���n7�tښ��+�#2w�A�w���7#�>O�	�����{�eY�{�b�u�ܺ�䙻��m����� �ٻ5���vƸa揍��������eŶ[���u�l'  R���o��f~1  `���g9Ͷ;�tn��ѷ���6�  �U ����lw @*�M�ՙ���x�斾A��y��W�d�'��>���o�r��Sg�h07�Q�D�w7�8�i;8"����We��o�]�T;��O�veƜ6>�/�Xy����Y4��s�3j���RI��vpD<���<��vƸ���w�紭����l����g��]�ɥ��_8뷃���{�ӌ}a�60� ���%o$�]�  ��	�:�x8�8,�c<�g�o؎  ��|>�mw @*�VQYC��q�Y�_T;�t��ۮ���t���_���ʶ����x��q��u�:"MU�6����vƸ�<�02���gny��m����:��m���V�`�y�L���Q������T~�M�5�w�Y����Ь�M+n��;�[��s�]���wW��?q�҄'��f��| ����j�Q�!  �Y�)�#=n�H�u�V9�2�А�  ��<�$9�j� R�;Vn�'���1���温_z��D��x�"�=����7_���S�>�U�?�v�'m�V��_呾���.O±�1�������?�k�����?��>;�ٛ�xt�i���,Οh�ǆ_�VnϠ��-yv��F3�:?�zꎟ��G�pmӺ���j�'<�l�ŭW>���;��'��ᤗ�kB��� @�q�$��v  � !�vI��;�t��;Ƙ�;_$��
  2�/���lw @*��ޫy��ΰ���������O}�V��ٶ{R���]����S:��O�xԛ��Mr{u�ն3�c��ѧ���ΰ��lRi�����?�����on����S�Y3�,�|���k;Ǌ`��N���Gz��=����ΰ��lR遹UO�~����=�j�KoI���Uw��ƽ���T�+r��u"3 �z��x���#  �9�H���5�@:��'�/]�x�s�#  �$FJ8s���� HE���V����kb>�98��C�Y��goZ��=�d�'���O��у�O��?��r�{lz������"5�������5�J?��ս��+�l�'�l��e��ӿ|�~��Y?�-���/ ,Y�]�X�vp�NٰG��a���|^spn�ձ��ݫn\�C��������>R����?�)���cӒ�;�2� �����ik�Y  Ƒ7�����;�Tǂ;Ǝc�`Z[[lg  �i��G���;  eE�d�v����L������]�I�=6U-;�����f~�����i�{l��/�i��lg I�iɳ/�ΰ�bN�f~�7���:W�z�-�{lڲ���+>u�K{�O{��b�t�=�Uֶh�ް� )�Ѹ��4υ���ꓦ���_�X�[.��v�M�>to����'Tnj��<Kyf��L�m��=!� �cd��D�l� �Lc��<�6I	�-@*c�c�_S藶#  �T����$5�� �T4kwH����+I]S�
�+��#_���ٛ�������K/��������^w\��Q/�H�#1�c%��p��V�K��=%����ʟ��K׵����m���?z���_��3��W~3���gnSYӬ�yiCze�0����u���t�M�{����.=q�W=����{��-�f�N��e� ��`\��؎   S�C�Mr��@*���+%�1�1�c; �LeZZF�����<`� R�;WlS�'�Q�ﳝ��K'���N�̓�~���[z~y�)�����1�]ca��\֓7�?�UN9���:}�N�mg I����<m��f�$u��w�������Z{~������-������0�_k��
��� �n�ʗ�4�X#��|I�,�/�,���������t�z毽��s��s��gF�),����u{��� �c��9�H��  2�/�|9�p��4�v��XpG���
�h; �L�D��W�"�}�[  ����������Sl�����'����O]�&g$������������]Z0���G���kv�M�ݓ�J�5o{��`L��x�.=�B�))�g��ܞ�����c��W���~�_�i��c�����=�z��kv���.J=%����v0&��#:m�Nm�h�픔�[8!��p���;��qպ�X����cU����ӟ� W��_�-�x�ޢ�"f��G:u��Z� �TcT����c; �LgB��hy�W%�[�TĂ;����8�j;  �z��d%���> x��ԩqN�"Ӌl����	��y�������m��=���Ĭo\�퇛m�����z�e������~�.o�?әOm�;lp��_�S��r�g�NI9Cކ�e�ǩ�×�m��5�����~����n;\U7/��EK>�?)������1f���E�:��2C�5oG�斩qv�픔3��6�)?�8�K�|��	��z��q�O�n;\��:��i�pK_^�-����S�DǛ�Ƙ� �7�p�;M}=��  �"����+n��	-�?0��
�j ��;��o �B�ߓ�;mw c�s�����7lg���G���v�����	����j8�o;%�y	���'t<�Q֏���#)w�����_<��181���҂Fr�,������읍�3R�o�V�(5_|q�nU����3��`n��|�9l��<O"��-=�	݃Ogy͏���G��n�G�n��(��}07pug��sY����{�o����3R��@���c;�9��+����HyC���|�9�Ͷ���<��&��4M�X!g�������ݸ�pD#��������������h����3���W�̛g;�9�����=�3 �!�ѓ���;  �������Ȭ��6��XpG2m�E§i�v  �g֬����>I%�[��Ă;���y�Zu��igb��P^W���Pt�|�{����;ƻa�ˊf躡�����&�&���w$f�i�{��r;LV���n�sʴ�w��H;z��v�FW{��s~�Ǘǻa�ˊ��6���??waWQ�䄇���Č�a��O/��H,��ChV����]<>Bz���GV�u��[���B����`�e�����f1������M�3�&Xp`�H�cN���m�  �׊VT�+G��� R��v ���3��  �S[�-��o2��m� @*��?�y�����S�J_~nN_~�i�N���{�qS<�o�-8���U9�����_�"���z�S�&Ƣ�0r��f-f���.�;1��x�X:Z�=�z���lg ��@���V��g�NI+��������J:U�����M�	}Cmك#�ޑX��FJ'=��������Ч�M�4[�u���Y���N�.ߛ���?��!��)f>2�����R�݋g�NI+�y�����"I�$��=߼)�j����D7{b���r����'��r��`N�,�8zG��}�H���Ĝ�Ƽ�`b:�4�`����T�}p �~�r;  �)n���s���� U����0�c�px��  ��|M�_��+>-�$�- ���X�C-S'��p�픴5����$�Iz�_���߾�����マ�h�7��&�nGRV|t !3�qF}	o��x<�qr�ެIq�wb�����]�@V��3w�$z�U�G�S�qw��j�:Y�S�l�����g����:����7���G��F�INV,>�0����|o��7+/�g��pt��U
Gm� �;�4}����Gm(��R��3%�)I��έN�?:��y����X�ǛP��a�z��2&�g�H�?'x5�꿞�0� o����}�v  xc�P(<R^�?F�7�-@�`��O$F�d;  �9#�ƌ�t=k� R�/׹�n��׽Wр�v���|^+�u�ĉ)�{p�ikv�$�a;��չܤ�\�>E��M����%M��I���VYc�����xB�>����}\�'Y��5��^3�N]�Kem�3  )�|���wۮ   o��~+���:X�x�p��@s�n�  ����U���mw @����әOn��%�ؚ�7�Ulg V�u��ǫ��p�i�M:����3 �&v�ǫd�>�mZu�N~��v  5��
�f;  �5���od��v�*XpǱ��ţ|�
 �t�8���� �jZuD'V� ����ӻ��f;H	��t�&�^y]�:�	^� $���Y�<��v0f�� ������ٵ+j�  �=_$�kI[mw ��w#����b�  �@S����� He��ݥ��V�@���1���M��l� )����5�����E�:��/���f�nܫ�Zg�}�� ���D"�]  ��F�mw ��w5#E���v  82>�㮝mw @�2	Gg��%�u��N��$������賝��8:�������q���fMj���{�9t�_��k;Hf> ��cX�  ��"������Ƃ;��#�U
��   G�<������ He�CQ]��s���$Œg���@�� %�����+���8c�vM���� R�$��yA9öS��`� ފ���/~�v  8
�狒��M,��hU�"��ڎ   G������N� ��&v�?mRV<a;8&'mگ���� Rڄ����s��Fm� �dA������ʄ�������S�c�� ���c��ڎ   G���Xe��h���w��+F��/  i���wG�c� R]I�Cg=Y%�p@�ӌ�a-^��v��4u��'63�*k�u����3��0��Kg��%�3鉙 x[����/��   Go�q�,v4��Xp������`;  o"�GN�� Hu3��u��]�3�#V�Ю3gY83��u���3�#V��ُ�Ȳ.p*k���g��� �3 pb�D��lG  �c���t����q�<	�E#%lw  �ccZZ��� �N|�Z��k;8lE�]:��䍏�N����-ڰ�vp�
[{t�#��c�G����:cK�H�| ��1?�ni��]  ��hb�k�Flw 6���#���9��v  H_A��%�� �`ц=:i�~���*h��y?'_4f;H[�۫�_`�#��w�邇�S`���U5Z�</�"�1� �i8��ڎ   ɑ��\/�׶; Xp�1r��   ������o�� �tqں]:~[���M�u�낇6({(j;H{���҉Ulg ojb��.~`�r�m� io��=:�E^lB�b� ��`(�]  �'.�?�)��@,��H���DV؎   ��e��� H��g^��|��'��_?�A�~�q�r����r���u&v��7(��EG YN[�K�o����3 pF��p�  .�D��7�;��Ƃ;�q��l7  ��3�8r��v ��8z�S[����v
���>]r�z��l� ��H�^���ܑR��u������#�s��:��j�%���� �#c~�9�  �盒�|/2
�8Lf��)���
  06|��/��'+�p9���k�s{m� ��ҭK~�����H��ڡ�kw�.�|^hƎ#��f'3)�� 8B�Qg�;�#  ��F"�2���`<�������ߍ���   c��)�|� �Ԣ{X~�U%�]t�zeqh0�N�T�̇US��u�C�=8b;p��7U�+��T�0� G�9MMmG  ��3�8���#����ñ�
=i;  �-���sI-�;  ݜ��ZK�}Y&���Wem�.x�9��q�)@�8yS�޹b3�njm�.z����t�{�Vy	�)�0�| �Q��:	1 ��r"���g�/,��m9F�m�  �=S_?l��v ����kuޣ����NA������yt��1�ہ�v��:�����0�1>��׹�>'/4�n���:���y�㆙ 8*����v  2CB�oI�m|d��֌j���#�3  �����XR�� HGSk[u���+�7d;n�H�6�ѻ���i��Eu-�������Xze�g�Vy�j `M��V]�����7c� ���$<߶  �Gv$���<f�,��%�-#���   ��tv�:2?�� 骰�GK�]��V�B�e�:��p�^�) $��j�k4���v
\(k4��>��REA[�.�w�&7w�N�1� ��H�Zw��   ����?m7 �w��_���v  _������mw @�
��߯��}�)p�ܾ!]��u��'d;��������׌}a�)p�`ߐ.��f�f��$80��ؠ�{����a� ���߶  ���B/�h��`����7ed�oB!�� @�1m�͒s�� Hg�hL�<�I������8FemZz�jqb(��|Ѹ��؋Z�j�<�|�҆v]~�E:m� x�h\g?��޵b+3ǌ� H�|��F�  `�yF/���XpǛ����?�  �HHߑēZ 8�t�j]����خA:����C�R�#ͯ�х�W� C�Qp���k�|~���wܶz]����F�Q`� �đ�_�  �Y͡�$���%��&�_���n�  ���Hd��h�� p���v-�w���8}�/{(��}��  i���CK�Y��p�����pL���-yv�<��� ��$Ԯ���RI��v
�3 �<���<n�  �a$Gr~`�K,��8	�'�#  �]�|�v �EnϠ.��:-ڸ�ee����6]�gUY�d;�Q���%����;�a��m�5����<�i���@:
����7h�*������ �$���FmG   {|��}�Zlw c�w���ώD���   v�"�g$m�� n�I$�p�^]��u��=`;)ȓp�h�]��F��m� 8&���Mպ侵�|�!O"qh�?�Q��!�9 ��qͯ�ѥ�[���~�9HA�| ���e��  �2�82?�����zF|�  ����v �MQ�S��v�f�n�����ѧ��]����8���EQs�.�{���j�����٧K�[{h�s�?�S��u�ݫ5wG���f> `L8�����  ����W�&��Xp�k��ëlg  ���f�+>i I����ǫt��Wn��X�I$t�j]q�*Mn鶝`�Gb:��:��)�����<���o���w�єff>�F�h\�Y�Uݿ���33 0�	��mG  ��`ZZZ��!��X`���0?4GH   I�|���/mw �[U�6�_=��7Usjw��ҭ��]��kw*+���`�M�m�U�^yh�s�k�)l�ѥ��Ւg�����0���u�oW1�33 0���_�klw  �b��N Ƃ�v RJ�/���  �ZF��3��%e�n 7���Z�v���4iㅋ�3y��$�1_4�S7��	[jYx2�76��kw��:�����)�|����Z�~�l�a��3���6^|�����N�c� �G�'�  @j�G"[���$-��$��;�ݦ�e�v  H-�H�1V^�#-�� nV�Е�yV�'Oז3h8�o;	��H3��u�����]���H����*U�<M[�3_����$$�_g�����a�����K��v53�͘� ��S�DVڎ   )��rXp�����W9	��m7  ��d<�N�a� Ƙ'��m���7�m�>^{�T�㱝�$��ԭ%���8�a;@��$�|���ܥ%��P	3�+�6��ڹ�8�<}63�%�� ��d���H	�   ���y0�8�#��v�,,��Gk��lg  �Ԕ
=�(�Z'93m� @&G���횷�^/�s�"Ӌm'�(���u�5kO��خ���~�t��
�,�������u�5gw3�
Ǵx�N��ՠ��>Q�Y��t�� X0���v  HM&�VT�#Gw�n��w�Z#�    IDATH����v  H]FJ����7m� @&)h�ՅnTK�dm=�5M+���Ô38��/Uk��e�9X��+h��?�֊�������Oك#Z�R��o��7>j;@��ޫ���Z����ǩqv��$&f> ���MKK��  ����S��g$�-@2��Ij��Q���  �¼���bY޻$�-� @�)	w�6�e�dm9s��+'�N��j���YxpԊ����C3���T9�v�ī3K��1f>�#W��y�<h濇ZS3 `�q8�  ���Hd_��b��sl� ���;���mv���   �ʹ����*s�>`� 2UI�C߿N��J��j���c�������r����� .P��E��WhV�v�1����҂�5:n[�|Qf>�cW:�Bkxf�v�1G��Ŷ���`ߐ�o����j��  ���"���#  @�sd~e��W`��3�[�	   =�,�'�� �U�6���Y%��k��ͯP�㱝��
[{�����Q��c;�M�m���Vu�k�isU7��0kCA[�N�Z�9;�O���Bu-��kQgq��.��'NӨ��|�� �Tb���v  H~���X4�%��vp�Xp����=�#  @z�
��N�W4J��� �&�t�'�t��=ڽx��O��h�g;��L�����������!
[{t֓UZ�a�v�6[�'N�H63��QE]��WPE}�� ���G�Z�U�<���u���5���z�| @��{}��lG  ��`�뇣�H��vp�Xp�t����  �>�4:"�wF拶[  3�g@g�ڮ�kw�qN��-��ȴb�~�*�?�9�uܶ:M��� C����U;t��]��1��?���u��u����`GnߐN_�S�����C�| @*3�rs�`��  �F��ȓ`�i���6�x�  ҋc�o��/�ǩ �r�F��/����<Q�O������Ͷ����F�ZӬy��UQ�*�8�� @�kg~o��?e�j�O������I�2�_>���-2	f>����3����^P��	\�-f>  ]$8�  !s�K���N���3��#����v  H/����hy�s��m� ���;�t��:m�.�V���
�_���a0	G�M���/�Y��=�� o)��_��٥�kw�:�돛ʲ�ax���R����$ xKy]�Z�v�N]������+4�u��b� �P��0�	5�lw  �4c��q}�vp,Xp�`�q��   ҕ�ɰ� i�8�JB*	u���;�4�H��U(4��%��㍏���]��G4}D�a�������g�ޡȴ���Rr�﫼�Q�6th����U7�"���3��r�ꏛ���%��c;/e�:�Ú�?�� ���̮]��  8b�x��X���Ď0�?�ʑ�|��j�   =����e��X[2 �F<��*�ZTQ�"I�T�25�.Us�%<˅�kb����[U~�Uu-�E㶓  iL�QE}�*�[%1�_;�[��l'@Ҙ���m*?�&�3�e��f1� HK����N   �ɴ������42�n���8��H��;  @z2���������m�  ����Aͯ����E�^�L+RKE�Z�NV{i��a�;�T�PI�S��m��=h;	 ��kf~����S�:u�Z*
�|��f~g��Ý7�l'��������\9Y���2�P����y]�*w���� p�_sc��  ���1���H[,�g,���  @zKs�qĂ; ��?W�&Uh�$�fy�^Zphٽd�����W��6'������G�[{U�PQ�Sك#��  %�Gb��iRe��f~Gi�Z+
�^:I]S��[8!mf~p`X�=*l�Qq�SE�N�0�@���TYӬʚfIR��Q{�$�VLV{Y��������[��.�;��  Wrd�3�c�  �/���c���I
�n��逿�7} ����|�Ec=��m�  �/k4��p�J���٨ף��y�*�WW�D�LP~���s��ƽѓH(�wH{4�{P�*h�UA[������ �*k4��p���~�gy�=%O]Ey��&�??�����3�Qn�&�jB��&u����W���| 8�DBőNG:_��Wg�+s�� ��u��\E���(����:�gP��{���^^Z dG	-  �Ĵ��E�+��A�-��`�=9��n   ����G�+�$�z�- ��OhrK�&�t����??�����r�5���H�_#9��'�W�E~IҨϣѬ�W���q�����UV<.4��PT�CQe�(0U`(�ʂ㐂�C2	����5��3$ۯ�I����`0[��@�g�(������Af> ������A����9Es��>4��n�K�����qe�G反*04���7��=�
�1� �ΩʎD�ٮ   �ϑs��a�i��4����v  p�x�wL�w �+�QMi~�R �]�Q����l� 0��Q��o��  Ɔ1��� @R������.I�[�#��q�5;��  �������v�         .����#  �;�F$��vp4Xp�0���  �=���c�;         \�ŜH��v  p;�HS,�g�D"��  �.�        +#�g.   ��rr��L���H���Q��@S��  �]�JJ���e�         ��feqh!  H*s����'lw G����/  f���<i�         �m�nl��  ��q��(����  ���:        �(��  Ɗ�$�K��	�3�Q�?~�v  p'���        ��h�m7   w2�Ƞ1z�vp$Xp���   �eB�!#��v        @�1�47첝  �ˑ�b�8,�g#=n�  ����	�         i��3  0�|��OHJ�� ���z'MZo�  ��ϟ��$�v        @:1�á�  `L���6I/�� ���y�����  ��<�$�-�;         ҇����]  ��=a�8\,�g ǈ7} ��p�u        ����B  0^��@:a����x�)�   3���        �ar8I  �8�M�A���`���^2--��#  @f�55n��b�         8�X�C ��1z�vp8Xpw9��3�  @�0�#9���         H�Mk+ �q�H+m7 ��w���Â;  _�p�        �6�L  �/V�JI��;��Â��xs�lG  ���xVHrlw         �2�,� �qe�d��v�vXpw1GZc��  2KnccD2{lw         ��a���v  �<NB+l7 o�w3��  ���        �7��D"��#  @��[�4����9�g��  ��<��/     ���ޝG]v�u����95�2��*U�y��"��!L����� A$�p	��(.Q�Ah�����A�!	AW_n�Ƶ����W��4��#d"&��U�<�9�w�(��J�s�{��z�O��Z�:ٻ�g� �}(aX ��r�E�]�p0��u�����rv 0��KK��     �6���� ��T�����?gw����T��|��� �|*��vW��Bv     @ݵ��|� ����p0�=U��Iv 0�j�     ���?���^��  �X��t�j�=U��g7  �F��/     �=j1( R��=�/"b_v��~�}�7|); �o��?��&�     �UJ5p R�k�Y��%�{�(Z�� �d�n�����     �"�G����� �Z���e��G�� Z��     �?����k_۟� 0�5���{�F��  5�ϲ      ڢl: �v--�EDL�;������u뾘 Q��?�n      h�Z��n  ��(��枈�Rv�����E?e ���[��6"n��      h����; �%\H+��M�>l �V)��      �ߗ[ou0 �~]��2p�6 @�Tw     �2 �]j�8T�V2p�:,� �v�9+      � m��替wdw�=���?l���k�#  �n���_#���      �TJ��� ��+5"�[vܓ�{��(W�� �5�7��'"���     �h:��bv �=�(_�n�{2p�Ƈ �V�S     �9V�g�馽�  �����1p�2 @+�(N$     �� �N���2p�Z�L �V��     �_Ŧ h�7��Ո�+�����?��p��dG  ܛQ��n      Hd� �R�h"⯲;�����/��! �:妛�Y"n��      �0*��  �ͯ��.��A h�&��
     0��+7�p{v �}���	pw�}Qꗲ  ��_     �N��?�  ��Ʀ�V1p�2-_�n  8�R��     `�� ��F7��*�=1���! �ݚ��!     `�hl: �V+�^{g��)����{?�Zn���� ��YW�_��&�     `�w ��j��i�>��A h�r�M{#��     ���֯��� ��UlQi�>(�[3 @'T/�     ���r�wfG  ܯ��t���x� ��a     �5�M �	�46���{�:�jv ��(�^��      0+%�o�  �he�M�a���Q�P :�ܷ      s�ֿ�N  8嶯�{�; ���&�l�.; �PL���     ���  �rmv D���ߗ��^Ɏ  8���#b)�     `��� �Q���h���>L �)MD�}v     �4�7m� ����h	��+>L ����=     `.\W���/� �Q��� ����j�6; �p��     �y`� tJ8t�v0p����  ��D\��      06 @�L�Z����J��  Gc�     ́j� t̆n������n��a �R�c.     �%�w" @��k�Y��[�;���ۖ��[oˎ  8�C'�     �W�C �*a�A:�.+qC�h�3  �׿~KD,gg      ����� ��Whh�n�! t΁�ʍ�      ki����  �����g��e�z :��     �c����ۿ�] p�J�m*��;�ܜ]  pd��      }V} tR��t�����J�[�  ���     �ϊ�B �N����0p�Z< �TJ�0     �V�� ���ǐ����J�C ���     ���B ���/�l:Hg��a�L}�  �TK�u    ��*��t  �t��n��&;��f��a+áa �I��w     ��ju�; �M%b����|3p﮺i˖۲#  ��t�E=     ��j8� ��^�T�U����^ɮ  8�ܞ�      �V5| t�]��;�~+�  ��}�kߎ�&;     `-4��#� �H���eHe��]>< ��*�����      XM�8� �Zý�ܻ���  ��xa     襍���u  �5p3��;���A ��~     �i�~��� �#UmTIf��Q�  �>o�     }tg���  G�TUr�wV�3�  �h��     �*6 @�l:�e��Q�?e tZm��     ��Wm: �N�a�A.��b_v �Qڛ      �| tڰ�3�2p��a �>�3     @� �4U��wU�� �6C     @Ո}�  Gæ�l�]5�0 t��?�     =40 :�{d3p�(o�  ]�~     �#߁  ]WKq?C*����  :��     �K� :m�`�~�T�Uk]�n  8*��?;     `ՕX�N  8*զ�\�]5-�� ��Q�2�n      Xu5l: �n��.�R�wՠ�� t[q?     �O��  �q��He��U�� �q�/�      =T�M �m�6��!��{GUw ���3     @5�; �ۮ����ܻj:�� tZ-��     �Z t��R�w�`�� ��`0�n      Xm�Rm: �N+5"��旁{w��  ��Q��     �^� �^�#��{w��  ��Q��E    �^� ��� ��j @�M�f��      �ښZl: �N�a�1&��|]5z :�ԁ�     �j� �u�gHe��Q�� �u�3     @� ��۵���ܻ�� �ZG�	      ��� ����� ��{W5C @�U�3     @��ph! �q++�gHe��UC'� �V�q     �6 @�w�M��;�Dl�n  8*Mq?     �O�  ���Z��n`��w�4bSv �ѩ�g     �>� �i�j�A.��*� ��s?     ���@ ��s?C6���� @�5�g     �j� ��+6$3p�(o�  ]�~     �R� �n+��t�����|x  ]�~     �#߁  ���B��wT�� ��sz	     �Oa @�M�ϐl���)����  p4J�j����r��QO=5;��3h�y�a��� ̷�:�- ��0� �� ��J�ǇM�ܻ��d'  ���se����ח �r�9��/���@�r���  �| tZ)�Z�+�g->������ �y'e      ��j8� 讦�Q%��{Go� ��~     �;v�� p�J)6�2p�b t��    �^ڿ�d� tW��eHe��Q�� �U܇��     ��á] �Y�:��\�U�� �;N��     @O�R�: ��*6�$3*���]�#  ��Ғ7}    ��j�rrv �Qp/C*�۷w�� �#1N�f7      ��R�Ӳ  ��{R�wب}�  ��DxQ     �� ���箋���;�o�6x� �R��     ��J�� :i�-�l�����|3p��� �Qe�w     ��J�� :i�46�3p��� ����x     z��_� ��T�T��wX��/ �Q%��      �� ���:��t�]Vckv ����     @��t  �T�M�ܻm{v  ��);�      �бuǎ��#  W��M�ܻ�� �z�t��     ����Ʈ ����t��6��� �ñw����>�     `-k5p :�:|�0p�Ѿ�ŭ�  �c]�x�     ��8 �&���w��۾ @�x�     �� ���Ǜ"��0p�8C @���     ́b� t̒�Z��������  p8��     �	��  �2t�BK�w\��3� �p��n      Xk�w" @��Rve7@��{�0 :��     �@�X���� �C�=Z����- tG=p����     �(����� �CU���
�Ww�ݻ�gW  ��۶m���      31�:� �Z�{Z�����Kw��T �F��!     `n"|7 tB�(Qï��
�=0*�� �	��     ����<(� �P�[XX��M�a��M�n  8��G\     `�� ��9l�1p�A���  ph�ò      f�F�n ��4�[h�>�� �n(��      f�Dl���'gw  ܿ�-*�a���b @���xSD���      ��IӜ��  p���;�a��'��gl͎  8��:|X��     �L�NC :�a˴��QOL֯�` �mи_     ���i� @�Յ�S"bKv�����x Z����7    ��S��
 �ۤ�_�U���ԇg'  \�0     ̝a� �Z46���{<*;  �`��n      ����n>ckv �}��n    IDAT���V1p�g�s�]�� po�֭�k�8�      �d4ydv �A��*���q��[� po&��!     `�9 h�1�(�3p�2h< -e�     ̱�TT ���ϊ���pw�� Vգ"�c�  �T�JQ����~��� �����Ell��~��|+ zop�F����I�����gg p�?+���3�5��v*զ��i��r�|�  m�>��7��߉���gg p?O{jk����c��7gg ���y?�ځ{|���[ �q屏�b���Au��˵�ޙ �]�xd���n�� VQ�GU�� -SO=���ؕ�     ��L�.?2; �^8���1����m{Hv ��M6lx\��     �ݠy|v ��Ոa�xLvܓ�QϔR���  p�O      J1p Zee<>'"���{2p��a h��O     ����8/� �8T��2p�b@ �K�x\v     @��m�x�=� ��9���2p���~. h��۷?("N��      h�a)Fd @�8��V2p��d���� ���2��      �I5p ڡ�q�"����7�}4��  ""J�/     �?)Q�/�  "b:�|_D���7�=Ԕ��� �ܗ      ��c�x�); `�46���{�O��� `��;N���gw      �ȺI)~ HW���Z��t�ʶ�̎  ���d���&     �wi�1 ��;�(snv����*? �x�     �{�Z�?� �o�R΋���p_���۾ @��G      ���gl��  �_����{�F�W��� @��y�qQ�Q�      -�q����� `~�Z�i5��:ye<~dv 0��6<)"F�      -���  `>���c���;�`�{�D�`v 0��Z���      �V5��R ��iyRDl�1p�1C @�Z���      �bO�'�|Bv 0jilKi=�~{b]\<&; �/{"�Y�      -6Zڸ���# ��d�N�����I�<1; �/�Z�%�     ���e ���-[N����;����\C �l�     pP�w* �L-�;��N0p��i� ���%�<%�     ��o<ޑ ̏-����� �|XY\|lD���     ��R���  ̇1�O��Ca��e�ĳ�# ��P�w      �Z��� `>L-�#��@-� ��(Q�w      ���:o��  ��qh!b�>J�S< k��oGģ�;      :䘥��dG  �W�L�����c��<9">� �׺I=?J���^:�\tQ����kj��|&�-�d�    0'���Gv �_{���qNv*�9�4q~� k������G'��O~2�#�]2?~��1������%    ́Z��5��%�W- ���r~T���� f��8��' `m���c���X}'��O}ʸ}�N9%FW^�q��.   `��m+۶=:� �z��d��9Q#V�� ���4~("��� �N��'>�~)0�������x��    ��:</� 觺s牥8��n1p�#��� �~*�q���N8!F����۳sL�~��^2    `͕��n  �iy��#bCv�9R�>�F�� �_�]"ʳ�; z㤓b��+������c���Eپ=�   �~;si��� @�J8���1p�/g��Ǐʎ  �e�o�S#����^8��]qy�ݾ�j�SN��G?q�q�%    ��`0q�; ���x��F}Zv.�9SK�& ����M_�Uq�)��{Xv	��<��1�ЯD?�   �ڨa� ���RΏ�M�p���L��m_ `��s�]�:���N=�������K8��ӟ�K.��    ����??$; ���B:��}�����xNv ��o���89���N=5F�_��.��-Q�{Bv    =5,��� �����vlD<3�����<j�e'  ���� :���e��(F��Q�n�.   ��j��� �~X�{nD��G��}�(/��� �R=㌍Q�s�; :k��]q�q{m����pĺu�%    ��Y��̎  z�8���2r�O�'۶�/� @�-//?'�����I[����WFyș�%�r�1���dg    �C�c4 ���œK�S�;�H�ϩZ� ��2� Gd��]��(�ve�p��xE����    z�D}a�� ��J�?�;�H��_�ݻ}x G���qR������ٲ9FW\�L'��B)1���<�A�%    ���ɶ�O̎  :�V��i����;�xzv �M+�悈ؐ��%e۶��Dy���SXM��_�qcv	    =R�E� @7��wD/��i�slX�K� ���/�. �2���WF9���@9�^ziv    }R��:o��  �gt`jL��<�j�g׭[7gw  ݲa�̈8/��+�������G~$;   ��8q�~8; �Qj��y��m�J�(; �R��"�dw tAYX80n?���f`���Dy�ò3    �R��. px&����e�>�J�߲ ���A���; ��,,��J����qc?|Y���g�    �O�ڎ�� @wԩ��w�^�� t�ta�5b1���ʎ1��UQNߑ���;c���dg    �e8��8; 膺y�qQ�y��܉��7v �CR�xiv@ە��^��(���W��>7_��   @�����  �`eݺ#��Xn���zq�7eW  �V�n�\K<;������1���Qv8�}�/�4����   @��N��dW  P�+�`��񀕈�# �v���+"bCv@[�>0��(۷g��6��×E|v	    ���� @�-/,<"J<.�V��;���� ��jĠ�rIv@[�>����۶e��"�3b��_��    ��j�g�]\\��  Z�'�`5��h��[޶��������) @�L�M}`v@��;cx�Q�n�N���~v��������g� ����@���Y�?���G"��Y�?  �cF���� �}ꩧ�R��������*"^�� �Om�_{�e׮]yEĖ-����Gs�g����E�f��o��s8�yO�θO�K/��߿��_�NX5��?=/~��������  ��&ʫ�羻\}�Jv �.+�׿8"����d��ݔ��?[���� �=����k�3�; ڦ<��1�⊈-�g{���h~�7b����o�l��R�U���G?�O�N�w6��×�䇞q�]�5    tP�ض��o<+"�0� h�rIv��Av ��ieҬݱK @'kyUD�; ڤ�y�wNn��^sML����������n߾���Q��O�K�Sٹ3��~wv    V��&� h��������Xm��C}]�� ���k׆R� wS�q��َۛ�~6&�|Vԯ|e�����c�җE�?�]r�</Ͽ ;   �������s�# �)��	����]K���� @;������-� mQ��}��SO��u���w1������u;gi)&/}i4�G�%�i��wGٹ3;   ��*M��� ��m�vz���X�|�A��g7  -Q�$��r�Y1���[fxr��JL��Ƙ���M3��v��JL_��h>���{w�1��_�X�.�   �N*?VO;��D @c���fw�Z0p��<yya�� @����i�g."�<�a1���SN��E���_�W��}���W���'��sΉ�O�tv    ݴa2]� 䪧�z|�xyv�w�]-?��  �jJ����6(�w���OE�|��.z�1y���ٟ��}���K^����K�����Dlq�    G��O�ݻ�gg  yV�m|yD���k����P_�'� `~-��-5����-e�~�m1���Q����]��&��������f�|���c���fW    �A5b�|��?�� ��(�u���ܹ/�#����*1���(� ��9����+"N:if׬7���]�+_��5{o:���*��~6��{^�N��    ��J�o��������pAD<(�֒�;���xmݹ�OX ��ٻ��Q/�� �TqN�>�Ɉg�HTo�1�ϻ ����sc2��k^Ϳ���%���c��WeW    �M�L�->=; ��R˛�`��s0'N��^� �֨�o���� Y��g�����=n�-�/�(������f2��k_ͧ��.�.�K.�ؼ9;   ��Q6� ���������Xk�\�7�ݻ� `N|��[��̭r�wNn�fw��o�ɅF���]s^M�1}�������iS_��
    ����,,��� �N��7悁;U#V���� `6&KK���Y��я����v�~�1y���Ͽ��5��t�7�t�F�X��8;   �.��g� ��X^XxdD<9�f���CP~��� �W��5^����<�11���#�?~vݻ7&]�K_��59`:�����g��~}^���
    :�Fy��x��� `�o�����`�̡x����� ��Z��+#���Y+�yL�~�c��7ML_��Q����]���4Nr����.����.�r���    �gPJyKv ����m;�F�q27�9$�ַ9� ���q��R��%0�c����l��1}�ۢ���q���^�ӟ��h>��쒈��)�    �/�??$; X;�1l8�#��s���充�eW  kceyrI�X�� �����w�L����oF��>2�kr���~1�����\pA��۳3    �� ��eG  kc���#�fw�,�s�J�ow�; �OݵkC�����Y*�=!F�Xı�������b��w����Zc�����#�/�F1x�s    誋�/,�� ��AӼ="��0K����{y��s�+ �յ�w�%5b1�`Vʣ�����M�fz���/���~*�ifz]Q�1�ŷF�ۿ��1x�"F��    :i8��w �����3w�9,�Էֈ�� �������� ������|���VL_񊈽{g{]O�1}�ۢ����kز%���w}    ����۷?(; X=�Z�NGb��s������� `u����*���������egp��oG4�]�v��eKڵ   �Ѡiޖ �����C���; ��;���xW�F t^=�c#�[�; ����'����38L�w�+�_��9s�   @�ոhya�� ��F�'l5�S��3W��dG  Gg2�!"N�� ��n��;.ͮ�M���h>���    p8��wdG  Ggy����(���,���uq�� ���;N�5ޘ��w���7bϞ����}��9;    Y�������; ��P��FD�΀,����R뫳; �#�<i~."N�� �z��\uUv�`�����|pvܿ4�k   �K���f7  Gfe��'E�S�; ��;G��[��'��� �z���J��dw �]�ꪈ�$;�U�|��1�����u���M4����_   ��+OZ���] �z��v�k��S�7�3� ��YYY�4"6ew �]��W�Xeͯ�JL����������/�سg�   �ܨQ�Wm� �S���ew@67��R�M���� ��YZ\<'��,�`ԯ�mvk��Я����^�?��;c򢋢~�����   �W�ZYXxqv ph����K��dw@�s������ �5���fg ��t�ￖ]�i~������Z�?pϞ�������3    "J����vڱ� ���|�[���]����/o���� ��&���,Q���0�7F,/gg����.����Q���A��1���~�    wS#&���; ���;v�Tk�%������0�A�� �ՈaS���; �ƭ�d0�o�VL���#��o��Ϗ�W��a    p7�ƛ��o��  ���d���89������Q������:; �w+�^5��0/ꭷe'0#�o�NL�g#n����Gw�ͧ>��?#�W��vq    p�q+++�fG  �n���#ʏgw@����A�Sw��\�暥� �_ԓO>a�Է�(�) ��p��t^��OD��ODl�e불㎋ش)�ƍQ��1�F|��K����={��   �;���[���������% �w+M�`D���61pg5������xov �/V6n|W��5�`��a�>�n��N﯉)    p�4�\#�X�� ���x��q~v�� ;�~�Qq�x�#� 8`i����� ����    �{���m�eG  �ݻ��(���md��j�4����%J��Z�+�����;    �>��ԝ;O��  "&��#���h#w�@}����dW ��[�_%~ �`.�    �t����_Ȏ �y�waa�����h+w�Dm�j�(� �Uݼ��A��gw ̫����	     ��D}�Ҷmgew �<��@D��me��Z9{����� �W+�ֿ�F,fw ̭}��     �˺R�e5�d� �<Z��fw@���fj�K��v��; `�,-.�?��0��   �V+OZYXxIv ̛�k׆�C��vM���׳# `�ԈAi�#b]v�\ۿ?�     ��j|�nݺ9; ���}o���dw@����J�Zڶ��� �+��OD�y� so2�.     �?����ˎ �y�<~H����w�^��Vw�<1; ��n>ckDygv ���w�Qr�u��?�[��YYH�]ϭ�4!(A$�(*�Q#��
q�N��0�Gp �2�+�����QA	*"!�&.$]�V���e��]O-��9z8F�9�J�s����       �9���t��  t:�,�}NR_��0pǘ3����0� `�����$M�� �4n\�       �����0��	 ��+��%��h��$�Ƽ2�w�
  :�H����;  �0p      �>��eْ�  t���O����h�ĭ8ӫ��C  �4��;��,v �L��        6��N��� �N����J��h'��LO�
} v  �&�N3�@� �Cl���       `K�����9}�C  �$Y%=��/����h*��=a��  t�z��b�^� �O�L�]        [�I����Ď  �S����>�hG��l������q�C  hw>m��E៏� xSy�       ��c��d�ʼ�  t�z��9I3bw 툁;b�%˲�bG  ���q>!i0v �_�dnp      Жʲ�L�;�7v  �¡�zy��]1pG&{g>P�'v  ��K$?.v �Qp�;      ����lݺ%�#  hW�}6v���#��}ѧO�; �v�3L�,v ��Y���	       ������2�w�  ڍKV.��$M���3��w�{{�;v  ��� �?v �1�i�       �����Ņ  l�<T�d�cw 펁;"��k���cW  �.�J���� xlB�       �F�c��wj�
  �E-�]$_������f��  �Ս�$s�~ �`��I\l      �͹��t~�  Z�ϛ�cҗ%M��t�h�Y�t�K; �V�R9i_��]� �汔[�      ���u�ϚU�� @+�V���dO��t
�h	�:0�T��  �Ue!�,�ٱ;  ��v�)v       ��yV���R�  ZQ^�>�d��t�h�d!�; �V��Љ�;  [h�α       `t��_U�_ �?�E����Q����O�����'� �U�A �Wr�aRoo�       YM��    IDAT.?9OS�8 �&.Y=)}��J���0pG�����}2v  ��B ��lpPɫ_;       FK�]�����!  ��z��ݥ�cw ���;Z�1Y%=2v  ��Cx� �����Vi/�      �1��z��#  �-|��>��T�њL˲4�#v  ��i�l��A ��;���Ǯ       ����,TŎ   ����GRo��S1pG�/�E>m���C  h6��)�Œzb�  �]�7�v�=v       �"?5a��  4�KI�h�/���[�N���l�|��3cG  �L.%y�|�Ki� �()�U���R�-      �=�]�3b�  �L�4}����t:�hu��
 �U�>$�� ����7Iy��3m�]Uzm       t��yR��K��-  4C����kI��0pG��ei���  ��z��7��� ���'׫���K�zS�M��f�Svo�       0�����bG  0�֧i�]����`��v���___���C  +#i����eI� �A��q�;%��Z.����H�&5�L       c.[R�T_� ������ʅ�*if��[0pG[0�@���}Μ��-  �6�>}R��5ISb� @7).�X�����gڎ;�t�i��<      ��af�������!  ��<�Z�g�� �	w��g��7,� �hr��=}gK�o�@��_T�O4���/Tr�	M=       ��$K_��a.t t�,T�,�kbw ݆�;���Y��.v  �%�%nzE� �f�S?�bYs��-��=�g=��g      �{B�e�T� �h�C�K�Scw ݈�;ڏ��@u��  l��1���  H���⢋�w`����>'͜ټ3      `���Y%=)v  �jCC.�����-@7b��v��_�a``8v  [�V����_�@kpW��w�����9s��_:W�8�yg      �3�{k!� ���3flW�}C�U�0�B��YJʗ����!  l)�1<`�_*iR� �?h4�x�"����iG�n�����K�r��      �1f&;'O�g� `K���{�Γ���-@7c��6�fYv�K,A  mÇ���=��%͊� xy����oڑ�߾*-�H��      �&�o��͎ ���C�Q��$v�������y�� ��p��,���g�n <�T?���~մ#��W�4�<       h��I���gϞ; �͑�p��w�� ���e!�1v  �'����� ���׿���#��}ӎ,��D%�ڴ�       `�����ȅ.�c�  �X���ޒ}.v����C�i�4=(v  �&Kӣ���� �-p��jz�|Ŋ�g���>��/m�y       �&{Q���� ����u+�!�7v����S��Ey�>;v  �,O���:C��n l_�Z���9�J*�~����9�      @S���P]� ����`��q����[ <��;:�w}k$M�; �ժ����5�/ �-���?\Z��9��*��L�߾�9       ��������  <ȧM۾�Q\.iV� ���fz"}�g�� ����a��&�n l��oT?�hi����ӣ�gȞ���       c��:3�WX ��y�z�q�/��G� ���;:�kv^._���c�  ���������n ���Տ9V�՚s���*�w����4�<       {=.�$KSƄ �h\�|՚�$��#c��eO�J���y�zb�  ����O�]ߒ�K� ���k�U��o����8~��眣��6�<       {��u����c�  �S���tT� ���;:�I�׬�ХR� @��y�z�r�bIω� �������.Es��Q��W�`As�      �1�R(��W��Y��- ��W������; <6��h�zY�O��  t�J��5_6��@�+��55޿�y�J*}�T%�Ӽ3      `l���Wx�:-v �;di�:7}(v��������Jzr� @gs��>'���- ��(��E5>���X*����U:��R�ܼs      `�����m�1c��) ��V�T_&קcw �<|G]�L��C�sϪUM\�  �I�KM~B� @s��.�~��׽�ig&�+{�S�xӛ�w�ٴs��٬!�3�;�c���c���Ųu��􌮱~���/�]    ��yO�7|Μ���j�c  �'� �_ ����a����S�J�Ͻ��>#v ���i�>w��� �8'H����WѴ3m�=U��﫸���~.5M;��5�*��=�=v	�QfO{�J�}"v6S�%�:��Y��   @;�����t�I��1 �ΑW���¿!�/v������d���R#w �h���m��`� @D�j��]�v���%�;��Oɱ�J�ۼ3��;NTqᅱ+      ��⮗���B_��0F� �ѐ�鳽�oI����Ib Mf2�\�R}u� @��Bu�\�� ��B�Eo�_}u�����O�>=v      �u���<��T�� hoY{��rI�b� �r�э3?���C  �+�5��� �B�u��V~�u�K���LQiɒ�      @�zeҳ�] `+ei��dWJ�����At��ɾ\���! �����1��!�b�  Z�Ȉ��'����.�6J^������      t�c�P=��~ `ժ���JҴ�- �wt��ɾT�T�=v �}d!'���Q �G�׿���W�o�5v	�Q��Ə��      t)?.���e� �\Y�>�
�Z��[ l�Y�v�f~q�R}u� @��*�$;S| x<���.���%�64����;      �^���z���9 ���B�S��%͈�`��� ����,M�� h]Y��N����O ����ܣ����'v
�A�p���O��      t1?.��.�c�  ZSV|�dW��ہ��@ب$��Y�� ��<����x�! `��w�q���ڵ�S���e�N9E*�b�       ��<����y=�C  �%�2�ZҴ�- FO6I$;3��=��W.� hy���]�� h_��[U?�0�/�X�~��9�
��S�y��sΉ�  �m`�>_6n\�`��-���yg�  ��+�k֔|��#l��,v  �<M�uץ�O��`t1p.��sy�{V��h� @<.Y�K��?b�  ڟ/_��q�Q��/Kj�R�]��W\!_�*v
   �R��Se�3�1�X�D~�bg  0����|����/����[� @<�4�_�.�4>v�ї� Z���ZK]��1 ��s�����ĸ 0z���T?�5R��N�֘4I�3�I=�      �l���{����C  q�B����51n:w�Q�lq^I?��:���s���!�@�b�  :���j��R�;[���T�����       L������`�� h�,�7��˒���`w��bz]��}�<�a ]�C���]�MI��� �\���V��wJ�S���W2~�       ��=�����N�K  ͑��b�>#��@��9���֬����O� ;^�N�eW��E�[  ����"5N:)v�R�?.�y��       �;��5�����K  cǥ$�t�/���9���\��5>sf� ���000�~����n t��/���bg`kL����?/M��      �z.U-i�8��� 0�|Μ�<��K�(v��a�l6{Z^�n$�'�. ��Z��[9)�X�.�[  ݧq�)*�<3v����D�>�I�,v
       i�'~E-��c�  F�M�ׯ�B�a�[ 4w`�������!<7v	 `��!�o�~�R� н��^;[!9�EJ^���       6�5���P=)v `ۭ�VӼ޸F��c� h>�����pH� ������}[��c�  �����X���.�V(��ݲ���c      �E�ɗdi�	g m+K�=z
����c� ��/䀭3!�}-�űC  [�%���Ir�-�'v  ��FC�7�I~�b�`K�J*�3����%       �zkVI/���'�N l��2�B��q)�nw`�\�4�L�7��$ ��3�/��&_"�b�  �0y��������%�RS��t֙���K       lb��}?��S @��*Յn�e�&�nW9v ����|��a^`wܱ.v ��y����.�sc�  �6lP���U��bٓ��[���U�S�X�(v
�G�׿��#vEǰv�&��%x�b��h����U�7v    Ĵ{"�IV<�w���ǎ <2�Jy��&��b� h܁ѱ��?I���V��5v ��j��O�U\*i8v  ��U�U�V�k_��S�l���/��x��sΉ��W\��+bgt��ҏ(9��1��/�|��1��    �ä����V�ٷ���� <�O�>)��������u$���s�6�V�; ��R��ĸ �N�_�#^%_�:v	�P�N�=��3       <�D3�$���v�b�  6I�'�}כĸ��0pF�t/��<T��n�塺8�}]Ҥ�=  l)��n5�R���)���g�!͜�      ��%n�p=���iӶ� ݮ>P=0q]/�I�[ ����+�|i�y^��� ��g�خ����|��z ���P��#�?�9v
���*��R��      �?q��|����͎� �����/�4%v��T� t.{U^��*��z���k �[�T�s���\sc�  0�׿V��cU:�$^��(l�,i���c�y�Jo�;5v
      ��[Rj�,��U��� ��g�خ^����_�@kc����&f?�+�W��^���1 ���i:�(�˒�/ ���O���_;�e���J_:W6���oK-R�ɯ�A�       �j�˾�����U��䱃 ���T�;��_��ɱ[ �>��3ـ�}���]u�L*b7@�q������))��  ��׬Q���U��b�.O���$Q���T��ҽ�Ʈ  �z�#��z{bg c��^; �vTr�G�!}��KG�]w�� �h$�C��ϕą� 6w�9�&_R�| ���3�t����  "�ӟT?�0���u��p욇찃ʧ}B�W)<�  ��rK�   �(���_d�z׬�Y� �.��N6�H��= �7�M���� :A^�<���n�ĸ  H�ݧ�GH����al�}�����3       <�YJ�f��[b� @'X_��yH�1�b1n����7KI�,����v��!��-��K!v  h~�]�{��aC씇)�k��)���       ������,�g{b� @�����ʅ�(i��- �w �񒝕��%>445v �����R�}TR9v  h=��_����I�z씇��*}���ĉ�K       <�cs�Y��; ډK�Z����I��@�b�D䮗���/�xR 6C���Փ�M&�  �6��j5����c��*��]�3       l�]�.�T��Ŏ�V�!��<�ט|��R� 퍁;�,�]SՓ�_� ����	�+]
�{  @{(�;_ŧ?;�a�c���_�       �g��O����=Mw� ��V���$�I��i��P6��<���Y�*�c ����W�k7=���.  `�4�.U��o��x��J�~L�:5v	      �����_���c� @+����Yg��W%�� ����Z����-�J�U�C �dizT�(n���[  @�rW���xc쒿��~�>���       �̠[qM��>gN_� �-�V����7Jv|� ���;�z���yyH/�juZ� ����g���Ε�]�  ��j5�_���U�K�.9�%/xA�       [�$[��_C�Sc� @.��P]��,�	�{ t&�@�riA^�/�4�/v 4S}�z`V*����n  ����8�8i���%���Ai���       ��͕��Z���R)v 4K-�]��s�RI=�{ t.�@krוY�~�C�; ƒϞ=9��E��6��  t��f5��v�=v�$��T���5v      ���c�%y���; ƒKI��Lv�dO����1pZ_"�[s�_q�;�NU����~%���-  ���]���bg�]r�����       ��흔7硺���t������^%���������5�]Wei�̧O�; F�O��tY���%��  ݡ���Vq��cgl�ӣ��cW       �6�]�4�j!�; F�KIV�.L�/%��@wa���ka���y�ǎ�m1���,�Y���[  @�qWc�"�M��]"IJ9X��      t�g�����������:�/�41v����hO�.�"ճ�Z�; ����!O�Kٷ\Jc�  �.52������.�J%%��?      �C�s��<M���t��1 �%|Μ�<�%�4n���{ t/�@�2�_����R]�����૫z�kw�<v  ��\���'Hy;Eɂ��ɱ3       �����Y��>}���9 �x�J�y���]v����= �w��M���<M���.�c ��di��<��n|u�o�  �A����q�ɱ3���,xE�
       ��,٢zo�oj�*��hI>445K�en�$�5v H܁����d����?}����9  I>c�vY%��\?����=   ��8�*.�j�%G-/�      :�K��/������4v H�K����y�q�\%�M
 -��;�Yƹ���u��izP� �m$���ޛez��r�  ���x׻俽5j�͞-{�s�6       ;�zY��[k�z�ϙ��@���t�<�?��I�c� �?c�t�9��ZH/��;@w���K-T��Ⱦ%iV�  �Ͳa����aCԌ���z>      �17��K��~U�V_;@w񡡩Y���sIܺ�e1p:�I�R��Y��������|xxJ��&���_�  `K�ooU���ڐ�"��'j      ��ع(�r./�.%Y�����l��R�& x,܁��+٢����Z��d�� t�JY%}m��n�T��  ����"��O�L�(M��|       M���k��\^`,��}��L�s%͈� ���;�=f��+y�^�W���3�!쟇�F�>/> ����H��η���       ��fz_�����R}�s��Q0R��"O�I{���-���6���?���ґjuN� �V�<��K]v���c�   �&��&�^/`;.i      ��t�����W�4];@{�juZ-��I�r��/Ж�]ʤ�I�˳J�qO�b� h�,�3͒_�4?v  �X)>�)��>��;      ��v1�E��[�V�p�f���qy'���d�%��n�����n�2�=w�Qa�O��}�  ����{{��$;^R)v  �X�+T�}v��m�       H&{�~SҋF�՝c� hM.%�4]�g�[\�1ISb7��b�@��3��|���硺؇������b������	��   ��q�'��k�����&      �Ve.-H
_���C�  ��%���<����"�w�� ���;�4��K�,�M���874]�����BuQ^*�����^  Ѝ��#�f�~r��      ��z�Z��(~Wa�W��b�'�T_������zb� m�<�Yr}1��e��B�ʱ� 4�ϝۛU���7�&��f�n  ���җ�{�m�k�y       ���-��3�t�9�?v���CxnVI��Ϳ#i��= 0V�x��̗�!e�t���׮��̗�T��  �j55�8��GڤIM=      @[�N�Ey��,��}��@�  c'a�,�׹�G2=?v �5� 6��W���    IDAT���o���y�zb^���BuQ}�?0l  xdŹ�J�S��8�yg      hw��=��j!|�C�;��W�/�B��])�Y�{ �Y��;Ivv�z��J�-����hS>}���R}K���$?ݥ�	  �e�_���_l�ye�)      �Ŷ3ٻr��Y�~i�Z�9v���R2��Y%��(�rIό� ����֘%���R��Z���i�C�  ��g�쯅�Iyo�]2?�a;  ���K.�ܛsX/w       [�O�#��S�Y�2/v���s��eizT�[ٷdzF�& ���;�m1��KrםY����R�;�#���K�g�垻L�DҔ�M   ��W���Z՜�z�      �f�I�e��j!�,�T�;�#󡡩y%}O�~�]r�+鉱�  6� F�D��R���ZH/�C�?v�������"��,�k$��n  hW���sP�ܜs       t3� ��YHo�*Յ><<.v idpp�,���zc��>$if�& h���Ĥ�.�2�Y����q� �d��*����G.-�T��  ���曛sP/�$      O���<�洞�I���A@7z�¤Q�V�E�&�n�V���X�S�s��ܞW�w{?Ocl}��Jzr�~�ݛ^Y�[�&  ���?6�+�0      �1�o�%��,�3�4}J� ��y�ĬR=��
`���k cʥ�L�K��~S�3ʫV]m��n:�KI=��$[�ҿ��g;  �X�?6g���      ��%;A��P�A�3z�8�V�Z;�#!<Ѥcs�	�O�� ��h�ލOڂ<��河��g�ʕMZ� ��g�쯗{�ɥ�J�c�  ��� ��      Щ|�L�r�G�4��'��g�ͱ��v�s��f�ֽ�\%��$�� 톁;������Y%����.������<6�J�4}�:&7"yo�&  ��R�]        cm�\�T�������c�Unu_�Z��܏�׮{�I�c� @;c� �	2��G�!]Q�_P4���s�b��d$M�`nG��c��s�   �Բ�       �,&i_��͕|:K�o���ʫV]���C|������P������ ���;�V1h�ťR���P�Jҹ����v�=�b𡡩y^�B����~   �d�      t#�^�#]vd�_��sr�&�\yw�2 �ʍ��E�G�#���4.v t� ZMb�HzA^*o���j���;e�7m�r�$�h><<��e$f�z��2M��  �P��.       �؞�Sʮ�d!�Nn��W�{����R�'��r١�����N��@+o�|���k��1�E��WʫW_kR;����Y��D6���  Z��y�       h���d�W^*4��
��ҷlժ����R�VwWQn��%͊� ݂�;�v���׻%��Czf�N�~q_��]��V&h+.��!<ۥ��Q;  @˳���	       Њz]:�d��H-�W��➾�o���9v��jCs�L�J�$�b'@�a��M���Dvd�z͟�4��p��o������Y�8�����Z���-�]�H��	   [��;       <�q&͗k~>R�e!���.�)��=��;x4�0j?\j<!v t;� �ݴ���׮[�����vYo�ߵ�+�;�����S���tP���'����  ����b       @;铴����K�S����L�7�Kǭ\yk�8t7aBM�?1;�\�i�& �C��$S$f��F�7�t�y�Ҟիo41-�ث�M�b��V�x�L���   :D7�      �V*K��]�&ҩY��.������S�g˗g���|������暟K&�vrE Њ��T%��4O�,�BX��~�nW�e�l��b�3x�̬\�Ǥ���bW��  ����       0*\�%-Ld���Bz�ɮro\ջz����<�	u�9���)�?��)�B h�t���@�z^d!��fW&ҕ垞��;Fb7�=���5J}�+J�����>�ɇ@   nҤ��|e	      ��L������%�Bz��W�ٕ��߷U�����R)�Ӭ8��r�9�z�� �� �Q"����4�ޝgy=�_���\�����Gv��bG�5���꽽�,�<��{��ޒ�n��c��   �D6cFs���       �i�dǛ��\�,Mo�t��kE��W�;���r^�<E*=���ʥ��b*Sv h�@*K>�d�L���{z��~$�������+V�����000�$ɳMz�d{��n��I^   Lߡ)�8w       x�k�����6��~�d?��k�(_߻�_�T�������)�Z�Y��Y&^.=K��Yu @�a� ��,�&�L�i�j!]-��nHT���$���wo��m�����SݓyJ|�\{K��  D6n�l��	�����?�.B���wo�A�      �̑|�d�Y�Pҿf��I~�����Ѹ�֬�/v$��K�l`h+5��}���g�SeJ,v `�1p��`RE�|��Ly��,To��涼��>�:[���حxd>{�����n��m�\���^��Gy ��J��v{��$�@���Տx�TpL���U����9+�7�       ��$�%�^�Z�'��]d(��j�n�]s�-�:�%��y=�����И������č�L������ �NY�]����Jd�%�Bz��~Q��"��2�u��ɿ��˳���«��yQ<�=y����溴G>R�L����  �̟�ҧ?%������Ȟ�<%G������쳏4iRs���        ��/2�K�x������~%�_���r_�-v�����-\*ժ��(�&n���\�=%_�fKT~h� �v�`����ܴ�iӈ�]��u�,���iyQ�7��w���r�{��wǚ����%ې�i��/��\�9���Үy�;J�ئ!;3v  �x�CU�c�J���,��������Ieh%v�!�;��      `,L�t�LH.w)�)��.�Z��r��I�5J����Xq�I���V𡡩y�s<i씘�q�]%R.�>N2�Iw� w {eI��k���$�)�ɕ��o�n3���ߛ��tgb��GZa+W�1r{4>sf^�tkTMɐ�g��Nn�S�Sv�swIƋ�  �VK�:J�H�͸d���8C��K���ǡeX���5����      �Y\�J��u�d�.|/��4Ϥ;\�{Sr���QH+���$�s��w�1��?�>}RV�0TR1T��.2��r�#Ӝ�ޘ�d��]b� �R� ��$��=6~D2%��R.)�zIwJ�[�5*t���q�{����XSO�{��Z[�j}Ŀ���3fl���gj9I*����}��x��r�!Y�����4N*����\�  FQr�a*}����ob;������C�ư�$Yx���ۼ����       x4=�v6�����q�`*�� ~���VI~������VܓH�5J�{�zz��o�sܿ���s������Y_}FR�'���w�7Y�K3L��M�SCŦ?������  ���; ��	��$�I����M�g*6�^^.\�LYH3I�$������L�V���}ĥ���䖻k�����Ö3I��E������Hz%��a���d���m�T��S2Q�rM�4U�)�ciJ.�˒T��9�^9��  �Y���T��}TJ�-�sm�=U����x��:o&�x�&)yի�z���oM=       �Uz$���/�����7�\�M7�7j�B��ɴVnk%_g�u�N�����Z"�wȓ�_��ٻ�(K������Vݪne��I�3�;�wΌ3�w&��(Q"q�F��hDp51nQ��ƨ��+₈��+Fc��(��ƨ	J#uouˢl�U�>�� *K/u�u��s��z��9�9�>�;O�6� �$7�Zo���a)�����a�/ex����z�R�\:90�Xk9����Cj�%9di�M��M�p�6����=�[�� �j�&�\�#v�u�0n���G?������x��an�$�S�s��5��{y_n�k�� �qS�s�̜��4n�E�aK^����L#�	�y�㓃^�K��;    ��)IM͡��)n�p��Uǭ���Ncx�1�s���3J���b�}�m ������ ��}�n>   �A��c�u�����#��3�p�Ϩax`fN>y��v�R-      ���  0Uʆ�]��:���7��t�+v&�s�����̪�[o��;      0��  �.7��q��?<�g�+9��=��=43�4x�=I�3p      ���;   S�̮�k��A��y�I�v�?�6f�������\�w      `��  0U�w�3�s��ϙ����=�1��Y=���N礓��pc��      3p  `�^���+�������.H9�ȑ���9�Iw�_��S�z/�      ���  ��r�5<���Gr|�W�*3~(�����V��SS~���\}ur���      h��  ��S��,����Fr~ٰa�K�~�H�g4:'<.3�M���T��      Z3p  `*կ}-�O|br�M��ࠃ2{�Y��������q��i������sZ'       4e�  �Ԫ��,�މɎ��`v63�~uf^��������2s���Lӎ��/����i�       К�  0����M�O>%YZ���N��k_�t�#��}S�s�̾���|�����	       ��  0��g>��S��,/��Σ����79�����)�7g�w'�:%���3�ԧ[g       4g�   I��(��>m�#��K�5���D������`|pf�>+eÆ�%I���ߐ�3       �3p  �݆�X����֑�Q6n������1�;���s�I��_h]�$��]��>�:      `,�  �m�����y#�g��̜��̜~z2;;�{�i��e�]�L��_l]r��g��'       �%�   ��睗��^6�{:'<.�g�����#��$�nf��?R���%�����?���       c��   n��mo����G~OyЃ2{�E)�����j��g��H9���%?Rk�'�pغ      `l�  �����v���)?�s�����y�s��?�����ޙr�Q�K~����~��3       Ɗ�  �����_��_4;��s������q�������?���.�1uq1����u      ��1p  ��08�5��_��]�L���I9�U�o�qDf?�����[����0�S��\}�      ��3�:    ւ�_���̤��g������ޙ�;ޙ���y�}���0��>3�=/��~�u�O��ͩ_�b���R���ԋ/��7�<��    ��f�   {hp���Z�yֳFY)�tbʯ����ן������kܾaC딟R���^��� �mx�Y�uV�     `uZ   �Z2xի3|��V�r䑙=��̼���ᇯڽkU���2{��rܞ��3x�3����%       c��   ����We��7�ꝝ�O�s��G&����kE9�̞����Z�ܮ��^�����       k�   ��<-�7�yu/=��̼����ȇS��Yݻ�\籏���ߖ�_�:�v�??����u      ��3p  �}4xşf�������?���~�̞~:���V�a,p@ʿ�w����f�5g$����nW����/l�      �&��w~  `���I��Γ���w���Rf��K�YZJ���d�����d��S��:��R��&��䚫S��&��U��c���a��zhr��~xr�a�����S��3�G��3��h]|�n�)�'?9پ�u	      ��`�   �i�?IJ'��?�M@��r�{'��w�]}�Ν�F�?�Ar�ɍ7�^}r�����v}|���u�'�oLv�L���}����7����KJI>x����ɺuI�rЁ����A'�r��'�xЮ�:h�����)���3&��E/N�ַ[g       ��   �/{YRJ:'��:���ͥlؐl�p�/��(�}2�������       kJ�u    L�Z3x�K3|�;[�0�w���=�u      ��c�   +��^��i�>�v����''7�к      `�1p  ��Tk���>�u	��������       k��;   ��Z3x�2<��%��������o�      �f�  �(Ԛ��^l�>E�7���K^�:      `M3p  �Q�e�~�٭K�����On��u	      ��f�   �Tk/|Q��~w�F�������/o]      ���  ��՚�^���i]����?~Q�      ��`�   ���^���9�u	+�^rI���u      ��0p  ��r�����[����2�'��,/�.      ��   ������\#��n0��3���m[�      ��b�   �m0�=r�`����?K��Zg       Lw   ha0��9�����.a/?�����       ��   Z2x��3��C�K�C���2x֩I��S       &��;   �4dp�F�k����tRr���K       &��;   �v�K��h��������n�      0��  `,/g�ԧexᅭK������      `�  ��2x֩~���%�F���^���       S��   ���rOyJ�}�u	Ir��<�����[�       Lw   7��<��~�Ƚ�n���NH���%       S��   ���r�<9�O~�u�t���,���ԯ�u	      �T1p  �q�{�^?��%�媫���Ǧ~�+�K       ��l�    �N,-e�I'��G%�3�k&_�~��ɕW�.      �J�   0�v����m]       #�i            ��;           c��          ��`�          �X0p          `,�          0�          �           �w           Ƃ�;           c��          ��`�          �X0p          `,�          0�          �           �w           Ƃ�;           c�Sk>�:          ��Vk>ޙ;�G��[�           0�j�Es��Gw�7��sv��>��\�:
          ��R��ͭ_�Ȳe�͝$)�\�4��=6��i          �t(5��m���r�;��s�H�~�	)9�]           Ӡ$�ݴ�w�%�,��k����A��{bj�^�<           ���f���'?1pOv��{'&y�j�          0-�y�~,�����{�{���#o          `J�wt��;nO�`��$%��~��I9stq           L���n�I%��g���=�e�����~��           ����~��;�'w1pOn�����׮\           S���{2nO�`������zϮ%��           S��/�������ɧ�����ދj͟�[           S䌹��s�tܞ���=I�{\S^��_          �t�)�����`o�n��I2�_xiIy��|-           ����>�_x޾|�>ܓ��_8��          �[�ԗ�����3��{r�Ƚ�Ӳ          ��QJ^����d�د�{�t��W�����9           �M����^��{�~ܓ���&%OIRW�<           ֆR��n��ʕ8kE�I2��9��          `J��rjw��g+u��ܓdn����rJ��J�         ����    IDAT �X�Iy����_��+:pO��Ņ�&���          L���g��^�����=I����ה�'��|           ��)y�\��(��=I��響'$Y�           ��AJN����4�F6pO��~����q1r          X�n��k���t��$���k�O�4�           Xq�Z��z��G}���I2���)yT��q           +bPS�0��p�j\�*�$���>��G%�y��          `��<v���պp��I2�������          `���5��p�j^���$�ݺpQ���Hr�j�          �]�9L}�|��j_���$�.^��2,�%����           ܮ���\�����M�I�ݺ��R;��;          �8�^R}]��?[4�'Iw�/���\߲          `�m/%�����n�t��$�~���F���-           S��Rr|���l���$����Z���[           �ȍ�S���z�k����=I���j���$״n          �ז�c��:�c3pO����K�zL��[�           L��S�����u�m���=I����O�1I�j�          0�~�Ny���[�����'�\�����nm�          0A~��9vna���=c9pO����o&9�&��[           &���S<�x�W[�ܑ��'�|����zTI��[           ְ��Ny�����Z�ܙ��'ɺ~�ۃ��J�k�          �m�Ù����:䮌��=I��z��<< ɖ�-           kEM�Z����~��[�Ě�'���[����I��u          �pE�t8�u�?��S��������oڴ��3)'�׭{   �T��S�<�u weݺ�w����9�� �ov��u�a�� �q�CZ'   0]�7����+��:do���b��MG���߻u  0:����9항3    `M�[�d���:  ��s�p0s��m��n됽�i�/����.u��5�T>          �*�2,�����'I�r����Σ����-           c�_�K�~۶�Z��5;pO����o�G��[�           4���N9�^o�u��X��$)۶}�����$_o�          ����f:G���k�����=�=r��yPR�ں          `}�۝=��+��Y	1pO�����;7wlJ�Һ          `���p�r�勭CV��ܓ�l���n���I�ܺ          `����zLٺ���!+i��������&�R�          ���ݒcJ�U됕6q�$)������1����-           +�\��cK�wu�Q�ȁ{��m�n���O��-           +���޼�貰pM�Q�؁{�{�z|�϶n          �۽����5�\�:d�&z��$����M}D�ϴn          �{�o�;wL��=���{�{�~���k���-           {�~������UW]ߺd5L��=Iʥ��;��G��#�[           �JM�T��yX���Z�����'I��7v�z�cJʅ�[           �HM��\'�Qnjݲ��j���2r��o���n          �I�䢹��GN۸=�{�{���?&��i�          p��|ln��G�-[nn���Tܓ�$�n�����Ӻ          �&�;`��˥��h����ܓ�#�^9�u          0�J򁹍5���d�����b��$�j�          L����{�S.�d�uHkS?pOv�������u          0U����W���!���}���n�����ٺ          ��=�~���1p��]#��g$���[          �IV����_�A�qb��v����J�_�n          &Q}k��prI��Kƍ���(I���N�%ֺ          � 5o������>�;1�뽰��i�          `Լ���{JIj�qe�~�{\S^޺          X�Θ3n�K�{`���Ғ���          ��SS^=���A뎵��}u���          {���>�_x^뎵��}/��W��          ���k�����^0p�K�~�եď           �PI}�q��3p��^<5Im�          ��R���~��;�"�}4��)5O��;          �[�yQ�����k���~�[�%���dغ          h�������i�C�2��4���֤�#w          �V5)��-�^�:d�3p_s���k��Z�           ��&��s��׵��+d���zB���-          ���I}�\����!���}����%���;          L�aJN�����:d����h��͏)5�&�n �iQ6oN����:    ֦��S����   k� %'��zg��4�#��y��Ú�̷n          V� 5�7��{w�Id�>B˛7?|X���         �$�Z~w~q���!���}Ė7��a�^�d]�          `�-�Z~{~q��!���},m<�?�d}�          `���5��_�:d������|P�ԏ%9�u          ��v������n2:��Ew���K��Z�Z�           {d�0�7��W��W�ҦM�)Orp�          ��TR�[���t�i��U����XR�K�u�[          �۵��>¸}��7����6�<$�Z�           ?��R���~�3�C�Qi0�vn���)�O%9�u          �K��]X���!�������6�Ǥ|:��[          `�][J���z�:d�uZL��~��SrL��Z�          ���6%3no��cb�ƍ�I)���[          `��0��й����:���cӦ_H��%�غ          ��2�<tn�_i�.����|����zTI��[          `�]Y;�������}̬���=(9�$��-          0��_;�!�_k+��}7m�p�����ܫu          L�mu�9f~���:����1�~��-�:|pR.k�          ���n�Ù���/�1�~q��A�N��-          ���d�v:�2��{�h��+��k�7m:r6��$�n�          k��N9z��¥�C�s�kD�ǽ6,u�?����n         �5�{Ù��뮸�;�C�k�kH=∟]���lR���-          �\>,�~۶�Z��g:��s�����]^~HJ��u          ��-������k���s��=�z�          S���)X�u��!��5�l�����̃����-          0f��4�9ꀅ�^��^i���?�s�.�L��Ӻ          �����٣��/�a���q�^�:di��'����-          ��7�Kݣ˕[��a�uZ�ʖ-?쮛h�/�n         �F����+��k��'D��=Z���hjԺ          V��wK�-��խC�^p���+o�./?<��Z�          ��(�t;����a�>Aʶm7vS�Orq�          ����l�ز�pM�VNi�ʫ�6����$Ǵn         �����7�Z���Z�����>�J���{���k���-          �¾�ݹ�8���d�>�ʥ��;��G��#�[          `e�/t�vW�����%����+�����CyLI�p�          �/%��.-=�\y��S�	�k�~�ǖ��n         �}QS?�-�8���WZ�:j2��i��I���-          ��j�'���Y�l��u���)Q�A��BJ�i�          {��|ܸ}��O�����Ssv�          �35��܁�e�>]ܧLI��މI�j�          ��Ԝ?�qãʥ��h���*�h�&ei��3�<�u          �������J��:����)U�������3[�          �n�3n�n�Sl��}�I}}�          �]9���`�>�ܧܮ�{�Y)���-          L��n��wv���z�Skɟ�n         `�Էu�O*ɰu	��s��^敭;          �%����b��-��1����;          �p5o��zO6n�J� ��Ҧ{�QM���          L����-���:���wnW��pzIy~�          &KM��v�ܹSK�6�aMyU�          ־�������`|�s��6o~n����          �]5���~���;o����n�wFJ����n         `�)�/3ngOx��=�s��SR��}         �*%/��z�h���`��^ٹ�OJ�o���         �����^;X;��k;7�������         p�jj�3��{m��w���M�NL�[c�         ���I9u����!�=���6�vIyw���-          ����g���oh��d��~ٱi�o��sb�         0�jR�>�￱uk��;�m��͏)5�&�n         ��aR��g��6wVĎ��|t)���         L�AJN����j��g�ΊY޼��Ú&�o�         ������{�n�d0pgE-o��q�N� ɺ�-          �Ԡ����ŅsZ�09:��,�[.*�<2�ͭ[          ����vV����M�~��\�d}�          V��Z�o�/.|�u�����Y�x��2�X��Z�          �"v������n�d2pg��6n|`-��%9�u          �e�0�1�����ar�3rK�6�rM��I�[�          �ɎN�o��zm�d3pgU,m����t.2r         Xs�������?�:��g�Ϊٹq�/�t>���-          ���׻��ŭC���L����K�zl��[�          p�n,%�����YUs���N�1I�j�         ���t���^�s�C�.�u �i����!5�Nr��-          ��kS�^�K�C�>�4�c����t>[���[          H��0�򰹅�/�a:���͛6�ۙ��k��u         ���a��_��z�WZ�0�:��n���oJ�*I�u   ���w�a������wU=U�=�g4A3��D��66�	�(la���8�����&�9��`��x��9�`���p c�<"h4���t��h���]]��+��骻���y�����5u���      ����f�Nn�d7�n�[K[S�D�         �!�������{?�;R� ���^����Q]��         `H쫺�[[�{��;"���2:9����#���-          C`���o1ng!�;ΉM���G�PD\��         `)����^�����ݹ[���΂3Z�{�Rl��{r�          ,A{�Z�&�v"/��`U���S�}(�zl�         �%bO�^�ed��{s������U��o������n         X�v���[F�����c�΂Wmذ�So|0"���         `������2:=}_�8�Z� 8�4=���uo����n         X��:��&�vw�45��h�o����         ��|�S�mk�'r���0pg�H{�<P��Q�'r�          ,_��k�,ۻ���*���U]uժ�ə?��o��         �@}�(��ݻ's���0pgQ������-          �g��nKey w�/w�jÆe�z��5w         ��"�m�ݾ?w\�Z� �Piz�X�#�ù[          �O��������<^DuGD|0w         @>i[QK��,z)w ̇��F;��O#��-          ����祃����w��41q��#E�7w         � }���y�q;K��;KFڱc�1��%)ҟ�n         ���bv�����#�K`�������g��JQ�I�         ��������������g�^�})Żs�          ̷*�_��s���Gs��|K��_��zg��ߍ*^��         `>TQ�y�V{q��8�����,Y)�[�ۯ���         �bU)>�l6�4ng)3pgI������{�[          .T�����i׮��[��R� �*��ٴ�7#���[       ��+�ĉ�?-w��FĞ�LT�ʝ�MQ�+����8p ��org  �0)�76n|yڶ������; !E�����Φ�'"�͹{       ��/zA̾�U�3.ء�?����G�3�;%""Fǖŋ��uqb�չS�{p��; ��"���q�+����QUe�-�M��"����      `p��c|ͺx��+z k�%�7�K_���j���  ,
�h��W��=�;��; )ETE9��H�˹[       ��7�k����q�e����1��7�ո �s�?����a��P1pg褈�h��)~)w       ��|Ūx����^�����ħ<#^��7E�52� Xl�oe����#w�R�����۪*~>w       �U4�q�]��g�����W����ϻ3�{�K�V3�  �l��,ʉ7��^����&�Zk��3UĿ��      �`���7?'���/�z�޷{��V��eo��~�M}� ������,и�af���k��UE�7�;       ����x�k�c˖��٫V���|���5�>v�� `	�����;DDD����)�O��       `�.���x��k/�0ogn�lK��M?���8og ����b���)��������/���e�       o|�%��������_�Y�?��׾9�-[1e  ���,�o6n�����e��)�?��      ��5���ޗ�!���g^�倫�۟yK��%��FQ�s  KQ��i�m�Exw�E���"�?�K(      ��S����8�{�K�V������x�_7?���R�c!  KE�/�ʉ��w8�f��_"ś��      `(=�)ψ����j���g�Ɩ��_���'<y e  ,��˟����;�F������FD/w       �w�5�ū��#�j����̺���~��eW\9�2  ��������4''~#��      `X�[i����o��߻���Uo��X�j<C  �QJ�3EY�������Y4ˉߌ��F�       CillY��5?��������x�+���H�2  �T�O������; �fY��̦M'R����      :�z#^�=/���blly<��ȝ ��QE��VLN�r�Xu�����3�6�R�?��      :)���gݖ; �ť�H?ڜ��s��bQ� �I�,�Q�xEDtr�          ZQ�H�4n��a���n���;         pU��'Ͳ��r��b�� �Q��~����'zU�qD�r�       �[�_�C����` Z���N  X캑�����������.P��~������ժwG�H�      �~JG�D����@q�P� �Ŭ)��l�?w,V����5�&>��tgD���         dխ��:�v�8�p��ɉ?OQ}wD_��    IDAT���         dѭ"��59�C`�3p�yP��_���܈���         `�t�*��*'�G�X
�a��{�.U��Gđ�-         �@�VQ�՚�xw�X*�a��IQ=/��        `���E��VY�'w,%�0ϊ����s#���-         @_���z�HY���!���Ce�����D���-         ��:���c�,ߛ;�"w���䶈궈�?w         0/��/*��r��Re�}�,�OG�gGā�-         �E9�R�Q���K��;�Y�����F��s�          �X�����s��Rg��l�?WU��"&s�          ��PJq[11�7�C`�À�&'�Qݒ"��-         �99��������!0,�a�Ze���C#�v�         ���Z��91���!0L�a�F��+�Zښ"&r�          ��@T�ۚ�����2���g�׽)"ݗ�         �&��Z��9��S�C`�C&�SS��Uwk�ؙ�         ���}U-�ښ��|�V������nUm��{s�         ������[[_����2-�=sQm���[         `UQMU��-��_���������[t��"�ݹ[         `��j��ZSS6|� �����*�fo���_         0{z��֑���C�������.��n��/�n        �%nw�[�:�wｹC�����4=���uo����n      ��R��F�; ��۝�:2�gg�����������͑⓹[       8�Z�W?��q��-j�z�  ��=s)n���/w�H�@�={(������[       x��يko��X9�.���+�J��rg pf_����c��D����aK�v=X��n����      ���Y���1�|�7��j͆���'d� �,�ҩ׶�ML�s� ��� �Yڹ�Pu�U�휜�@D<#w      ��[�bu\��o�F�|��.ٸ%fgN�Ԟ{�񵪊81�H[��E��y �S�RQ4nm��=�;83wX�Ν��n���7��      V+��ŕ�?5���O.6m�.:�3q�Ԟ���UU9>;��ڲfԛ��� ��|��uoK���s� gW� ��4=}��ͽ0">��      `��py\����q��uW\sC�^�q U  ��g��������a�0p�E$MO+��#">��      `�l���r�#�s�Z���Q�=9��\��2  ��3E�g��<�;8w�Ȥ�<^�ҋ"�r�       ,u)����'��+�?�߭��q�c�#c��P ���mE-=;����.Ώ�;,Bib�D16zG�xo�      ��*�j��<9�]��>�Q4�17<#FF��/ ���>U4j������K��g��Tڱc�1��%)ҟ�n      Xj�"��o��u�.��fk4���7EQ�P �Y�}q��iϞr� ����}�lc|�])�{r�       ,Es$���;b����v����O�Ψ�L5  ����������s� Χ&X����K7ܕR�;w      �b72�"��g�貕�~��K��O��H)���  TWtf��8���8����K۶u���:�6�^Dze�      ��h��5q�c��Fѷ;.�ty�Z#1;s�/��Z�j�gO���}w�� �%��s������N.��;,)�[��k;�7���W��      XLV��W^����}�k��u}�#"�ı�Ѿo W dSE��T�3MO���̏Z� `���n�n�>"~/w      �b�v�q��Oȸ ��S��@����41a�K��;,1)�[��7D���n      X�6\vMl���H)�N �<T�oŋӮ]'s� ������+��#��r�       ,D)����c���N �<U�k��~�q;,M�D���(�o�H���      `�_�)�n�"w  �)U��_�v����;,a��'�Q�J�      ����v�/�˝ ��ygc���m['w�?��=4r/,R�R�      ��db��x��d�  ���,��+S�\����a����n�����s�       ,UUŮ�|&�>�; �3��GQ�_e�����Hk��3UĿ��      �P�zݸw�'�ıùS  8��[EY�:Ets� �a�C�U��U����       X(�s���ŏ��̉�)  |��7�r�RD/w	08�0�Z�ĿN�~"w      �Bљ=;�����ur�  Q�+���a��Ð*ʉ_HQ���       ���G�޻?�� @VU�z1��a�vN�0Ċ����?��      �P=t��ʧ#�ʝ 0����͇���AC���\Q��1�����      ���x��d����  C���������e�D�n��H��0r      �����cj�=�3  �F�/�ʉ��������f���Q���^�      �s12���痻��O���  |}�^�D�`a0p��99��G�#w      `k���5�����ϊ��X_��s�������z �0KQ��q;�p��7i��Q�)��     �&��7_�?��X9�.j�z\q��zgUU��˟�c��� �a�R�lQ��6w�����,�߮�zUD��n      ��]�2��g�eW=.j��7��r|}����׻{�n�{�'���}� `��*~�h��}�`�1pN�U�o7r      r���q���uO�)Ɩ�>��\~��Q4��1י��?�ٓ}� `TQ�ۊ���,L��i���U�WFD'w      0|��Z�?����+���N?qh��|�c��3{�x���ǣ;���
 p����c���/�.w��Z��;��#w      `@�"�x�q����e��;k7\+����,�ıñ��OF����. �%�����,'~%w���g�j��UKqgD��n      ���K6�㞺5.ٸ���kn�Z�ч�ov����뫟����w ,UD��fY�j�`�3p�I��~��^'s�       KO���������D�h]�͑���k����_��_�]  �\/�zc�,-w�8��11�g�Jw��;      0�.ٸ%�ԭ�z�Ƌ>k��bl��y�:����bz�ށ� �Hu#��e�;�C�ţ��XR�ɉ?�l���U��D�h�      `�]�"�x�l�����R�-��_��G��z�v���;j��7�g��������Q�����)�7s��@  N�U��Y�� w����(˿�l��yU�z_D,��      ,.)�b��bӖ�D����]�2�o�*�'v��٧�w����>t�'g�r�ʱf���� �<t�*��59��s� ���J�B15��=?"��n      ��+���O~Vl�����ۿnӖ���X���f���h�~  N���]�����)�`���GRTF�      �Y�델���ǵ7~G�����}�V�+�����|��n�^5��j)E�n� ,(�UTw�&'ޝ;X�|�.JQ�MQ=7"��      ,L��l��>uk��teD��ݻ|��X���1����ZDfL p���{r� ���;pъ��XT�["�`�      `�i�(�#Y�������������c��KZe���C���'`^4''�ET�E���[      �����=q���Y�7������\o`w���� p'RTw���{s� K��;0o�e�鯍��n      ���|>z�n����m��k7��������{J)���@� 8��)�e�W�C�����WͲ�L�xv�      3{�xL��j��/��	Qo}�cv�U5��{��"y� ��xJqGQ��,-���k�۟��޳����-      �±�}o?z(��Es$6=꺾�1�̸="��0�  �:�R��h�?�;Xz|���59����Q�n      ���b�W?U��r��K���k�v�l�۷��U���v  �C)�mE��׹C�����VY~���Ƚ��      XN;���e�=����Z��A��^�v ����-���,]�@_���W���5EL�n      ���_���ǲ�=2�<6\��y?���EUf�^K)�5/� �`����v�s� K��;�w#����7E�\�0       H�׍=�|>��/�&F�V��ss�{��h�{  �@�j�7'&>�;X�|�btjjW��n�;s�       �y�@�?�7��)�b˵7FJ��
�L�;og���; 0`DU��9����C���00�����U�5"���      ��޹=:�3Y�^�b<.��Q�v�\�� �������jN��T�`x���hYjkD���      �57׉��۳ݿ�Q�E�5z��t{Ut{�y(:��Rus ` ��n�����r� ��'`���ro�)n�Hw�n      �z`;�?���z�W<��G|����ɓ'�СCq���q��ј��=�9}��^��v 0���^�����/��O#w 0���]S����t�E����      ��{�c��K�^��a���_�)�O�����w`|���u�"{kd$6��$֯��W}�띹���Q4��������^���T��@^p�I��M��-�O�      ���9������^��f"��������8p��S��#"fN��={'�S۶Ŷ�|6>�s݁�S ���V��M��)�v �z�������׽5">��      �g_�+�>8�;�?���?����#����݃��?��عsWt:�{��Q7�  �fO�^�:21�#w0�|��KSS��F���S�[      �\��s���f,~��}��w�^��7��h4���RUq�Νq�ί�����Z�] �������<�wｹC ܁!���@�l�U|"w      ����Gcj �?v,>��?��G�|��G���H�7 �UU�`_��}�|&�R�0�  �bW�׽ytz����8>� Fڵ��b�u{D|<w      ����{���#g������/���8z��#�W��cdt�y�W������jǁ����x:� @|u���9:5�+w����,(i��C�H�9��[      ���z��s��#����_��s1=]�����eQo�|^�a�{��nw�b�Ψ٨��l `(}�S�m��h�x8w`�I;w*�s�E��      ��������~n�Ӊm��Ynt���Hg��^Q=l�ߙ���������R4�f ���rQ4�.ۻ�?�x�>� R��>V��^��      ^yߗ�3sr^ϼ�ޯƱ�G��s�z#Z�cg��^��W��OOFu��_�F��z� :_*:�ִ{�d��S1p�4=}��ꎈ�P�      `��ݹس���z殝���϶F�G�^?�Ϝj�ޙ��ѣG�7�
�� ��ET�J�wM�8�~�-���"�E�_�n      ����x���<,ZUUL��u�?�R��e+��3�ީ_T?����I;'͆� p�>S�xv*��C �ħ`�Key��#E�7w      0X{��Bt�:}�ɓ'b�3s^��(ZQ�FO��S�����f�I)Ea� \�O����nߟ;�l|���c�Lc|�KR����      Ngv&���}��?z�~otlE��#�UDTq�������)�� �PIۊZ�-ML�����w`�H۷�6�W�4EzO�      `pL�#�.�ѹ|>�j12��_��N��{��]�]���z; p���8y��v`1�	XT���K7ܕR�;w      08{��\TՅ�ǖ-���m�F�Q���k����F�u��]�F��� ��h1;�t����! ���XtҶm�F�}WD��s�       �1s�X�8v�tlY�t�C���+#��gطG�l^�=��,��z 0�G����ҁ�(�L܁E)Et��|m����-      �`�2z�ш5k�]���j�}��^Q����/��GܛR�k^p �C��-:3�O��͝p!܁E+Et�v���{�[      ��]�2���E��+����o�.�z����oO�b��5u��� ��UQ�E���ہŬ�; �b��nU���ٴ������      �c՚}�Տ�.>������[�:�N'�4g�߰)��Ϻ��U�^�z��^p�=y"���=o- ��VE���f�δk���- ��X�RD�k#�����=      ��[9����X�v]\}�u��/]��Z=Z��i������K7_����ı�Ѿ/w 0U�l5�׸X
�+`IHUQ���~5w      0���F,[�z^�z�3n�z�?�^yգ̸ U����F_l�,������}�կ�n      �ϊ�u���LV��gm�}^�z��+VƳny p&��w5/�xgڱc&w�|1p���F��E�_��      ̏Uk���y���	q㓞>o�5��x��7FG���L �s���d��i۶N���d�,9)�j��o�R���-      ��[9>����g<sk|�M�F�tQ�,_�2��e����o 8�we��)b.w�|k� �V���3�n�?��      �0��VF����Ox�Sc�������U9|�~7�W]����cdd�/}  ���^��1n�*w`IkM�vf��z��'s�       �o՚�����QW�e�o�/~�3���o;�нV��e�o��>�;c��M}m 8��)ʉ�O��! �b�,y�v��f6o�R?��      8?+��;p����q㓞7>�iq��}�g׽q�Ѓq���9˖��e˖Ǻ�����*Z���( p�(����ہ���
�v��g6m��H?��      87�z#���k/Yk/��� �<��(ۯJ��! �V� 0(����*�/��       �͊�u��i 0�R�*��+S�\��A�)*�r�'"ү��       �nո����R��1�~�q;0L܁��"���xkD�Z�      ��V�1p �W��O7�̸6���yh��~KT��[      �S]�2��H� �,�h���<m����0h��PJU1��'Q���n      i����!U��@s���I;v��n���Z)�WL�����      |���� �P�Xsn�i����! ��C-Et��կ�R| w      �z��V���  ����iz�X���܁���o�mV�K"����      D�_)�4  C�+Ew�9i׮s� ��� @D��<^�<yGDږ�      �ݪ���  ��N�vK��ޗ;`!0p��t���"zύHw�n     �a�b|]� ��H�nw�e{���[ 
w��Iey`��G��r�      �0]�2����  �p����>:=m��0� �blb�ݫ�۪��r�      ��Y9�>w � ���sZSSw�.Xh�Nad��{�V�="��      �d�w `ɛM�{i�,?�;`!2p8����R-�3�[      `��X�r<w @?���.��/s� ,T� gPLL�M�k#���      ����"%S `	���[��;sg ,d>�E�,�)ޒ�      �����s'  �MU��7'ۿ��`�k� X����ټ��T�O�n     ��j�����5י�ٙ�/��Gs'  _���e�gsg ,� ��n�tg�e�#�7�n     ��ft��h�Fv��{��/v 0����5��ק�*w�bP� �X���('~����r�      �R�r|��*�<�`� C��Q}_����X���1ל�����L�      XJV����ؑbn�3�� �a��+�:ߓ��x������<�����+    IDAT�E��'w      ,�z#���}���] ��:؋��Ҿ}ӹC w��vz��Gă�[      `�[1�.R܄��� @_uR�����Wr� ,F� �5�g{�j/����-      ���_?��:�3q�衁� �*�xc�n8w�be�p�ɽQ�P�      X�V���]^o �)����d�rw ,f� �Y��UE���      ��ht��h�Fv��; �?��v��� X���A�,*"ޙ�      ����vWUUq��� *]\��)�����̃Q������[      `19v䁸zOtfO����G���l�� �M���ꮴm['w	�R�� �T���Ֆ-�3י�DqY�      X��?��?""Z#c�j��X�f},_�6R��w�=�o^� ��#U7�(M��L�<1p�Gi����M��;"}$"�r�      �b2s�x�k�}�Q��cŪKb���r|}4[�}��� ����R��1����C �w�y�,�O�l���T�;""��     �Ũ��ơ��q��tD\���s��8~�p?R�a��5����� Xj����n�����OLU�T�      X
.�u�C�ED��P `X�n���/�# �"w�>i��?�ٴ����+w      ,%����: X������ K��;@�����̾�S4���r�      �Ru��ݫ��#ȝ	 ,��^�δc�L����������GOl����Z��qI�      X��u��e+cl�����f. ���Q�^�����X��7� �W�SS�RT/��n�      6'�������  ��?ܜ�ܖ;`�3p��,?���W�;        ��◛����� � Ҙl�_)�rw         ��c����"w��0p�Q5:�o����n        ή����k/M۷��n� ���?�K��q(w     �o��>�����sf���B����=��@�`K����_k�K��իz�Zl����K�բ�zY*
?�FE�&��$ �$�	�YB 7{sΙ��fI6�ݝ9s�������������y<��u%����k�Ȝ����  �1ZQ�������! ���`�m���<������-        ������~��� ��� ��~��5�+�;        �GR�>��}cv�42pH2��,">��        <D�[�/�� �V� IJİ�:�����        DD��:]X��c�! ��� Q9p`�U�'#b��        S����/.ޖ�0����{�������        S��s��˲# ���;����_^�^��        S�v��4; w��P"Fs��OF���        �2���3?Z����! �����.u���f�        ���Q_�ei�]� |��;�i/.�X��<�        �B�����wfg �����\������        h���v���]�73p3%b�Z�qov        4�r����?��73pC�z�n���        �L���z�[�+ x8w�15��}oD�Qv        4I���v���� ��;�kϵ)"<)
        �D��J��Q�[ xd� c���s�[?'�[        `���K�(;�Gg�0����ZJ�,�        &Y��{�^�� <6w�	0��&"���        ��T�877�� <>w�	P"F����jv        L��(�'ʞ='�C x|� b[�۫��Bv        L�R�es��-� �w�	2��}[D�3�        &C�q��{Mv '��`´��/��}�        0�����K�0;��g�0aʞ=���/����        c��K�..��� ���L�v����zqv        ��q�\�wiv ���`B�O�xiD���        �1s߰ċ�# Xw�	U>RJ�����-        06j�d[���� `m�&X�׻>�^��        �F\5�ػ,���3p�p�'^��;         �}�/ʎ ���L�r��R�?ED�n       �45^����fg pz����]Q/��        �5⪹��e� �>w��h�8�����        �M��0��eG �>��>|dT�/fw        �檿���ߟ]��0ph�������        �M��v��G� �w���m�_�ew        �[����)�� ֏�;@Ô�{�įew        �F�Q^1Ͼ�� �/w�j�zo�(7fw        ��}nn���# X� T"F5F�%"��[        `��Jԟ){���`��4�|������        XW%.n����� `c�4�\��""���        �uro�֗eG �qf� �8��=>�q�k]��     �d=��x���eg�	Jݚ�  ���J��eW �q���������{j��n     `r�3ό�mO��`�f' ���d��Kv �� �����"�hv        ��j���Q�C �X� S`[���D���      �t'��Ǐgg ����^�s� l<w�)1��:"n��      �I��Ç�7�..y����s `jԈ���y�;L	w�)Q"VKԟ�i     �S��ww\���Ž���6t����oϝ�Y 0%�/���?���a�0E���'"�]�      0I>��O�;.y}{��7���������8���$��T��\�yv ���`ʬ���x0�      �]�5>qõ���]���a�|8Ɵ]������F�^� `u�%��h���;�����uK�Wfw      �8[YY��\�����>�����1���V6� ��Es����# �\� Sh��zUD�;�      ��G���+_�������>���u����6� ��W�Q�Wv ���`
�n�x��߳;      `���{�o��XZ������^��5}- ��o�~�Pv ���`J�/v��F�Pv      ���v.�~��������8����?� �Vuw�߿(��� Ӭ/��av      d���M��>����bu08�뭬,�{/k���ס �O)�K�jv 9���|�������      Ȳ��W��mq�uWE�uݮ;��뮊�?pE�F�u�. 4]��@���Hv y��\{8���r$�      6�ѣG�mo������7���)���7���v h���h�ײ# �e�0���ҁRꫲ;      `3�����5��۷�������7�&:�����V.��g���
 r����nDl���     ���+�ş�������m�=�{0.{�����wn�=`�<�^]�?� �3p J�{<J�Fv      l�������_+�˛~����w^zQ�z�_n��`ܕ�//,ew ������h�zQ�I      �4�Ϯ|g\w͕QkM�X�?��q�uW�v ���?�j�~v �a6; ��P"F�R~�ָ>�     ��Ӻ�p����X�Q�Go�P�gl߾#;'""��q[l��������Ny�r�� �L���J�{<���P� /˝��%�ew        0>�����D��C ��  �L��?�        6A��_1n���&����#���        4]�x{q��� �w f8�,"V�;        h�Rʯf7 0~�x��KKwG�7fw        �L��{ڽާ�; ?%; ��T�o?{К�3"��n       �Q�u4���{��bv ��	� <�r�=k��fw        �4��v ��; �jn���_��        �1����� �/w U���K��dw        �o]Z�;;��U� o�쳟8h��gg�        0�V�u���..��`|9���T<Zj�:�       �IW/2n��8���U�9�	��ٻ"�of�        0�N���3�u��� ƛ�x\ei���U�        L�d���p�; '�v:�V"�,Q�g�        0Q��W�(,e� 0����I)���Vī�;        �0%�h���r�; '�>��g���Fę�-        L������uqqov ��	� ��r��5��;        ��R�v N��; �d��k#�hv        co8*��� Lw NI���gw        0�޽���rv ����S�����       �8sz; ����S����F�K�;        O�������; �<� ��hf�#b5�       ���*�� L&w �d���wFğfw        0n�����'�+ �L� �]�WDD��        `|��rz; kf�����z�Ԉfw        06>7�ؽ6;��e��i)%^��        �x�%�o��� L�� ��[�t>Q�?�       �T�����]"F�! L.'�p�J����        ���1n�t9���V#�`a��Q��- �T�_��/G-�G��m�z_D<Xk]����2=iT[O*Q���Q�������xzD̦�W      4@�X�;�)�ݻW�[ �l~��i+ueT^��!� h�k�[�����`wYZz�t/Z/�����=�����@D�ӈ8�k     �L+��������;wn������- @3���(��ZW�����k�`��Y#��9������k��������     h������ʁK�! L>w ��r���W�; ��v�D\5�z�|�u�X͌Y޾�oGk����#��     �1v�\���# hw �ͱN���(wE�lv 0Yj�b+��ͮ�\Tz ��[Ո����+5�gD|gv     �x����7gW �� ��Ag��� `b�Z^ݞ�7�n�xv��t:��F�͈���-      �ʍs���gW ���  ���.�  ��G�_l�������k'e����������U�#���     �L����n �Y����[YX����=� �x�W��ܶ~v��睷eee�WK��[�{      6S��������k� ���p�; �� ��tg)�����i¸="���sb���ߣV����>�     `s�?0n`�9��uW�����c���(۳[ ��P��wvv�gʾ}_�n�(5�v�|I����hg�      l����^��� ��	� ��r���7dw  ca9j�o�~�G�<n��(un���R[��D��{      6T�ˌ��� l����G�Jv �j_��Gs���f�l������W�+J|,�     `��R� ��f2p`C��{#껲; �4��F�'s���C2����[�D�y     h���w�_Ȏ ����8��:; HP�3�߿��ߟ����q��l����g�      ��Q��e7 �\%; �f[�t>Q�~v �9j�k��+KKf����//%^��     ��������av ��w 6V)o�N  6�M��l~���Q���;      NW��f�v 6��; �}���#�� ��ĭ�V�7�폮��{iD\��     pF�:|Kv �f���*���wew  j�j���t���C�Y����_XK\��     �5ꇶ..��� ����p%��� ��9Z�������C&Aٵk0��raD�bv     �)�- 6��; ���҈ �ċ�o�Θ$����uԺ0"�e�      �����9�ώ ������7g7  뭼y�׻4�b�߳owD���     ��U�\Rv�dw �|� l�و�F�rv �^��v��O�\����     `2��[� �� l�������  ��0"^P��c�!���|�JD?�     �Տ�/.ޖ]�t0p`Ӕ�o�n  �C}�\�svE�Ç����rv     �c���� �G� `zԈ2�,|%"��n �l�=�~Nٳ��&Y�,\�<�     ��ߎ��v_ 6���4%���dw  kWk�e���7j�E�rv     �Õˌ��L� l�A�["b�� �A���-vߞ��D[�ݯDԋ�;      ��7e' 0]��T�z�n��&� 8u���*5���VKyUD�dw      ����s���+ �.� l��f'  �춹~���M����F�K�;      �Z���Mg����k���gw  '�Fyy�ew4�h8�����     ��Օ+�# �>� l��gω��2� 8i{��]x�	�,�+"ޝ�     P�~�8�����1p E��wd7  '�F\Z�*�iJm�5�     ���� �S� `:Ո��N�[�l�n �(�s����gwL��Z�,�;�[     ��u�}��9���#�! L'���DK�� ����q��*�Q�wfw      S�}�� d1p O���� �q��,;a*�Zo�N      ��(�M i�H3��~:"���  Um��^�1���ٷ;��     �8<��dG 0��HU�x� �V���ݻ�]1��G�     �)T��e��� ���; �j+�$� xT�gL�a�     l�2tX! ��H����JDٕ� <\�֙�ÏDD��      �G����ӽ1���f�@�R�'`�ԹV�Xv�4+KK"��;     ��1��1�� `���nvv�1��  �����ݛAܒ      L�0�HW��]�'��x�=;����      l���z��eG ��; c��'�  x�bX=F�     �&���n �w ��j�ueD�� ��F��c�      ��D}ov D�0&�u������ �kJ��Jv�Z���      L���~�s� a��)Q<	 c�����"J�,"�gw      W�=%�fg @��; cd؊�d7  _3j��n�|/     �Ub�PB Ɔ�; ccK�����;� ����9���7�      �����gG ���0Vj-��qp�S�Ǉ�     ����J�0� �����RJ5p�|5<���Uw     `ôZ�+� ��+s������ �r%.�`&;��+��     ������>; ����S��� `�<����J�3�     ��*W�={NdW �C�0vʨ��� �v'VW���E5p     6F-�F��c��ؙ]������ �f���	���I�     @#-�-/_� �����S"F%�� �fefƨz|x�      Xw5���С�; �[�0���; ��;���g��="��     @�Z>��  �����47^�� 0�Z��n buf��     ��^��  �����T����?�� �iU��B-�9�     @��[�fW �#1p`l��Wg7 ����	�     `�k� ���0�F�w �R��5�dgL�Z�oe7      �S��0��[�K�o��}� 0����}��gGL��*�0�     h�g�m�1; ��; c�~(�  �Ui�~ �a�:��fw      �R"�/wܱ�� �����Vk�+�  I)�e7L�R�     �uWK\��  �����6�|��1�� �iTk���sc�Q      �n�:smv <C �Z9|�HD�Tv L��;����iT�������     @�ܾei�]� �X�{��k� `j�яg'L��O�pD���     4L��� ���0�jˇ+ H�S5b6;bڴJ<?�     h�2j9d��g���k�z���~v L�s��w���iRw�<�Fa�a�    IDAT���     �q���ԏgG ��1p`안ZK\�� �j�r��f�F�!"�;     �f�Qn,���� x<� L�Z?��  ӫ��z�y۳+�A�(�fw      �Ӫ��� 8� L��p��� �b[Vګ��1V:�7�     h��
�0��[���{�; `Z��?W;��fw4])�f7      �t��}��� 8� L��N �)��ՈgG4�`ǹ?5�'�     h��e׮Av �w &�We@��%u�γ�;��F�ZF�+�     h�V�n�n ��e����z}v L�����#�h������     @3U�
0AJv  ������q^v L�Q���z���C��>�igV�_�����     4��~��� '�	� LO@�V���1�����¸     � �ƍ�� Lw &K�� ������?��+�(J���     ��Z�ސ�  ������Z��`��;+��wggL�z�yO�Z�>�     ��[ &�_�0Q������]� @�G���Yg=);dՈ��������     ���o/��lv �
w &O-�,�������eGL����/�Q�]v     �l5��1�� �Sa���yv �?������I2ر����Wfw      �תac��1p`��Z?��  <T}�r���+&��9�>����"b.�     �3����S� �TՈ2�,����[ �o�������k�C�ձ����_;%���     `*ۃ�����f� ��p�; �D��/�; �oҮe���;.�Gu���gk\��     ����q; �����Ԋ�)� x�3������}�!���s��Z3�Eĳ�[     ����  Xw &�a 0��RK���;v�Xv�8Xޱ����ѧ"�;�[     �)Sm+ �L� L��'n��Qv ���K��������L+;w��RZ���e�      �g4Sn�n ��0p`"�Ç�D�۲; �G5�^�����z���Ͷ���L�����     `*�;��ޑ ka��$�*- o�D}�`q��O��gd�l��s�֕N���ؚ�     L��Q�; `-��d� 0��o�o^^Xx^v�FZޱ����ED���     `��Jܔ�  ke��Ī��c 09�\j\��Y���N����Tw�ܺ����Ki}6j<7�      �+� �V5�:�Fę�- �)y�D�?������q����V�^Q���     �WF���,����p�; �DԈؕ� ��'Ԩ�=�,|fu����+߹�Y�@+����    ��R�d��$3p`��(��n  ���Z��+��[V^P#f���J��]���Q�%⇳{      �ԛ� �t�0�F� 0��#j\2�tnY�t�s=�'e=T�����N�GV:�(7׈�ED��     x$%���� L��N�9%�m� ��:Q">0�z���ה]��۟�w�����?F�9      ����?kw�7dw �Z�0�jDk�Y�?"��� ���������l�#Oؿ��a�z�3��|����*���Eĳ7�^      ����g�={����2p`�t>ߛ� l�ۣ�Ǣ�/���Wk����}%���E���g���Zf�Q�5�/J\3�     ��J�5�띟� �c6;  N_�9���txv�xvD�3�Ġ�p|%⎈��Z��R�h��/j<%ΈZ�X�<�~�/gEķ"�����j��o     �J�g� �t�� ��Z��T�7�D�����-�v�;     ��Ů� 8]��  X�>       �bC��3p`��<swD,gw        d���0���xe��bv       @��+,ew ��2p�!�b       �^��	 ���f���	        iJ�N �� 4B)���        iF�v�F�� ��0h�vώjv    0�f?���'<1;cz:�?��f�  ��+e�;� �C� ����Y�jD<%�    �\�/�q��S��yg�waԥ��  �d�v�3J�,; NW+;  ��m�     ��r��1�+��sNv
  L����h
w �z�    �2r ��S"���  �����(Ň5    �	e�  k7r(  b�@c�Q��    `�� �ڔ�P@ ������F�F    �pF�  �#w �������u#���     N��;  ��Q{4�Rv �w ���      N��;  ��{��҃� �^�hw    ��0r ��WG��v ���F)%��n     `�� �c+��Jv �'w eT��     �/#w  x�8�F1p�Q��;    @#� �#k��V�F1p�Q���^�    �PF�  �p��� 4��; �R>��;     �F�  �M��O~��� XO� 4�'�    ��  �aOٽ{%; ֓�; �S�    ���  "jT	 ���Ʃ�ܙ�     ��3r `ڕh��8�� ��j�%;    �j�E���+�Ny�3"�������������/�8pp]�  c�T� �8� 4Ni�;�fW     �l����#;c��>7f/g�S����}ֳb�����.������ �q6��	� 4N+;  �[{u���     ��zk������u�v9���y�Q�9gݯ  �g��n ��f�@�,-����     <��;  ������� `���8%�FD7�    �Gf�  ��r��� Xo� 4�'�    Ƙ�;  �6� ����ڟ     �c3r ���� 4��; �T�xJ    `� ��'��P� 4R�2    ��0r �SW�m �d�@#�yJ    `�� ��E1p���h���p    L#w  8y�(� 4��; �4g�    0��� �䬎V��@#��H��?��;     8uF�  �ꖧ>�� ���+�d     �6F�  ��-�w�dG �F0p����;    �����?�G�����������x����  ��J�D �X� 4��;    ����|>V�w�Ɯ���gE9�����  �����ޝ��Q�y~�����8�	
�#��h�O���(a�M��OQt$�(�
�H�	�� 2���8"�BP6���	T���q�k�Tw�r��奞������C���iw ���; �+e�    ��~�(&�ܖ�{��G @�%� ���; }+��    �E[K�  �s2��[
� ���%O�     �H[J��
w  zOf�; }L�����6�    �����D���  �J�w ���; }+5lp    �Ks�U7�,��  �yU{ ���; }k�s�<�    `�R�;  ,����� �-w ��#�4"�f    ��Sp �o6�; ���; }+�("��s     ��� �E+��X� �]��s��u'     ��)� �s�e���\�! �]��w
�     ,��  �] ���; }.yR    ��� �{t! �k
� �;O�     X<� �=� �5w ��'u       @�Ȓ. �M����<�    `Ilp �Ǥ�. �M����h�ug     ��)� �cRJ� �5w ��'u     ,��;  =��'��  ��@_KY6��     t1w  zL�rn� ����kMw     �D� �^�@�Sp���V�]�     ,��;  =&��. }M����ܵ    �)� �[Y�@_Sp�������    X<�v  zMf�; �-�;  �ӈ���=_w     �U�p�f�ZkE��J�1:���#=�@�)�.Wz5{ ���; ���~�    �X
� ]+�l|䧟1bD�Q:�O�b��n���$@+��w �Z��  �V?<?"ʺc     Х���@��#"F����3#�tӺ� ]ld�3ug �vRp��e)"��;      �t�ܾ��;�bR�_w h���  �"bt�!     �B6�t��/�/�Bɽ��G��n�;�4|xd����؈Q�#VZ)���{䈈|XĘ��uw�"�>����̋��ܡ�?�HO?��EQ��Cg<����# @;)���RĳY�!     �NRp�^��ȶ�.b� �����Q~�{�5�~���w�䞭�nd��6�׾6�ш��H���"�����6�8[�'����+׌Xu���X#bܸ�{�H�=���{4��G#=�x��n����U�Vf�b ����^ 0����     ������e��m�h~�3+�Tw��k�|s�94ҽ���s��hL��V��z�E1gN�;fFy޹�~u[�	Y���4�'Gc��#�pÈ#"����}��x\�_���m�ܾRroL��/�ȯc��E��^s�Ԑ�ÆE�c���G��j��jd����G�#�����]t  �{�� @����     �Ej���>����gG�������F~�5�x�uG錱c#��������rˡm���O������m��g̈|���fú��׆�Ɓư��$�Gٛ�1fLD�}����"���h�O�I�F��E�Pr�6ݴ�$m��g�h~���go|c�ӯ�l�;�l�e��UWF��C;Wn_�aâ���F�C�Nс ��)�0ܽ    ��E�	�"�t�ȿwmd[l^w����o~3�'�8T�W��2T^�ۗ��l�M#���h��g"F��P8'{��#�������|#J��c���c#�l��A��K�OK�	�y�1/�}���f�_�&�t&X�l��鑽�uuG�[Y�#��9@OJ�t  �{
� w/    �h�Vp��h~X��=?�5֨;MWiL�1�gt_Ѱ
��ox��=>ϣ��~�Ϙ�F�7�6fL4����"[����1y�PɽO(�/�>+�g�ͯ|y�o�;6��΍쵯mo�5rd4���h~��+�\w��j�_4?�ɺc�����{
�  w/    �eYw��d�|e�]���h�U�d���WD���s�<�����e�.�p�ȯ�<��7nC*�$?�;ј<y���7v�=[nنT��ܾ�����˿D���]4fL4�߿=�*��3��Zw�����A�G��e�\� ����; ,N���#     Х�d�{���=���&����ͣ����S#ƍ�;M%�M����g�F)��`�?�k�]I��(���>*�/�쟗��*:�ϯ�1h���C C�      \�V�	VL�G�������)�-��)�Mo�;
���p�=[o���V�;�_���}.�'�1fL�i  ���;      0�z������_ta4;,"��ӓ�W�2�K.��>{��r{����ht͖�l��#�~U4�ޫ�(  }E�      L�VDJu�X.٦�F~���6٤�(�o��h~���<��c�N}K��M�䞽��uG���;G~�Ց��5uGY~�VDY֝ �(�      ����7���������W�;M_il��ȯ�2�6�;
���6��{���GG��_��W�1jT}9*���g#�}��  �@�      L�Vp;6��};�XDïz�![�ȯ�2�n[w���2`%����g���WDc��r~�Z_:>ʩ�� `���      0����K-�h�ȯ�6[mUw��7fL4�uJ4�:ʍ����;l�J�٫_�lv��ƶ�D~������)�h}�(O<��$  ���8      0�zd�{c�"����^�V�QG�E�#?묈q��N=I��&�Rr1"�����Yy���L4�����c;sf�̟������NIu �v��       P�n/�gY4?�h|䠺��l��#���h}h�H��}�q�gd�o�ԩ������7��w��tn���l̓�Xu�ꆎ��gD���H?�ius�L��#͞��CV_=�SN��mom�9m�~8�-��t�-���6ҽ��	 �E)�      ����F4��}��$/[w�ȯ�<��{D��/�]/�l|[��匫�u�O>Y�ܺ��(�K/���'F6~|u�G�����������v�_1}F��go|c4O�vd�xE�ΨTJ��?�oq�o#͜��_Ez���� ,3w      ` ���;¢5�����ј8��$,�ꪑ_8-�=����ם�V[6�E�>�Q�}vu3�ͣ�F�ݣ��OD�����ܳ�lضٍ]v��c#�o�+�("����~u[��o�t��fΌ�7��d  �Pp      S7np6,�'��m��;	oaQt��#�xc�i��es�3�Dq��������ݪՊ�珍��C�<昈F���}��=�`���y4?��ht`���W�i��H��:үo���n�x�ٺ� ���; �/�,"�;     ݦ�
�#GF>ujd���7GQDz챈G�x�HO=�ԓO?�ɧ"��7T��;/�x>��s#,z[Q��iV+�q���W��GD�5T�;6bĈ�F��Xi��a�"V�ؕ#ƭ��ʑ�<.b�q��E��C����>�F�����]����CE�C�G���f��r��O=ͯ|%"���ӧ�ܳu�ڰ��s�|�ꑟzjd�lRͼ�U�n�5�O~�O��?��ӟ��D�Q� ��)���R6��;     �AQԝ�/ƌ���3#{��k�P^ye�_�b���H���驧���e6rd4v�)���T=e�#"?}j�8 ʫ�����eڱ�==�@�&N�tｕ��%�EGzxN�SO�3������=�#[w�H3g������N���� �r*�(O:)Z�uJ�ܹ��T�R Н*z=# �bY��;     ]�U֝`�ر�������G��#���CeҊ��{��(�9'�wo�'?�'ða�<�h�C=�C��6��W[n�=;Z;�`����(���"����F�L���ͬY��W���Ƅ#��Z������S��t�r;KC����� ��    ����+���߉�-o���4kV��.��~���WD���(&N���G׳�?ϣ�����Ν?�@��f՗��+�'Dz��f��t�QL���#�5*�3Ϩ�C*����m�ͣ���'V�}��ʫ��b��D���k�@��t  �{
� ��,bd�     �B�{���F~�E���M�_�~[oi��ZίDJQ�65��w���Ý?�ٌ��_��?����F�f�#�:��r��~��w����ҝC���3����GG~��}��=[��p�U"?��ht`���ł�:��h�OēO֗����{
� ��d�;     ��?�w���F>��6ڨ�g?�L�>8ZGY��B�?���[F��:x��/~!{������f������Ѫ�F��fώb��s*��~֙=_r�^��e��5F>czd�zW-�4��(��:�Ӧ֖��6,E�u� �vRp`(�    ���ϯ�܅��׼��G��o��=[Gyɥ?��<�ɓ���/FEg�βh~�?mr��e�oV}����֎"=�@e3�Q���(v�5�駫:jT�g����^����]7���������WD��W�1Ւ��Ŷ�F���2�V[M����� Yw      �O�c{y���򢋣�~�H����;�,���7�>������Yf�;}-�l|�S�VZn��s����H��_��>��#�=��X�����GG~�ٽ��}Ԩ�^��\�ͣ����1fL�s-��Gk�����OF<�l=�ͦ�; }M�����_D�y    ��t��>vl��=�������־�F�c���\�t�Ql��H�_�كnr�4���B�e���|s{<�|�/��W7s ���Y�>�����n�Q��uf��_����H0��    IDAT�ꪑ��ht`D�u&��I?�q��2�k���|�ϳ���; }M���V��    �h�,{7������6ڨsgFD�����߷�r��=�+<�x����~>�(:wn�E�K�E6~|�΄6�6߬�r{J�:��H7�X��R^uU���R��Q�"?�����j�v@��z���9�k�����`���R�_�F������@_jd�. }M���6��]w     *����fγ�V3g)d��G��wu�H)ʓO�������;�ۤ�)�t�������;w�I��G>uj����(O:9�K/�t�)O9%�+��v��ё�}V�ȑ��m��U�Z��v���#[s�'z��y��o�hw\D�UO�V�Ҙ�3 @;)������ug     �:�;���������٨.�|ꩡ���N����.������=������cQX�1c*/����/}�ҙ��uđ�ڡ�GGV��6��^�o�0bD4�?>�'�X۟�鮻����QN�^����,�^Rw h'w �Z�QxR    �'���#?�̈��⩃�NI��m[o�����}�|2��'Gk��t�&����V�g���~�a�+������kG~���u���W\�{���k�@�+��s
� ���'u     }����"?���ͲU�B`y�eQl�C�{�;J�J)ʓN�b�]"y��40p�O&b�ܺc��4kV�>l�1j���ZDD4��*��#�x�z�E��L��F<�L=Y�@Sp��5�    z[�G���G��"����Rp/�h}�3���G"�ϯ;MOH?�I۾7ҭ��;
���+��c���"�xc�1��J����9���q���0gN;M���9���e�@_Sp�����    ���V���s������'��b�ݢ<㌺������QL��7��_YF����NѿR�ַ�Uw��dY4��+"�j9>��7Q��}�n����Le�� �5w �Z��    �'e�xG���"{�;�w�3=��|Μ(vx��n�;I��ӟ��s�(����$�����{���ҏo�x�Ѻc��ˢ�~�H>XwL�Һ3 @;)��ײ,���     ,�,��>{G~�w"V_��G�9s�:����Ŏ"͚Uw����s��o�(/���$з�k�Ww��W>ϝ�jEkʔh���g��;(�L����@_�Rj�o?     ��*�D~����g#������G��.�چ\����!�Dy�u'���~���#���;7Z{��I'ם��R�Qw h'w �\ց߀     ���׿>�gD��ww���zv�{�яE�뮺c��V+ZG�;�N}%����j�P���EQw����'�m����� �B����      Ԫ1aB�^�Zku��t׬����y��ﾺ����t��u����~�È��1�΍��_֝�o��o�b��{ �Pp      �1bD4�||4O�ZĨQ�;7�(O�ڹ� X��GuG(�7��/��9?��&F<�X�Q  ��*      :.[s�h~��������R��>:�s��� �(�(��S��?�Sw���jE��<�亓  w      ���w�;����*�=xa�}��=`@�;���ү~Q�J�
�7/Z98�뮫;	 ��i�       y�����ӕ�@�я�0x�������/��Sn ���;      �v��kG~��8찈F�M�R�>��v�+��#��_����[n��}�E�󮺣  ,w      ���n��3"{�:xYF�ȏGy晝?`��_�Vw���n�u�zVy�Q�41��G� 0��       }bذ�V[-b��E��zd��w�+���ד�(�u�aQ^|I=��y�"{��)�yg�zOJQ~�����	u'  �     �zcW��Uk-�c�Q�/���կ���Ǝ��ǌ1r�߾m��Ϳ:�ٌl���G�1jTĈ�Co�G�1|DĨQ��1lXĸq+�1T�(�u�AQN�^w�����Y���Tk������u��Q^zY�I  x��;      T�1a�hLر��k��h���]Ww�����n�?�I�1`��<Ş{F��ֺ�  �W�     ��1~{����N t�4sf�&��� �ߩ�      ��SOE��.�� �����Wn �R
�      @��H;N��_ԝ �b��E1yr�ܹuG `1�       ��t�=��탑�( @�*�h���Q�uV�I  x
�      @�J��jh룏� �V��Eq�G"��ם ����      ��t�Q���y�� t�t�}��c�Hw�Uw  �R��        ˪��(>��r; �X�[��n;�v ���      ����߈�!�FE�Q �.U^~y'E<�h�Q  XFy�       �JJ����G��o՝ �V�?���ԝ ���      t�矏�!�Fy�eu' �QJQ^|I�>�����;  +@�      �n��G��G���N t�t�]���'#��guG �
�      @�z��(v����;	 �m�"�o��/9���N @E�     ���x Z��i�캣  ]&=�`�&��w��;
  k�       ����6Z��� ,�(� �)w      ���n��;F���   @�)�      ]�<��(v�1wn�Q    �A^w       �h��u�qQ�tr�I    ���;      P���������ں�    P3w      �>s�D1y�H��Vw    ���;      T$�zk�ܹu��i�3Q~�3�z��( tX�㎈矯;��j՝  ���      i}�(����E[o��  ,R��         ��_(�  ���       @ǔ�__w  ��)�       �1����  �b
�        tD�93��w�  �b
�        tD9}F�  �.��       @G���   t9w        �.�sO��w�  �r
�        �]��ں#   =@�       ��+����  @Pp       ���y&��o�;  ��        ,��##{�#[m��g���裑~��矯;K�n�%�(�  � w       �'d[l�	_�X}��y{��(��7b�#5%�Ŕ?���  @�h�        `��,�Yg�C�=""{�["�������gc��}w�	  ���       t���$�sΉ�QGE4_s��X#�K.��ĉ��J=Tw  �G(�      ��,�;A���*�����D��fKw������	�<�?"��XF/}i�	  ���      �C���\Ĉu��K��Gc���ct���u'X�Ƅ#����^��e�����;�ug�z��f������#   =B�      ��d[l�ԩJ����u��t\��C"[��c�E�G󳟍�'���y�馑_=#�׿��p+(ϣ��"��;I�eo[4��c   =@�      ��d�o��^�A.�GD�j�E~��6ؠ�$/}i��'��]ɸ��)��.�Ƅ+��B����W4��޺�Ԧ��O�s  xQ
�       =Hɽ_n_�e/���K#{�[k��m�Q�ӯ���v�ȑ�<��hw\D�W;{i��r���N4�ٺ��D��:��ԧ�  t9w      �6K��}Ă���6�,�o�����[n�駷���m7n\������э����#[k������"�pZ��Vo������_|Qdo[GϭBz��9�T:��מ�m�E�3 ����      �f��ۣ�cψg��|v��o�g�a��2ʶ�<��~+bذ�g���C�|���9?�,�6|x4���h�o5�^L��O*�'�1jTۏ���_#�>=�׿��gEDdo��#�h��f���4cFe��'��8�ڒ{�E~�W"V��  @�Pp      �t�Q�W{J�D��T�-6�|���ln��Q�W[6�/Ny��:���J�F4�9:���lV3sQƎ���3�q��;c�5׌��K���v�=g���/�8�5֨lf���hM�)҃V6�EϜ5+�	"=�puCW_}��'򼺙  @�Pp      �%���[�}�rڴh}���V����}����#V^���ek���G����^*�FE�䓢y�Q���]w���"VZ�����5iRG��>{��h�4�Ғ{��&���Q��  ���;      @���~�����k�}���ˣu�G+-�g���|����_����_�����\� Y4:0�Ό;���������W��<�������l�2ghCɽ��Gc��*�  �w      �kk�}�%��#+�����ܾP[J����E��w���w�l>n\ɪ�m�E�ӯ�l��Vl���ќzZ4;��`/H��]����Z���2{v�&�1��f6���^W�<  ��)�      Ԡ�%�ӧ*��`P��������y�F�����ãy�W�y�q�n6�J��z�_q�r���5ֈ�⋢��V��J��������t�H�fE1aBu��G����gE����  z��;      @M���o�����_�#��(��6��<�h��e����\3�K/�ƤI�ei�UV���s����tY���D~�Ց����I��3Tn��+�[�4{v�v�XY�=[c�h�qzĘ1��  z��;      @����gP���ӦE�#W��="�&�7��E���O���Xi����hst4O>)b��}x・E~х/{Y�1�=�Ȼ�ܾP�=;Z�v���H%�׽.�'}3�٬d  л�      j�����\�}����e�{Dd�~u�W^�ɓ#�lȢ����_pA��V���Nhl�}�W]��_����������y�qÆUzv�=�k7���4kV&T�ɽ�����*�  �.w      �.�֒���5P%w���UN��Ï���c�Dsʱ�_��������W�l�5"{�y���̧#��3;(�p�ȯ�2����G���"�h�h|��1���Gc��*?3�}wv��0�	i��m�U��w�5�?��Y  @o��g�       }faɽe��]�����Ї"�ϯtv7Qn_�rڴ�����G4����6�4�gT:�k�y4;,�������њ8)bΜ��U�4{v�&���i�l�o|�c�y4�3Ψ   �klp      �"m�����F~�9�GW>�(�/Yy���:���V�Q�;UoA�C�5+�	*�����h�O%�  �ޢ�      �e:Rr3���uRn_:��G�##ʲ�(� �}wv��r�B���,���C]�Y  @O��       �?J7��^{G~��#FT:;{�[#?��H7��ҹ�1"�w�6�����?�b�#�{���u)�M����W���ѽx��G����1�#[m���#�N�\ҝwE1iR�#���2i��hM�9�i�"^��
�kqxd�FE�_tc  w      �.�n�!�=�*�W\��6�$�M6�tf�I?�!�}��r�B�ZrO����<ҝw���&D�/�T�=ͼs����uG�\�5+�	�y���Xc��5:0�׾6���x��
  �L�      ���o�bϽ�Rrg��o�b��",�;J��Tɽ,��կE���-r�wy�E�fΌ�O�l��j�l�̙QL���cuGi��7�g[l���Q~�C����OD����S  @��      ���{gB�}��(�ϝ�C��k������D��6��tRd���P�e�f͊b�]��ܾP�5+���+���N4O=��d]�(��s�H��~�I  �6]��      ������>[w��6H����iӢu��܌^�4sf[m����?{��(v�=�o|3"���[�;����s�;JǤY���0!����7�y���Fd�|e�I  �6
�       =Bɽ��ܾP7�����G���#�{߲]�jE�_���D̟ߞp�!���QL����uG�4{v�&�<P��2n�Ы*  ��Rp      �!J��1�������R�'��{F̝��cʫ��b��#ݷ��6H��Ť��ܾ�M��&{�;�����  j��      �c�ܫ�������Ϗ�~�EkʔJ2�;�b�m#�tS�3�r���ٳ���D%���8��ѣ�  ��      Ѓ�ܫ�����*����b�	QN�Q��'��b�ݢ<��j�.�?�۟x��gw+%������<���c  @�)�      �(%��ܾx�.����<����t�m�9�(�5eJ�>�ю}��o~�ܾi��hM�9b�#uG�z����/�;  t��;      @Sr_>��/��6-ZG���{y�9QL�)����ˋ/*����t�mQL��ܾi֬(&L���Ō��u�  ��Rp      �qJ��F�}�\о�{QD�GE���(���/F��ϣ�f�H��u{����(v�%⩧�2���ٳ���D%w  �o(�      �%���ܾ��.���GT[r�(v�-ʳϮn�2H�C���EW;�W�E��n���@�  �{
�       }B�}ɔۗ_9mZe%�4s����n� �
X� Z��)S���n�9��#�|��p�E�  �k
�      ����_-������{+L�G�}є�W\%�t��Q���H��Wa��R�'���="��]�1?��(>���y��6`���њ�s�#����̝۷�~�n�-"�忾�d  hw      xA�##{l��K7��v�G<�TR��Sr�[���Y���"�{�P��]���?�U~��e��?���x�6$,i֬(v����WZS��\�n��wD넯.��E�)S���� @WPp     ��������?�.h��<唡2ޜ9��H�}�r{��iӆnZڒ��y��o�hM��B���-�sO�������놾����*�Y���qB���;J��SO�����V�W��E-�����G1qR�'���T  �M�      �J���E��N�?���ͼ3��w��~>�(:��͠�ܕ�ۧ����*��ٳ�x����>�C�V�OD�ݣ��7"RZ�C��ӣ��#�{�C�G�=;Z�v�M�)Ey�	�����N�~)E�C���iK~\YFy�yQ�{�H?�Yg� P���  �Nϯ��+R����    ��l�5��OGc��#ƎzcQD���(O�v��]��N��Ə���'FVw��)��h��q�5&M�族�h��~���k�u�s�֐l�5��*��)b�U��}�9�F�S��h�jH68�W�:�g��*���1�駣<�(/���(��v�hqxd���Co�7/�3�<�Hw�Uo@�.�;��K�! �]��k
�    @%ƍ�h6#�x�E7��Ǝ��GD��Z)E�5+��^婧�����������l��#,��I'Gy�	u'���lF��҈��"�����@�Rp��)����     :#[s�Hs�����5v�P�֫w P?w �Z^w        ���?����կ�}  �.Ө;            D(�          �%�          �

�           tw           ���;           ]A�          ����          @WPp          �+(�          ��          �

�           tw           ���;           ]A�          ����          @WPp          �+(�          ��          �

�           tw           ���;           ]A�          ����          @WPp          �+�u     �3'"�ϤȞiDz*E67""�4��l\iLD4�ġ    IDAT�����՘     z��;     ,�3)��"K�dwF��9,���~��'�eHZk��<_�DJ��#eo�"�[D�nSn     �Y
�     0�Y�8K�q}���ܜ�~�s+:4��'"�g/�'""��/����ٻۘ������߹�s]����8�9N0-2�e4�Ӯ(@ԭe+E�`t��:�Vt�Tc7E�Z��A��Ҕ@"5��MQ�
���5M��BӐ�!�ulb�I�:7��@�4ʍ�|����|���O�y��R���F��E���~     ̻�=  Φ�`��5�-�;   ����Ԉ_��'�:�`Ƃc�]6�O�uQ��qU�   `nܵ6�ܟ= �'�    ���G�ǣčk���=�%?<��"��`�7#ʏEĻ#b[�2     8�z�     �z"����J�k����mn���ϴ6}im���~7��F�PD�y�&     8W�     ,�'k��WW._�~�['�7�:�������{��kć#���M     p�	�    Xh5�f�쯯��\y衣�{NU9p���h��NK������=     p6	�    XH%�@-q��h�-�z0{��ڱ�y�p�.�?����     �� p    `}|u6}����x�m4��?�^5n��     g��    �Er<jy��h�����c�cΖr�𱵃����w    �|�     ,��kԫ��1{ȹ���yS�f�Q���     g��    �E�����_���r��:���d��5�粷     ���    0�J�O����9�X��,�G�X{��o��_��     �c5{      ��_\�~�Dt�C��{�׈wN6�G��?��     /��    �O%nXm�W������������-{     �w     �P�������+Z��~*jܔ�     N��    �y�;�����۟[�����?V�~6{     �
�;     ���������������y�dm2�."���     'K�    �����t��r���!�<����?G��     ���    0j�������!�f�h�P�G"�fo    �"p    �}%nX?x���3�ն��ֈ��;     ���    hݗ�\����cۿ����w     ���    в�����{��C�]������#�fo    ��"p    �]5n�on~1{Ƣ�F�E�'�w     �s�    ЪG�������_����     �l�     4��l���gX��|4����     �l�     �����Of�XT���#��     �Lw     �S�ʝwN�g,�r睓��d�     �g�    Д�P��Od�Xt����Q#f�     ���    Д^�Gʁǳw,����'zQn��     O'p    �%��R>�=bY���ƈ���     O�    ЌR�7����;�E9p�H����     ��;     ͘�zs��e��p�    h��    �V<��җ:M�[���[#©�     4A�    @+~��s�8{Ĳ��5����     w     Qk���˪�    �6�    hA�V������f��GD��     w     Z��2}#{Ĳ*�=wg�      �;     �j���ް�J�     ��    ���dOXv5��     @�    @�:���	K��{�'     ��    �l��m�����"�]�     ���    �l�<�=bٕ�G���;     Xnw     R����o�Q�     R	�    HU�ތ�C�     Xnw     R�R����T�    �\w     R��U7��     d�    �JT�     �M�    @�*poEu/     H&p     W���	|K���	     ,7�;     �j}I���ە�     ��&p     UU7���^     �J�    @�NT݌��     ��    �����Q��     ��    ��e��K�     ��     dۗ=�����     ,7�;     Ɋ��5�D�+�w     ���     d�U/�{i��ew|8F���     ,7�;     �+S��'�G�     ��    ����2{��     @�    @�R���]W�M�     @�    @���5b%{ǲ��%�5�;     @�    @.�ll\�=bYM�ë#�y�;     @�    @J)�foXV��    �&�    hB����˪�µ    �	w     Z�O���G,��ᾨ��;      B�    @CJ-��ްlJĻ�7     �S�     4�D}W�(�;�E�(����     �"p    �%{�{��!{Ĳ���F�Wd�     ���    hJW��doX���7     ��	�    hJ�����eWg�Xt�={�+"�N�     x:�;     �)�9Y�,+]�`�     x&�;     ͩ%޶���ײw,��={^[#ޒ�     �I�    @�zQ�G�G,����Q�g     �3	�    hR��}[{ޖ�c�l�(Q�?{     <�;     �*�~�^|�����^tѮ^����     ���    ��]6�����b�_�P�f�     ��"p    �i%�OO��g�w��ˮ�?��     ���    �֭F�[�`pQ��yU/���(�/E�J�     x>w     �W#��K��F��-�F�ƽ��5b��     ^��    ��Pj�y:�?{Ǽ�n�D���     p2�     ̍�?l��0{Ǽ��QK|8{     �,�;     �Wj�<�n���M��7�(��     0G|�    ��Y�Q~m���?{H���]]k�FD�go    �S!p    `����֞=��Қ�pxe��3�+{     �*�;     �jw���M6.�&{H+&��yC��BD\��     ^�;     ��Z��m�?�=$��`��W;"���     /��    �y�^j���`���!Yƃ=?Y��zDl��     �C�    �"X�(�}2�zݻ���1�J��]���zCD�d�    ��%p    `a�o��'_��󷲷�m������]��-     p��    X4{��_�������s��������D��#��{     �L�    ����(�ir��ݓ��{�ǜ)��ˮ�:tW�����     �4�;     ��U5����O�K.ٝ=�Ū/��x8����Q��=     p��f    ��9�wo|�ߚ=�9_�Z��S�Ξ�)Q���j�����ӈ���<�=�d�K.�=^]}�d2���ؑ�     �6�;   ���W���]�3���C
DD�z�x�jď���_�"�������G=��^�w��{�$�{JĶ�=     p��    X6kQ��"~x<~1j��?9qK��7�U���>���G��K�����    XB�    `Y�"�uQ��&k�o?��ů�lm�޹������m�z�\7���J�K���    @��     �3J\�ո�[[���;j���"~wu}����ř���w����ꮔ7��N"��E�F=;     �?�;     �U��=���Ԉ59����p��7j����]-ktO���D��VV����f�^��Y�;K�v��Ԉ}Qʾ����x�;�D�    ���    ��5vG�7�Q�F��FD�E��V�^zQkD/JDԨQ���v     8)��           !p          �w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	��    8sݶ-Ff�h�t:͞       ��;   �y�ߏ�G�f�hN��E�      0��          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4A�          @�           4a5{  �����j��5�ϞA��~8�����=        x�; �t�\[�+~�G�g�쫟�L��        ���            Np   X(;f�عsg���w�D� 8�f���_|q���>~<^����3    ���   ��'���_~y���x { �SO����G?�=�d����kn�9{    ��^�            ��          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          ��;           M�          Є��   0��O����f�����3�3;~<��'�����      �  �I��J/�����++�S��}��7ޘ��M;vd/���6��O&񊚽     �=��   0��5�N�o�Ǳ�*8u��͢7ފ?�]�     �f	�  ��Q��6ފ}3q" 'g="�O&񿧓����      ���   N�����l�'��g��i�w]�lk+n�f��(     �&p  �aZk���bc<�a'Y��E�U�i��d�S�     N��   N�}����8��N�d��	�t]�bk�Ϧ1�     0g�   p�ND��i�O�e�)� ���i����v     �c5{    ,�?���p�����VV�� p]Pk&���*l `�}�g�k/ّ=�D��7�s�/g�   ��   Π#Q��t�9����~/%{ g�k�.�N�.o�  `I���s׮�$z�ǲ'   ��=    ���m��7s�/���WM&��8�     �w   8KF�Wf��?�x���������㸽���     ����:   �E�Z�:�}�����<k0�Vj�+���_�,��c      �_�  ���v1����4J� ^�Kk��'�M�     p�8� X:+ǎ�;�g� �ۻ.���=X2'"���4����H5��;���r:���Y�5{
     �B� ˧�8t�p�
�m��q���3�%��unM���c*rh�t:�?��      KA�   	��G�����z� ^�K�͞      �4�      �L��я},{ɮ8�-�    ��;     ��)�Y�z�oe� ���wD�~�    8%��           !p          �w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           � p          �	w           ���=        ���ɽ��c{���ײ'   L�       ������h�e� ������.|Y�  `A��           @��          �F�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&�          h��          �&����w7=v�w���}��x2v\�Nl�q��*8}�(bK� � �-kĂv���G���] �HTm�� TK	I�3��9s����*iK�p�\���?�7��"���|��          A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A���6    IDAT          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           � p          `�           ¼�  ��V�����?�z�=�����3        �� p &�?>���?m=�ƾ��/E��[�         ~B�z            D�          �y�      lV�|��w�z�}�o���z    </�     dSJ�@	�    0>^p  �3�E�+�Ǳ<؏\.���/t4�ū{{��Λ!      �$p  �3pi��������i�9 <��}ߺ?�=x�������ͽ�X�     ���   ��\��������A|�k� �wRk���q��q\������n=}1~�X��     ���   6��2vޏ;<�7��� ����:�88�88�W��慽���^ͺ��      FM�   p��㥃��{�ժ� ��7W'���9�������������]_�      xw   xL]D|��(N�⟏��U�0eǵ�W��"����lw�z*޽x!�Y,ZO     �;   <����x�� �������u�9 н�:���G�����ĥ���ޅ�X��z     ��	�  �!�j���?�?�Y.�[� <�>"�u��X.����Wvw��ⅈ��5     ��-
   <�?Z�q2?�ܥ�S~lu�||��?�zF3���/D���3 �/��m=��,�����ϛ���qS
     �g�  �C�+%�Ji=��Xv]�vvZ�h�ٮ���Hf��3�?W�Z�Ο$      C�7           ��          �A�          0w           A�          � �          �;           � p          `�           ��          �A�          0w           A�          � �          �;           �0o=    x<��899i=Hd�Z��l�zƙ��U�	  0J����Fw~������7���   )�;   ���|�~���3��.��o=R��{�b=������ `�~�7#.\��z}�_�  [ӵ            w           B�          � �          �y�  gmo���~�g�����n�	        �����[��w��K�g         �]�           �w     �t��u�׷��z������    ��	�     ��[��w��OZ�     xd]�           !p          ` �           ��          �A�          0w           A�          � �          �;           � p          `�           ¼�    ����>._��zF3��� �+�<�٬��3�X�[O      ��   0R��:�^��zF3wؼ�}6����g������      ����            ��          0w           A�          � �          �;           � p          `�           ��          �A��[�e�	        t�z  l����j)Zo        ؔZC@jw r�ա       H�x���� �VJ}��       ���� ��[ �m��<��z     @���ƺ���AC7��� &��; �	�ȭ��p     ؘ����� ����; �u� �6��9�       ix���� ��uu       @� ;�; ��u�^�        �2�� �	�H���u       @����7 �6	�Hmg��       i�R�[o �m��[���        �)}���  �$p �w��       i�#�Zo �m��Z�XG�I�        ���l�? R�0n.       9��: R��^�ps       �`]�|s�z lӼ�  ضR�(j�  �7[�������fJ��<شW���X��i=���O�   ���z; �� `�N�_�Z�x��       �'���{?��z lS�z  ���      �[ �m�0w       @� =�; ��Z�       ��G� HO�@z]q�       2�� �	�H��       @�� L���)�       ��E=n� �M�@~����        ��J�ZO �m��_�       �Wkh  HO�@~���       ���� �; �U/�       x��	��_�;       ����� �W��       d��  ?�; �u�:�       	x���� �W��       0~�b��ȯ��       �_�@ 0w ҫ���       @^p`� �Wz��      ��+w ���_��       ���J�@ �������       dP���� �W}�       H�� L����j�n/       �W����ȯvw       @��HO�         cPJm= �M�@~]-�'        <���  ?�; S�p       d��  =�; ����       ����� L��       �@��  =�; S�p       d��  =�; ��2       �@��������w       @U�@z�? �+w       @�����v ���<       ����� L��       0~�W��O�@~��y       d p =� S�p       d��  =�; S�p       $�i  HO��8�       )h  HO�@~��;        �Z� �'�`�       �4 �'p ���       H@����;         �	�ȯV�;       `�j����v �W�E�	        O��n�z l����J�ϵ�        ��4 �'p �R�       ��+Q|���� ��W�;        ��? ���_�w       `����������       �Jh  HO�@z%z�;       `�J��= �	����       @�� �'p �"p       Ư���� �W��       0z}�E� �mw ��y.        � ���^���z       ��+�[/ �m��^��T�        O��m�  �M��8�       h  HO���;        ��W�HO���      �ѫ�k  HO��T��      ��+�b����;        ������	p{       HaQ#�G �6	���*p       r�|Y@jw R�ѭ�E�        1�	�HM�@nn-       ���T� �Mw rsk       H�������Ԏ#�Zo        ؔRw R��Z�X\l�       `SJ�k! HM�@j]�P       䱮U@jw r��C       �F�B ������έe        ���  9�; ���       �B �����jy��       �M��HM�@j��:        �R� �&p ����       $��  9�; ��Z�       �D� �&p ��P       �QKh! HM�@j%|�       ȣT�; �	�H��C       ��ӭ �6	���R�        �\� �Mw �s�       2�B ������       �L.�;wε �"p �1���w        lԻ�>�z l�����]{6"J�        ����|���� ���:�9        ��M i	�H��p�       �)kM y	�H���V       ��K��  -�; i�e�0       �S|���� �U��      �|4 d&p �һ�       �S�&��� �ջ�       ���  /�; i�p[       ȧD\j� �E�@Z%��        6�F}�� ��; i��9        #��������       @F� ������       @F��;wε � p �z��ND\l�       `J|�� ��; )�       ���z��  %�; )�k��z       ��t}��  %�; )�:sK       H���F �������q       @Z%:m )	�H�tw        �Z� �$p ��3\       @bE@Rw R*�\i�       `[J'p '�; )��˭7        lK���? R��R-�Z�        [�B� �w R*5^l�       `���  � p ��U��      ��v�[϶ �&p ��o]��y�        �tr||�� �4�; �'o       @z]�i$ HG�@:])/��        �m��; ��H���       ��J�H ����tJ��       ��j��r@:w ҩ�8�       �y���� �SJ8�       �U� 		�H����       �$h$ HG�@:5��       0�jDi= 6I�@*5bV"���       p�ŵkj= 6I�@*�/�t5"f�w        �����{ R��ʢ�o��        pVf�j% HE�@*�֗[o        8+�V�d� ��Ew��       ��R������Tj��       LG�z�� �$�; ��w       `J� �"p �R��       LG�����d��n       �Q"^��n�o� 6E�@�ƍKq��       �3T���7Z� �M��ƪ�}r       ��Y��	 ���F�pX       &��z�� ��; i��	�      �ɩ��  �; ���       0=E3@"w �(]8�       S��  �; i�Z�       �	*� ����H���        �^�Y��9�z l����/<϶�       ��ly����# `� �p:��n�       ��y)�	 R��B��!       ��^;@w R�n!       ��k' HA�@
�!       �0������C       0]��v�� �P�       �I�p�{w�z <)�; �W�_�PD\j�       ����^n= �����[���v       `�f��P 0zw F�:�       D-�����0z��       @D)
 FO���U�3       ��54 �����s8       ��� �I	���c�        �+����# �I���7�G�s�w        ��d�w FM���-���[o        ����q�0j��;�7        F-w FM���u�j�	        C�E�0jw ƭ��       ~�
�9�; c�w       �+�w�.Z� ��%p`���/��Z�        ��ɽ{�[� ��%p`�NOO}R       ��4 ����Ѫ��i�       `h��
�-�; �U뫭'        M�!p`�� �Wq�       �g�T 0Zw F�8�       ���Ոy� �8� �R�r�jD\n�       `�v�ׯ��z <�; �t�X��z       �P��|�� xw Ʃ��[O        ���� �q���       ���x  �$p`�:�0       ����x  #UZ �GUo��]�������       0T������j� ���U��C�       ��:��?�z <*�; 㳮���        0|�����0F�j=        `�jT� �#p`|J�]       ��i, �; �R#f���;        F�#���/� �B�������G#��;        F�;],>�z <
�; �Rf>�       �j���Q�06�j=        `D� ����Q)Q�*       xh���Q�06�l=        `<�k���E� �� ���՛�D��w        ����޽O� K��h�Y�k�7        �N)� FC��h��?�z       �蔢� `4� �Gu�       ����\ 0��  x�����у��i�       `d�"�r��;�� �/�w F����n��       GYwݯ� C��8��SY        �i��gZo ��!p`j�_���M����S�U=3		Yg��2B��-A�M�[T""�\Xr����Gp?p	�x����9G�	��Qnsk0�$�]=�$��LWU����$$=���Z�?��yU]S]5��~��d       �0���d       ��Q�f�)�� ��}�RD���        �b'��9?; ; o0X���       �iW�Ge7 �=1p`���
       �x�b���3p`�_��        0�J�` 0���h5�Q.��        �_]O=��� �J��h�N�qbv       �h�v�|Dv |%� L�Rʥ�        �b\�%� ��0�j�R       �IJ�/�n ������U#5���       ��QU{��� pw��X�N�qjv       �Y�zQv �w &W)�f'        ̚q-�d7 ��1p`b_�        6])��� �;� L�ѨQ/��        �95.����� �+� pW���i�0CF�o5�q]�r]-�O4">Sk��;�K�L���h�P�'����qm�\�xwD�_������.�      �f���GE���C �K�0����(5��ٝ5�W��|_�ԓ>Z��v�?��z;G���Z�eQ㢈X܌�      �����0p`��  �+�N�j�gdw���%J����?����r�5��x���/��xvD\QOڎ�      �8�x{u�� �R� L�Q���-qzvL���(����=o߮Q�ݩ���X�Ќ����he�       p���ڭSʍ7��/d���Y��R���;`��Q��j�~��t�jv�]9��tv���(/����=       |�2.��. � �P#;  �Tǥ�0�>Y�����<���_5��������7����Z�}5ʫ#���&       �@c|Iv |)w &N)՗'�r��5���~���W��o�5;��*�ݲ�_~Uk}t^D�)"jr       Q�\��  _�d ���a�{KD�����|����Y<t���K6ðӹ�F��xpv      �������'>�� �<'�0QF��Ea��w[�x^��|ɬ��#"Z��_��+��?k�=       s���j]� _����2����0�5�f�핕7���]��JĨ��6�>:"���      �W�(�g7 �2p`���KD�_o�r�w8��씭�����5X� "ޖ�      0�F�d)� �y��3wZ�p��H��hkQ1    IDAT�W�� ;$à�{yD}]D4�[       ��8��;���;  �	2l��~71�n+u��y�GD���o�Q�����-       �Q�g7 ��09j�e��T����VW?�ݒm��{i�'G���-       󢖱� �d @DD�h;݃qzvl����������C&ɠӹ ��YxO  ��D��KĿ�Zo�w֨�n���(u�h�c|J�Ɖ�����~q^D�ʎ   `�i5�iey�Hv �0�ޣb\?��۩F=X�͋w8���I����?���[  `��Q#>؈���h\;*��n,��A5�]ZڻP�y5,�~}�qI��   �/��oX8���� 0p`";��Q^�����(qi{e��C&�p�wy-����n �-T#�J�?��x_ke��J�h�1�v��Z./Qͭz<    �E}C�߿*� ���N�����&��)�~�=�!�`�ӹ�D����n �Mv�F}Km4~k���fEԳ�^ֿ9J���� �   �tk�W� � ����i���iq̋�k���9;c��uz�*Q<�  6A-Q�u�u��Q>{z��t��WE�s�    ��x�y��n�!����L �jyR�3?�hܾq���OD�{�;  �8�k�G�G����h��~h���핕h�W^��܈���8��   ��i4G�g7 ��; �J�O�n��Q�mE}iv�4*�ְ�܈8��  ��m�f����S����g��;������U�a뜈��X�n   `��(O�n �� �|��a�ۏ�3�[`����#�|mv�4v:��Q�,\�	 �t��D}i�ߟ����.�h�r�xdv    [�p+���?���2 �hO��0ng��Ÿ��}n���  p��?�ڵ�0n��h��^�Z]�ڨ�]qkv    [fנ6���|3p Um���� [�^��g��+fEk��+k�jv  ܍�j�\�ZY��r��k�1��D�۫+�6*����    �Fi�gf7 0��HS#JDyzvl�Z���k�f�̊r���?��  _��ﴆ�G,./4;e+�ZYYn�W.�Q^��    6Y������� �/w �{������;`��vky�����������  ��#Q�핕o/���g�c�C�-��_���Dħ�{    �T'�>u�c�# �_� ���[Z1���Ɏ�E%�F#^��  q[��'�WVޔ�a���j_�[    �<����� ��2p M�����bo<���~vĬj//�MD�'� ��U����VW���B����<l6.���f�    �Y��k�Bv ����k�ރ#�����Ǎ��YW�姳  �S%n���׵WV�!;e�p�@��м4"�2�   �Mq��׻8;��d�@�q�������X^�>;cֵ. "�"� ��R"��k��g�/Vn����`����    �_���� �|2p E�����Ju�xmvüG}Mv  s��Q��߿9;d�O~����"�_�[    8>%�3jD�� `������}��xhvl��w���SvżX���U���  `..%���߿.;d��C�nE}\D�n   ��Ոް�{dv ����m��l^�� [��;��D�J)o��  `歗�xfke寳C���~�@�xjDܙ�   ����xfv ����mW����,�F��ˎ�;���N  `��(?�Z=�g�Ӥ����e�    ��M� �w ���^���R"�Un��PvǼi��^Q���  `f]��/�dv�4j��o�o��    �X����zɮ `����>{몒�[�F}Gvü��x� �
�Z��甈��i���'"�9�   �c4�Wd' 0_��f����J������U#�}�  ̞F��\n�i5�c��C��WF�(�   ��+� l+w ��ѳκD\��[���n�!;b^-�ZG�;  ����ZXY���Y�^Y�Ǩ��    �s��#�# �� l��x��Q�;`��f̳r�G�Ƈ�;  ��G��Ȏ�%��ڏ����    �A�Nq`���mju�*f\���N�w�ԫ�  �%�v<xcv�,)����ߟ�   ���Z�]#�� �w �Šӹ "��[��ov¼G|4� ���KK��1���ߋ���    `cJ�=�N�� �w �I����b�U�ǲ#��x�5  `ԟ-�\3̮�U%�'�    ظ��� 惁; [�F4Kĳ�;`�(����y�>��#b�� �T��u�)��1�Z��{#���    lTyV��vfW 0���r���jD7���u�D�k�D�M�  L����}�d���Lv    UO��� �>w �\-�y���5;�Ϫ%>��  �Ժ��h�Vv�<X���8">��   �Ɣ���n `�����9�O�V#�=���*�~*� ���;ey�Hv�<(5��fv    ��#���� f��; [j��veD��ֈzGv�W>�]  ��*�;�	�U�["b��   ��4Jynv �����U���	�j)��n�j  �q%������󤬬�{�xwv    Sk<�F�� f��; [�h�{^D<*��CUO�Fq�>  W"ޔ�0��N�   �F_5�t���2p`˔Z�svl�2v���p�  �bX��g7̣�Νwfw    �15/�n `v��%��������mJig'�Y���  �:����dG̣r��k5�_fw    �Q��u߾�fW 0����[o}FD���ۥ�z��>k\�� ��z_v�<kD\��    ����WfG 0���%ʋ�`[UO���  R��u��p�   �T��]�	 �&w 6�ѳκD\��۩4���>��I�	  L���>�1�Z���D�m�    l�C��#�# �=� l��^�3"Jvl�q-F��T'� �%��:tKv�<+�qMv    �`/�N `���������y���JԽ�|Vm���  L�q]v��     �E}v=�T�����T�[o}VD���	����8/; ��Q�'C-^   ��t�pǎoώ `����J��g7@���V����D���  L��	�B   �iV^��� l&�T �4�N炈�(���:��t�#�ݨ9r�>  bX=F��   `z}ը�y|v ����M��v�[+���z~v  �e\�jv;�s�~v    �n�e� �w 6Eݳ猈����4�ƣ��  ��hܑ�@D�����dw    plJ�7�v��� `6��)F��#bGvd*1�,�aޕ��n  `��<|��}r|&;    �cV���� f��; ǭF,��K
D��j��+�b^�vϫ��  �J�O}����ç�    8%^Xw�>!;��g��qt:�gew�h�".Ύ�W�pz;  v�D�gG���   0��;l6_���3pตh|vL�q4���0�J�� ����|�qv     ǩ���� ���; �e��>6�^�����J_ַ_=眓k�'gw  0uvU�G:A�I�    ����gfg 0�����2�xEvL��u��fw̛���D���  �N#�8cWv�W�]    ��+?�� �t3p���u:��gw���5���0wJ�� plv�2��^   �YP�k�KK_����2p���(?%�&���3N̎�G������  `:��FF����ߎ���    6Ii~v ����cr�Ygu"����P'[�oώ��F��b  �Qs<ޝ�@đ�n;3�   ��S�>u��9?���d��1i�Ư'��WP��ϝ@����i���  �W-��"Z�n    `S5J�ʎ `:��a��=-J�(�&�Y��n���Y7�����  `z�hVO�Z��   `�<�����ˎ `���a���;`������ΘU��SO*%^�� �tk�a���:    ̞V����� Lw 6���w�R�%�0%�,��̎�U���/"�� �t����F���    �(�ý^7;��b�����×E���05J}M=��f6���{�)Q]� �f8�g�\5��(dw    �%j��� ���; �Zݽ��Z���0MJ����џ��5���E���  fBs��ѯώ�g�^�#���    �H��ݻ�� ���; �ڨ�zYD���ӧ�d��<<�bV�u:O/O��  `v4j�,�a��qx�   fۮA��w �5w �z�9'�p�(8Fͨ�W���C�]=眓K�_��  `Ɣxlv�<+��   �u%��Գ�^�� `:�p���7"N�U⑃�C?��1�FG�~3"���  `�<�v:�X��F4k�K�;    �r����WfG 0��Gu��SJԫ�;`ڕ�?p���O��j�鼤��"� ������y4Z�=!"��   �v�/>�{���+ �|� ܣ�h�C�ͰJ#��,-9�|��z��D��fw  0�J<7;a�2��   ̏v����� &_� `��3��=\h}<"N�n���V�Ǖ~�pv�4��w�9l.�UD�?� ��VǍrގ���C�E=���ۋ#bWv    �f8n��8 �'��^���.D����2����g�l�i� ��JǷeG̓���¸   `޴��# �l� ܭ����Q�+�fQ�xʰ����:w������ �^�� �|(Q��B�mT��    �P�t:dW 0���[����DD;�f����͎�D5�9���7G��[  �+�K�ggG̃a�sqD���    R4"�k�# �\� ܥA��Ȉ����u%�:�_�>���z�N�-�-�-  ̟R�+}>�z��n     ��F{zOΎ `2�C wm\6"Jv̇��Q��?��.f�d�g�q���?
�  �灃��ӳ#f٠�yx����    r���k�Bv ����/s���O����'��3�����qƉ�-Y���[�E��[  �o���.��2%?�_    "8�t����1p��Ԉ�F����yT�>q�j������[�۰�y̰5���xXv  D��N���h��<�F}Zv    ��D���{�	� Lw �Ȱ������q-L��Ҹf��{Qv�v�e�Ի�F�:"��� �����v:�gW̒��F���    &G���?���dqX �Cݳ�a�y]D���DD�[룗�C����
uϞ3�ƛK�˳[  �.������wfg̊�R����Ogw    0q��כ�w���� &����F�ø&��ͅk�:��e�l��,�^4l4�ٸ ��V�;��E���Ȟ=�j���    `"�h6�?���p�; 1�t.�(.~�I���/���_�r<��â�/Eģ�[  �^�xk���n��V5ba��?"��   ��*�<������ �15�D��~/�${\#�Gֺݟ�����1udi���R�W��߅q;  ���ãk��1���O�q;    �����zᅭ� �9��t�ϋo�� �;#�o�Jy���옯����4���"�wF�bv  ���^]1tߠўޓǍ���z    �R��[++���  ��;���{��2��sD��n6l-j�)���n//�Mv��Ոƨ۽��xqD\��&  �G#�c����g�L�#���f�k"b��B   @�;F%4釽����ܠ�������q��Fy[]o�yǡ�o�X�tΏh<���ܨqNF  l�O�K\�ce�c�!��v��k|("��   �t)Q����?3��<� sl���u�4>~�,G����k����F�/���x�z�'���qI���F��Eă��q  `�\�/.��r(;dR�ݻO6�e�    0�j�g,��o��  �A#���������������`K�E��8��(וf|l�ټ��t���5�]ZڻP�y5⼈���k"��ܺt  �Xi=ri�ԧ>�2i����o/%�!�   ��U"�k*����- l?w�95�v����� K�tD�DD�-j����L��L�h�K�Xj91��%N�{"bWv1  L��l-4�Zn����IQ�=wqt������n   `�7�����+ �~� s�h��U�q�hD��n  ��U��Q�/����.�V�8��Ak���O�n   `f�K��[++���jd ��jD�Q�o�q;   ����(:��< �$S=����V����    l�F��7�}6. s��`��z/��dw   ��8��/���c�C2�݇[�����g�    0����eW ��Jv  �����4�����[   `���5�~�GJ�zv�vt��5~%"ve�    0�F�(�i//�Mv ���`NԈư�{D���   �Y5�?\h<���)[��~�}���Q��n   `n�K��zx��ƣ�! l�Fv  �c��~�q;   l�����Y[�=���#å��4l/~ĸ   �mv�`0zuv �c�����[�t�/Q>;�[   `�\]��%�����r�w���8^_K\��   ��Z��WV>���2p�qu�������:".�n  �94�Q_�ޱ�g�7ܞ�Q���9�_Z����81�   ��w}k�vA��'��`��̸�N�%�+�;   `��Q��j�~��t�jv�=��w�0l������5���    _�����gG �u�fذ�yB���hd�    qg���Q�����Ȏ�R��9}T�w�WE�i�=    pWj�o]��ߚ���0p�Q��9}�%b)�   �2����ͭ�ѷf�R��{�����OlFyn�xZD��Z    �^�}}}���[v ���`Ո2�t�Y"���   ܣ;���Z��=l_]>q���~��w�)���R��Q�"�ԭ~L    �d��\R"F�! l.w�4��^Qߐ�   �zmD���������KK/�\3<��\;�}���k���؈���hn^3    l�Z�WW~,���e�0c�ޣb\?n'   �b�V#�+%�/���|����Qo��-�,�q�o4�%��Z��R�~���#���	    �M�Ƹ<e���C �<� 3��z�����ؗ�        �����х;��� 6G#; ��Q#���-a�       ��8��\������`s�̈�R��%ʓ�;        `�=l�^_���(� �Q�����.       0������+ 8>� S�h�{^�Ƈ#��        Ht$j��۫�.;�c�_�)VO=��F-��        ����;w��� ���;������ηF�e�        �$(K5�Q;�]�- w�)5�t^_J|Cv        L�F��v�(�! l��;�t:/�(/��        �ITK\1�v4���su��v���5���        �`��x�����g� p��L��^��e\?��n       �)0(Q����7;�{��`J�v{�]#z�-        0=ʧ��K�++��]�=kd p�j�{�B���       �FՓJ�?9��tvv	 ���`��^o��;"���        �F5��,�w�^��� �2w�	V/��5�ߋ��d�        ��{�p\�Y;�]�! �=w�	U#����7Ո�f�        ��x�0�;�};�C �k� �F�a��+�[�[        `�<~0���{�bv _��`�|v�������        �E%�G����^xa+��/f�0a�������        �YV�>}�?�������f�0Aֺݟ)Q �        �A-qŰ���jO	01�!L��N�ե�gw      5���    IDAT  ��y���3r�%; ��a����        0��o������]0�\m�l��~�q;        d+�1�t~!�`��$,������         ""�����+ �Y� �W��ދ��_��        0i~��_yEv�<r�;@�A���(�Wø        &���uz�ʎ �G�� �l��>?j�V��        &Z)�c������ �'� �h����R�-��n        �Y�������fw �w�m���^Qj�5"�[        �{�D��V�����y`��֖z�,��^�       �4����~��e� �:w�-���<�D���he�         ǬF���WV~%;`��l��R��Z��#b1�        8n5j|w{u�ײC f��;�v:O�Q�;�[        �M3��o���Nv�,2p��N��5�;#bgv        ���k-�[\]����Yc��Ɇ���5ʻ"���        `ˬר߶��-;`��l�a�����q��        `�k�oZ��ߑ0+�6ɠ۽(j���zRv        �m�W����(;`�l�A������qJv        ����\XY����ig�p���C���"���         ͑R⩭��?��f�� �i���=$j�7��       `��5�9�v/��fNp8FG;�����({�[        ��q���7�. ;`�����y���K�Rv        0q�,u����ꇲC ���;����m��jD'�        �X�Ǹ����0M�6�������xD�KN        &�mQOh�����ia�p/�t�Z��"���[        ��qkD}|������i�� �����B����       �:%��{m����! �����3�ܽP�=q��        `*�Q��[۳�A�! ��d L��{���f���%        p�ը�.����0���p7�=g�ܸ        �$�Q�st��s�C &��;�]����w�h�;j|uv        0;jD��\�������n�D%; `��}��;�Q��        ̬��������7e� L'�|�z�9'׆f�        l�����;�:��0I�>���}�������#�[        ���U�����쳗�C &E� ����5,�O��%�-        ����ְuY�č�C ��s�v:��Q�8".�n        ��G[%[VV�=; S#;  S��v��3��       �\�xo��N��d�̭�{0��#"��        ��{�޽�d� d1p�Rݿ�=����Y"�1�        �<|8Z��z�����`�̝zᅭѭ��~�xjv        �]��a{����3N��n��\�����7רO�n        �
=l��Uw�>!;`;�s�F4���oGĳ�[         �ͅ��^ogv�v1p�B�h��7F��d�         l���x{ݷoGv�v0pf^�(å�/G��f�         lT����`����s�[ ���;0�jDv��%�3�        �X�(��~k���Vv�V2pf�g��_����n        8^5�3F��F,d� lw`f:����/��         �,�ƳF��[�܁Ye�̤�n�gJ���         �l5⛆��oV;P`ycf��R�'K���         �B�3rf�75��ٻ�7K�����9u���@�]]�}z�iDi��vB6��B��QDVA�eT��`��$�lt��F�y���ˌ^s]>@�:�,��5��:w��̓ ��KU���z���9����-��r����⍥;         6���`�H�C ֊06��~u���         +��t���� k����~e�xg�        �"R�{zaᕥ3 NV�t ����u_n�        L���W�;Jg �,w`����OG��*�        0^�\u�t��H� NT��^�./�         |[J�+����.�p"܁�ԯ�K#�G¸        �{���Y\xK���e����~F�qyD�K�         ��u����Jw w`�,��%)�1U�        `�����^�=�C ���;02����?��         �*G�N�z�+p,܁����{Ѡ������-         #&G���^\�`��{b��fn�s|6��        N� r\:����! w��jMU]�#]�J�         ��՜��f���t�]1p�V37�؜Z�Gĩ�[         ��j���^��C ;0���zt�tCD�V�        `̬�ϜYX�T�����:M]?2��|D�^�        `L�����׻�t�w3p�J��9}>"߫t        ���R\<��pm���`��~U=,"�g�n        �˭Az�����K� D�C�_��7G���n        �0GR��t�h� X�v9n
�v        �N�9�i�u_:�w���Uu�q(E�V�        `�ݖ�����_�&��;P��n�~i���"�J�         ߌV�pz~��J� ���(�h���=ȇrD]�        �;�5r���/�u�`��n��v�#}!"v�n        �N��ϛ����t0YZ���r�����u(��        ������,L܁s���S9E�}K�         pL���O�9|��J� ��w`C�[g�r��v        �Q�5�����J� ���Xwyvvk35} "~�t         �m��ƣ�;v�Ɵ�;���m[����#�J�         pbrD��^=�4;{��-�x3p�M޵댦վ!r<�t         'mG�=upi۶]�C��e����{���~�ƈxx�         ���v�}�m۷W�C��d����{�������J�         ���tV�Νs�C��J �%�Ξڴ;�G�ǖn        `]��N�9'}틇K� ���X3��Nir�6R�S�        ���禅�+��V� `<�:��t�q;        �Dyp����U:��I�{���S�LD<�t         �� ߔw�8�t0�܁�����Y�L�qQ�         �yX��z]>���K� ���8ay���[n�t�xJ�         �{D3=sC޲��!��2pNH�h7�����c�[         �j:���'��8n9��TݏE�3J�         0t�t�������!��1p������O"�O�n        `h���Uy׮M�C��b���j���"ҳJ�         0�R�����yϞ��-��0p�I�H�\�����-         ���I+G�\����nF��;p�rDj��=��ť[         -9�SW�"GL�n���;p�n�w?"^R�        �єs<m��/7r;p��U������         ������?��W���ܥ�~s��K�;         �3rp�����J9^_�        ������~(G��!��1p�GSU��R��t         �*�����+]o� w����s�w��         `�x����+Kg ������\��H��         L��^\xu�`8�J á_u_f�        ��K����3����;�����C�         @!)ův~�tP�1+L�~U� "]��         ��o�,.��tP��;L�~]?/r�a�        0$R��uz�o+��a�j����r\��-         ��R��tz�w�� 6��;L�庾$�""�J�         �����ӽ��J� ��&��\��)�OFD�t         ܍)^2�����!��1p�	���{Ѡ������-         pr�������J� ��&D3���9���M�[         �8��.�Y��x�`���h����0n        `4���ϙ���(�/ws���csj]��n        ����#?k���d�`���k���9�qZ�         X� �%�z��K� ����TS׏�9>��n        �5�o�x����5�C��g�c�_U�H7Eę�[         `,�Z�����J� k���L��9n���J�         �:ZJ)��YX8X:X;�������C"�Ma�        ��ۜs\�t��֎�0&����A>g�n        �t[ʃ�:��Q:8y�0�V��Sġi[�         (���JN���U����È;��ޯ=ȇrDU�         
�f���Ӌ_���!��3p�v����q{]�         ������^�oK� '�U: 81KU��5�7�        ����nX�����!��1p�t����S:�J�         ��ْڃ���m{@�������9R�ݩ�"⾥[         `�}%��f��tp�\p���n��ʱ?��        ��̶Rk����m�`��Èȳ�[����#�K�         �(���������}J� �&� �Y޶mK�n�,�         #�K����o>|���C���;��k�Mk�z�v         8a;ڭ���m�^�;��{��������n        ����:8�w�+�5wR�����,-�?\�         ���7����e׶�!��K���ggOm���"��J�         ���N��R����!��Ð�UuJ�ӵ���-         0����J���o���U: ����nn"}θ         ��C�A�)��qf��;�aH�{����3qn�         �kVV��g�}z��v�0�޽��[n����GJ�         ��yD3=s��;w(,���Y���O����n        �	��fz溼e�i�C`��CA9��,�X����-         0��t�������!0�ܡ��n���"⿕n         ""��� �ʻvm*���
���8"�T�         �;R�����yϞ��-0��a���T��#ǳK�          �+Ez�ʑ�����uJ���1p��#R3W�/"��t         p�r�X9|�9b�tLw� �_n��)~�t         p�r��W��r#w�8�A�U�m��         ���Oo��d�[�~h����)�kJw          ' �s���6����~S��K�;         ��riSu?�#R�g���7S�_.�         ���¦�>h�����ISU��"~�t         ��ҋ��~g�
W��u����r��-�         ���^\xu�7.����կ0n        �1��U�U�wJg��1p�5ԯ�/��*�         ���5M]�J�'�t ��~U�0"]~W         0QR�7t�\�Ɓ!.��~U=?"}8�W         �H)��;�����Qg�'�_�ϋ��         0�R��vz����Qf�'a����r\S�[         ��rD~�t����!0���-�u��R�D�         ߑ#�K�>P:F��;����SSʟ��N�         `�����Ӌ��Qc�ǩ��>)�|UD̔n         ��j��ҙ�����Qb�ǡ��s��FĦ�-         ��[͑�3��]Q:F��;����ϑ>��         ��[͑�5��}�t�w8MU=&G�!"N-�         ��f��M��եC`���=h������V�         Y�V��M-,\S:���;܍���s|>"N/�         ��~���:5?]�V�p�U���tSD�Y�         K)�S:J��02p�;ѯ�F��#��-         ��9�Z�ɝ��C�C`شJ��Y�v9n
�v         `}����fn��J���q���rU�@�t("fK�          �.�{������*]��w���Uu��t ��        ������?���J���0p��8��ޯ�@��+�         L�{G�؟��W:�A* �-���l��"bg�         `b}-��Ν�ʗ�w�(�����TU;ڑ��J�          �y����Ç��t��* ������q;         0��V�������RܙHG��z*��ȱ�t         �w�m����۷߷t�`���ɳ�[��ƈ��         �N��V�fg�S�6Z* )o۶�i�F���[          ���V���|��K��F1pgb�:��t "T�         ���J+�s���B������]g4Ѻ!��        �Ѳgj��;�J��F0pg��ݻ��4�����t         �	�_Ӭ�[vm+�-�����:�^ͦ��#⿖n         8I�؉|n���^:֋�;c+�Ξڴ��E�Ǖn         X#�Iq^ZX���!��K��Nir�6R�S�         `���N+����Q:�Z�t ����nn"}θ         Sk��|�Y�*k����������DĹ�[          ��#�M���g�}z�XK�t ���w�t��[�,E<�t         ������������!�\pg,�}�:+���i�v         `�<��L_���ͥC`-�3�rD�Y<���c�[          
8����]�6���e��H��>?Y�         �����UyϞ��!p2�Y9����G�g�n         (-Ezbi�J#wF��;#)G����9�]�         `X��,-]�#�J���0pg������?S�         `�����W�3�R� 89"5U���xI�         �!��No�)b�t+�)����0n         8�h����f�����X����ȯ)�         0B.m��eF�
_TF�r]�)Ez]�         �ѓ_�T�rD*]������\տ�r�r�         �ѕ^����JW�=�C�����H�S�         `,�x���«Jg�]q���������         �P�W.Wݷ�΀�b��P��կ�9~�t         ��I����_-�w&����_u!"�^�~         ���⍝��7���f@�P�W�#�e�	         ��R��wz�o-������ѯ��G�GD�t         ��H�_����^�"���~n���0n         �h9"��t����!`�Nq�u�����*�         0�r�x����J�0��)jy�����'¸         ��9������J�0��)f��~"E�TDtJ�          ����f�?^:��d�N�\�I9�"b�t          w��#=w�7y�&��;���s��FĦ�-          ܩ���3��'J�0Y��PMU��#}.��         �]3�|ɦ^���!Lw6LSU�ɑ����J�          pL����t�����Tգr�χq;         ���Z�S��וa�����u��ȱ?"N/�         �	YJ)��YX8P:��f���    IDAT�κ�W��"��qf�          Nʑ�JO���*��2pg��������8�t          kⶔ[?�Y��a<��.����A>�W�         ����=Zq����_�.a���斫�"�`���t          ��1h]0}����t����5u���?�8�"�J�          ��n�<8zq�oJ�0>Z�G����s4n         �gDjݰ<����C.��&���v�S���t          �y�>w���O�F��;'m��v��u("ߧt          E|%��f��t��U:��v�����         L��Vj�?�}�}K�0��9ay��٩7F�ݥ[          (+Gt[���Ggwؖr�R� FS���ڴ;#�J�          0T��:X}��Ç�X:��c��q�۶miZ��io�          �ҿ���9���/�a��J0Z�g6����          ܍=S�|��۫�!�w�Y޵�fepcD<�t          C�~�����e׶�!��T:�ѐw�w��|c����-          ���D>7�z_/��s��{��:�^�����         p�D�)����a������UuJq}Dz\�          F��uZ�4?���!/ܹK����5��          ���6�|cޱ���!/w�T�v77�>O(�         ��xx��zm>���K�0���y���� :"�-�         ��yd3=s}޲��!�T:����^�����-�         �8K�Ym.J_��m�K.��my߾��-���q;          �/?�iO]�w��T���a�NDD�v�x��9�n         `b\�����{�̔a8�s����>?Y�         �ɒ"=���t��;�/G��������-          L��㢕���s�T��2p�`9"5u������-          L���╹�
#��f�>�rDj�����gJ�          @DDNqIS��#ڥ[(��}�>n��AD�\�          �O��T�����D�O�~�}kD���          p.m��eF��>a���-)�kKw          ���/h��9"�.a��O����S�ו�          �c�^����JW�q�'�r������;          ��xy�~g�6�s����_̑�^�          NT����kJw��\ps��~�q;          �.E�Ŧ�~�t���1֟�<R~w�          X+)�;o*���0pS���"���         �1�"��ӛk�֞���W�"�e�*�          �!E��N��;�;X[�c�_חF���q;          �-G�_����[:��c�>F���)���.�           G���^Xx�ֆ���X��KR�+"b�t          l�9������J�p�����\���'ø         ��4�9=ofq��C89�#n��~"E�TDtJ�          @A�9�sgz������f�����U1S�          ��j���^��C81�#���s��FĦ�-          0D���3��gK�p��GPSU��HWG���-          0���ȗl��>W:��c�>b��zL�t}D�V�          �X���⩅�kK�p��GHSU�ʑn���K�          �XJ)��YX8P:�cc�>"�u��ȱ?��         �xI��������!�3�Я��E��#���-          0�nK��#��/�y������C"ǁ�8�t          ����ъ�����t	w�U:�����>8r���          p��b�?�߶��K�p�\pRG���)�P���t          ��[#Ο^\���!|/�!t���?�8�"�J�          ��zn�sg����tw�*��v��s4n         �usv䛗���[:�;r�}�,���l�֡��U8          &�Ws�3���ϥC���C�HUmo���0n         �����Z7ݾ���C����8R�ݩH#�}J�          �$�ukup���ݥ[0p/.o�:;��ƈ��          ����^=��mۮ�!�.��dyvvk����(�          Ŀ����7/.�k�I�{!y۶-������          04v�S��۶o�J�L*��g6���づ[          �;�_gup ��9W:d�o��k������xx�          �NݿiV�[gK�L�T:`��ݻ��,-���t          p����⼴��o�C&���ɳ��6������[          �c�w�V:/���t�$0p� ��NiR�.r<�t          p���3�>?}�K��w���.W�)M�k��         `d=�YY�6�}��CƝ��:����&����-          �Iyd3=s}޲��!���}��{�����8�t          �&�tf�˳���W�� ��;�r˭�IO.�          ���ئ=ue޵kS�qd���}��[����[          �uqA�߿��}�����n4G���-          ��I���o�����)�2N��H�h7U�'�[          ���r\���ty޷�S�e\����j���"ҳJ�           '�x�w��1U�e�������}��9�[          ���S\�T���v�Qg�~rDj�����ť[          ����T�G���I��;A��ۻ?W�          
�k��eF�'�����[#�ϗ�           �I~ASU��t�(2p?�u�����;          �a�~���w��E��iy������;          �a�^֟��Y�b������)�Jw           # �+�U�������5u�����{�������{��g8�z�oZ�%QR��֫�:����(�] H
��&m��i�)РF�I�4E�^P�]4��8�^�+���^t[�V�V���;���~��y�ɱV�.�g漜�|������ ��{�'�G��          �W~����!W)�u��A�P�/#�           ے$����q�sd���]���E$�?�u          �����&�~��9�L��g(勿��^��          �$ҿ�0>�?�:GV)n��|�7#�ߏ�\��           �F������k��d����(
�i���          �4�������Z��OX+����/#���Y          �}+�4�ۍ��W� Y���1k�¯%i�QD��:          ��U"��h���Z�
������$����          ���H��כ&F���A�@�="��_���?���Zg          ��4ҿ�4>�ǵRk��^��4��i(�          �SN#��������Aj�@������H�MD4�:          p��*��Z�����:H�؂{yp��4�}5"�j�          �R.�_���Z��Yp/��?�F�8T�,           ���$�+cc/�:�^;p�r��4��GD{��           �˷K�/�:�^:P�R��L���#ҎZg          ��夒����їjd���{)�<"�fDt�:          @u�����GGP�${�@�K��c�Ʒ"�H��           l�|Tr_j�y��Av۾/����$���u          �m������:�n����|��$��I$��          p�f#�_l��AvK��v�j��@ɋ��          �>q8"����чkd��˂�j�x�����D�:          ��Mr/���u�ݐ�:�N[���E�RD�u          �]2�F�Ŧ�����������P]���          ��֟������'jd'훂�r�P���ň�x��           �4����xq���t��E�=���O�q��Y           ��Ѻ��W�kd'�������\��BD��u          ��Kr�/�k�^���t`��\_����L��           �������Z��m�==v�����Z�q��Y           2�3���i__��lWR� ۑ�8�Y^]�fD�Wj�           c�nH�&cc7jd����':�+k�Pn          �T����fZ,v�:�V�W������Z��H⳵�          �a�ʕ�����õ��M�=��[˹��>[�,           ��'�������:H��Z�F�Ϸ�#�����          p�y��\��dzz��A�&�;���N5���_�r;          �v�\���i[���M����7��W�U�Ɨk�          �>��r]���ǎ5�:�ϒق{��Í�s�o�+��          �|�TZ��,��3YpO#�ʳs�F���          �_$�>W*��$=u���Y>M�
�iD]9_����J��           �7I$�����G�O6�:�'e��~�ܞ��#ҿQ�,           �U�__����4���Y>.3�4"W.����o�:          �~�����?�R�=�4")�y���:          ��r����<D���I�'��          p �z9_��,��k�V����D�Z�           [���|�_�I-SԴ�^��7"����           @DD�[�|���2A�
�k���D��k�~           >)��R��Oj������]��]�w          �3���J���T�W�y������$��f��          @�~g-_�o����^��\(�N�FM��           lM��?l��{���zQi���"��W�          ��%i������ݓw��KJ��oG���^�          ���D�_5������]V�+"���x           �"�H�q|����Kv�t^��3"������{           �uiD�w����n�`�
�B��#��3��          ��4��;�c�b7�+��B�+I�2"�v��           �L%���Ɖ�?���x�}�P��$�?����~6           ����ɯ7M���N>tG�k��_M��#�a'�          @�l�������?ީ�X�}}���J.���hکg          �i�4ү4����x؎�˃C��&��;�<           ��J���<>�g���{.����/����Pn          8�J�$~�~l����!�Tp/>�&��FD۽<          ���Z������ѯn��.�����K#�ZD��3           �W��$~�al���ܼ��{�P�\���#�};�          �o-'��5L�����\p/��OD$ߌ��[�          �a)I+_n���w[�iK�R�p.��VDto)           �|��GG_�����B����#ۊ          �A3i�K�#�UsqU��b񑤒�=�          ��f6"�����7�v�]����Iķ�Hv&           �tZ����ɫ?�Y�~�W���"yA�          �{Л�6^X8�.��;�����*�ӈ��g          � �J#�b����O���ྒ��U���          �A��H�_�?z��~��
����P]��v9           LQ��m������?K>���B�X�Ʒ#��^�          �@���V~�eb�ʝ?���=���O���          ���Kr�/���A.""���+��+"N�,           ��������$�-�սi��u2           ���_HJ��X��           p������)            W�            ��          @F(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�          �	
�           d��;           ���          @&(�       ԅ��    IDAT   �	
�           d��;           ���          @&(�          �	
�           d��;           �P_�  ��ب�����X���ήXik�Ֆ�Xk��}��-J�MQnj�4��4I�����r�mlDDD��jD�PZ�敕h^^�敕h���}v.��E�͛Ѱ�V˿2 pIs�X>t(nvu�RWW,vt�ZKK�����~�+Mr��P���0J���DDC�u�rԭoD����1��qJ��J4--G��B���š��h]\��� �߬55�bWW,vu�BgG����jKK����ZkK����zCCDQjn���J]]��qm-�4�$M�a��|I��J���D㝹���h]Z�5�27���7�c  �j��%:;c��3::o����YZ���4�(��l���z}�_�]*�hX+EDz{M�֘es첸���o�]nތ�� �i��r{���e��cs�rg�h��5*�X#*76F��ֈ�ף�������4/�D���ͱK��RD����l]R��_ ����������}1��������ˇ��<K��J�������==�SS�}�Z�..�y  6��b��7f��b��7f������X��Jno��[_����蘙�#���=u-��]����H*�=� d�Rgg��퍙�s+�==���kMM{$M�ui):fg���tt_����hS අ����5n����#Gb��3J{<vI�4Z�cf6_��y����6D "��F �==��,��]n>�Q����,u��qh~>:gf����>��ttܸ9kD�I
� p٨��냃1U,��ѡ�����ZǺ�������ѱ���Q_.�: ����B!��ŵB1�t�y�}���ף�ڵ�������= اJMM15T�k�BLō���/�oá����������)�� p ����T�׊�[c���=/�oY�F��\�E��X\���_��   7��o�Y���Z�sG�d~��nc#O]�5�2:##Ѻ�P�X@(�@���\\��c����냃�G/��r�J����+W�x�R��8� �S��b���;q<��Jkk�#��ٹ��ŋQ�t9���k	 ؆rCCL;�'O���p���D�$��u�J����GE���虚r�6 �����8~,F�����1w�H�>�4��E����˅螞�u$ `,vu�ȉ1z�D\*�J[[�#툶���:�K��x�r��	jB� 2f��-FN���S'c���Xki�u�]�P*m.��p!�nެu$ ২������=y*FN�����ZG�uI�F��D]�C.F�Ą d���#q�ԩ�R��y]-��Q�t)�.^�Ѵ�V�H @�f�zo�]N���P�w9�	mQ�p1�.]���K�P*�: P�J]]��ة�q�ĉ���u�]��i����K��������	w Ȁ�������31~�h�;<y��������������а����w�������Q�T�\.G�T�r���뵵�X���4����8��{q���~���r1v�x\>s&�<�`���Q�uuu������Q__����c�;c�\.�9n�ccc#�ۓ��||�����y�Ni����'�{/z�'v�� �����O����L_ߎ>;I�hjj������[��=����'�V�4���'�mll��x�Θeuu5�����؈¥Kq����?�Few Ȝ�ޞ�|�L\<}zǋaI�Dss����θ���>�n��$Iu�����.���c��Ϸ���l�����(~x!N��~}�a���� �7�\.Ə�K�OǕ�����}~]]]477����;㗈�ֈ>�g)�J�����kD�q���q����l̆H����F6����Ň�<�ǎ����������hii����hnn����N�T*�����������p��I�F��H�z��8��,���V(����G=xϧ�$I������)��4Mcmm�'�*������+++������8����3o�33;� ��Jkk\x�Ѹp��10p��kjj����hoo���֟��)�����O�[Y\\��Y��z/^�ϼ�N}�a�*�J l��C��s��Ň��lｗڛ����إ��y��.w>������˛�,KKK���/����o��K�"1v�����o��~(Vwh���Wkkk477Gkk뮯�J�X^^�Kc��(�������ߏϼ�Vt]��C��;�`������?>rv�E������舮������,�e���j,..�͛7cvv6��涽0�P.���(���76��I�;�ZZ��#g����c��w[ϸ3Qyg�r�Ծ���۱�����������������=,M#�j<������Qw�� ��K�$Ə����+>�O�<Z����ͱJggg���GCC���7i����J,,,���|����͛7��͢W��b|歷��7ߌ���N |�4���'�'��S����QSSStuu��Ç7K�Y�,//o�]���b~~~�ű��7��7ߌ�|+�n��� ��Ykj��><���O�K�$���~b��5�����M��Y��F##��?����;|�T
� �*�\\>}:~��_�k��ﯯ��ÇǑ#G6����5�4���Ř�������~���
����q��Wぷ߉:�0 �q}` �}��|������/I�D{{{���n�v��ݴ��sss1;;������ye%>��[��+�Z������x"�?�D,tum�������������ꊶ��]H��*���F7n܈��٭��4
}��j]����`ǭ����O>�x<��۷|SSS�����Ç���Ù���ԛ������-ޓJ%�.]��_y5
�.�RR 8�nĻO6.�>��X���舞��8|�ptvvf�x�*�J?�gYZZ��3�����[o��W_��ٹ]H	��; �RSS|p�\��٧b��sK����Eoo��?r���#��4�����~�zLOO����oYZ�ӯ��_{-Z�ᓴ p`%I\=y2���31><��[���g�k7�������ͱ���̖
d�J%���~<���G���.���k��+�}����cQnj���$I���3zzz���7:::v1e��o.�^�~}���~=���w޵�  ����x�����G�R9,I�8|���<K�6J�������q�Fܸq#�]�kkk[��{j*����{�E��y po�$FN��w�y:Ǝ�ҭq�ȑ�N�~^#�q�F\�~=nܸ[$�J����}?���v1%�_
� �V���g���O<�-,����EơC�v1a6������DLMM��-�vZ����v<��w����.&�����ŅG��?�L���T}_CCC������@9r�<Q�^���ǵk�bjj*�_����{�������>ڽ� ��������|\y表T���$I���+���?��0'�_������dLNN���j���,-řW_��_}5�X4 "�����?Wx �*�K���������t��l�499SSS[*��.,���g^=���]L	 �O��Ņ�g��=s��U�������188x`׈�_�[^#���^�n�pa���� ;h��%�y�x�OE�ʉ����(
188�ow�؎���������Ѫds����r�..�rB ���I��>�?�l����$I���?��|����	˟�\.ǵk�bll,fgg��o���x�b���]L �����x����ӧ�.����E�X����Yj�i���c||<���c���ٛWV��}/μ�Z4(��]����k?�����U�]��ۣX,�������t��4���٘�������wGm]\�G��r�~�N���H�$.�9o|�٘?r��{�$�����5�\���w155ccc133S�}}����K�_._��t�(��(55ŻO6�}��vlO�$�9�B!����~�4M�ƍ122��ӑ�w�ԯ���7ވG_�n�,-�AJ ȸ$��=��٪w�hmm�b��B�b�],..���X���E��"X�ҥx��/E���.������������ųGZ�bi]]]������Ptuu�A�������&sssU�Ӳ�����8���b �)�z{o}(�*�������`EGG�$�������d���T}�o��B��w߉�|3r[�M �$���L�����پ����y�	����r������x�'��	��� � ���s���_�b���������(�144�U\�OZ[[�����R�t������w^�����*w� ��f:�����sq�P������8v�XtW��;�R����T\�|9�~C�����}�h�r� ��RSS�����ݧ��J]�]�oii����(
Q__�	����Ÿz�j���Uu�����x��ߊ����A: Ⱦ���x��<�xT��P^[[[G>���*�:���7oƕ+Wbbb���:o܈g��f]���  �����瞋�b���{zz�رcq����i����T\�r����� ���7�}����Qp�m���=������MMMQ,cxx8� ��V�Tbrr2.]�KU���1;O��b��=H ٰ|�P��/�����.;��r���ǏǡC��(��6;;�/_����^[_.�ï���h��C| ��IΞ�W���+U�?:::bxx8���J�R���ŕ+W��]�o|<���7�oll�@�Tr�����/~1V������+�����CJ�R\�z5�^�Z��y��>������b^ ���5�s�����$Ibpp���ʇ�r�J�~��x򥗢����Pp�-Zno��>�\|t���^���'O����K�4����p�BU��._����עcff�@mTr�x�s�ě��|���������cǎEcc�%<X��ŋ155u�I̶�����>���G� �6���/�rU�tww�ɓ'�.�K666bll,.]�tע{����ߌ�^x!�VW�(! ����c��/�R�����ڞ��8u�Ttvv�A��gcc#�^��/_�k�=W�ęW_�'_zɆ �\.�y��x���G�.�>uuuq��QkD�hyy9.^�XUѽuq1��ַ��;��Q:�>w �V�ćg�����R�����K�����ɓQ(����yp\�}'�ﹽ�@7���  �$@-$E�vK�i˒��e�H ���o�R3U�^ޛ�yy%˲=���Nfۙ�%oZ(�)�ľ;�h��z��
�Ⱦ�"ٷ�流U�s.ȯJ���9��;�,l��ӹ�BwM ��'N������(�#""����l�q��r7}N���|TTT�`0D)]rs����������c߱7`��|DDD�$���܁�x�[v�Z�(--EVVV��%�P(���IlY螲����}��.E)�:�>z���j�8�Z�����KyQ066��Bw��*���&�{�P����|v6�{�q�n󌨼�F�1J钛�����0&&&�,t/¾cǐ���tD���DDD۰d��wO<����M����(//Gaa!�U �2�����ߏ�-:�e�������T���>�gރ��{ڤX����[^^F__���6}���b�o~����-6;�����XE9��Q�n��4--UUU�o�C*�z�`�/_���0�[4(��ž7ބiu5J鈈��g��|�3�7}�b����QJF����122�˗/o�v)�ԁ;�k�x<QJGDD����wl댈���Y]]E?�N���|>4���>:�3"Jb,p'""ڌ��҂��߇�V��c���(++�N��b@R122���a���I�O|��ǏC
��������q����>��-Rm6jjj����d��Ӊ��^x�8TͿ|�����NDDq�o0��GF_c����zTVV�6���z��ߏ���M;��^���_��"��Qb��w�?�ᚚM�3����D^^^���f�����ۻ��yF��Cq��Qbp��]9#���͆��j���G)mfnn===Xݢi@��8���O����dD���DDDxRSq��'1^V��s����0�7��Aѷ�����>Lmѥ�19����ߐ>?�dDDD7O�$�߷��ߴ#GJJ
�������t��,cdd������gX[��_CiOO��<gA�~�i�dX#>æ�myy���X\�� ���������dDDD��DI	�}�)x6i��hPRR���h7i�D�XXX@OO���7}���y��_A��G)ѭ%K��}7��s`�3"�Ʉ��J���D1m�,���� ���It^/���Py�b���)+/�{O>��Փ�555�"���	���m ���B����������Y�X���Oc��0�3B�����1������g�.c/aߛoB��E)ѧ#K.�y��{驪�iiihhh�3q`rr===�����p�O�ܑ�(&#""�y!I����p��ț�$����;v��QGOO��`�g�q�����QLFDDt����Q���������k���8v���(%#R܉��>!���ÇDWs������_�H0��� ._�����e��8��_�kŬ�5�8����IOOǎ;x�d����Aww7��t>��������(&#""�>Oj*�z�YLF>d�h4���Baa!�&Ed[�^/���133�
a��Ǳ��	`��""�X�j��7�{�M��t:TUU��� ���f������.W�=)���v��ŉ��j����gDl(�\.�����I{�����}r*�Ɉ��w""��yRS���=��M6(SRRP__���dt+-//���+++��p����QLFDD�9Y�p��A\��. B!�$I���Dqq1�����Goo/&&&">���p���Ү�(&#""��ta!�z�YxRS#>c��QWW����(&�[��t����Mn�)�������M^�#""R�xy���g��ɺ$++uuu0lRDF�mjj
��ݛ�DSq�����͏��(Fɒ�3��gD())�Q�
������h���4� ���KT�?�dD�`�;�w ������:�t�(&��A�ebhh(b7w�׋�?��{z�����(�zJ
�y�/+��Ljj*ّ#A8�NtttD>|�e���C4��D(�pDDD
zv�GAH�Q��!kb��|������L��<��ᜍb2""�m����$)>��h�6�������/ba��FV���ǰ��E1��xF�|�����с�����T\�t��@ �Ɉ�K��ҏ����HM=�w�瞍x��N�CCC***��pHK�E���Պ��9���g�Z-�kk �ccюHDDt�B��x�E�rs#>STT���&��(&���l6#77+++��Q
���B�����DD���F��O>����G,KMMŞ={��������h����^����ޔ44 cnVň�(6t:���3�ji����b�����#���v�j���˃F������3�&�a����DD3�{F�s�N�%�Ʉ��<��nx<�g泳1YZ�~�|���܉�(i�B���G��9�&��jEKK�Vk��Q4�L&���ceeE�K��*)�J�E���.eex�����N�]�v�����b	h��U����V�V�TU�hp�M:y�^����0R]���B�ڵ���	�b� ++��|a�!�õ��y�Ȟ�P!!�ﭥ���/}	��%�)))�Ν;��룖��C���8���+ޚ�j1�cL+��OO�������&JK��6?#jjjBqq1�M(~}���\�f�����A��e#��3�QR
j4x��г{w�g


����N�dm�fˮ��٘,)Fq?�
�DDD�C�Νx��g��IOOGKK,K��Q4m�fdd��r)�<�5�0�Ѐ��q�./������ъՊc/� W^��$I���Cyy9_�Kpz�����x��P    IDAT<X]]@L��Ó����A6 ""U,:�ŋ/`1BWv�F���F���p�����"6?���hU�����H[�����(IX,8���!�p���hDC=2g�a�-4�`X�NDDIg�d_z�������<�M2HOO���B(
�w[,��DQ� �^�
	��(i�3�݋�>񖙼�<455��XIIIAnn.�UX�t:��@���K��ѭ2���c/���7ޥ������d�x$IBNNΦ\�9���Aq_$��""��e��o���O�f3���a�٢��Բ�U�刷����c9ӆ��~��GDDѳ�3�]�v�(����byykkka�!��uuH]ZB�өBB�ۃ�DD�T<��8�⋘��Q�7�hii��n�r2�f�999p�\�WS��L��AQ� �
_���n�8�Gp�;"L��֢����M&!�V���<x�^����͇$	�55H[�&�>SE�x����MIQ���lhii��d�r2��Z����Ul �����B���B�p3ѭ6ZQ�_��
�����g���('#�	!������t���BV(b_�ʂ+7%=�|A���n?!p⑇q��;#L�����(Ii4������cii)l^�$�TW�����
	�n=�Q�p[,��K/bɞ�8�q���l�r2�%:����X^^V���o0`��×��v������,Ix���г{��V��Ν;����dK���ʂN��ܜB�v!0R]�wY��$"�[k������7�7n��h4QNF��d2!;;;b�U�e�(��Va����V���o?��Z��|AA�vIrf�����a��6f��Q�������Q~~~��Q,B��p�h4��r)=���r �##Q�Gt�������ªՊ_��"Vl��v�{���N�ʵڹ���z�X^^����Q�ܑQ���ݨ�$���O�g���`�U�t��
�٬�aL���A��#{|\��DD�pF++��C�G@�S�///Gmm-D��)��t:���aqq���a�4�VT���:�O��DD��w����>�P�����r���p�B �����`~~>��ɪł��R���@�PODDt3dI»O<���;�yFD�KOO��b���T��f��A����*�#�uX�NDD	o9#?��?�ے�8_PP���Fv�kltG�������V��Z�]�ye5��(��$	�}�Y�S�OMM�޽{y��IMMEFFfgg���l!0QVM0���1uQ����o?��b��(..V!�2�F������­p޺ٌъ
�u�@�N�DDt�56���OA���9I���Ԅ��B�Q,�j�������2�����=ii�,+Eig���NDD�HH��ֳ�b(���l�)2�L��̄��DPam2SX���E��X�NDD	͝��c/�w�rq{II	��Ѧl6�z=�����Z-.�ա`h�U�э����O?��Z����4�ݻ�!��(^����n�cffFqs��:;�ѧ7QV��|�s�ۛ������B2��$!''���XQ��k2a��e]]�JDD���j���ӊ��Z��v���P!Ń�~#���IM�tI1ʺ��a�;�$Y���S �������gD��hDVV�N'
�*3��2�;:�B:���w""JXkf3~��X�pMSii)��������b�^����
�j���AQ� ��
鈈(n	��}�;�-���������`@VVV�"���R�VW`��V!ų��B��_@@���h4,�mٸ%���cii)l~�l�TI1ʻ�Y(FDD7e��oEx1O��bϞ=�E83"� �@vv6���_�s��c6?e]ݐ��Q���h��������v*No����(�x��둝���}��Z���(.�����ҺɄc/��E�]q���
QNE��b��d2��t��t:�TW�����u�Q<����ݼGq�f����Z�b2"%z�YYY�����c���#cvV��DDw���x�K�ïp���j�{�ndff������@0���b؜'-΂�uu�P���>���2����T�K��thii��bQ!ţ��"�B�b�b>'�]���BB""�w<�0�[��xFD7J��!;;.�~�?l~��&�*�Sl�D��DD�p�Z-~����U�������QNE� ---b���`�XY*:y�6m�¾�q~�>�9�͆ݻwC��m�h3:�YYY�����.F���=6�4�ΩDDD��d�ፗ^��h��(ng�S�4�v;��b'�U�vʺ�!T�FDD�k.;o>�E^���thnnFzz�
�(�mU�d��m����_�tDD�.�}��߯8�3"���Z��N�aE�B`���',ss�$�X�NDD�E���S�Н���eeeQE�$--F�Q���k2�Y���NH��ADD����GDxَ�jŞ={�qI��F����LX��,I��Fa?R<�Q�[OI�/��B��v�b�v�)v�^����asKv;=
��THFDD�ȓ��c/��u�9ln��<�ժB2J�n����ass�ـ,#wtT�dDD��kk��c�gD����<#�O�E�J���TW#o�2�
/��"�QB���ѽg��\qq1������Qzz:�z=\.W�ܪł�LJ{zUHFDD�n6/�>�y�6'���x�$�:�������F(�f.��b���]���|*%$"�X�j��/=�P�:B455��p��������Q,s������I�Q<�8��XVx�N��`Ϟ=���P!%!�������BÀ��"�-."S�1�'񌈢A����p(6B
IF��P�����J	����DD�0zv��G�߯8WPP����('�Df�X ����|�܂�Y y##*$#"�X����c/���6g6������U�D���`@FF���!_w���h�tQ*.u@�� �����x��Oc��\aJ����
��D��YYYXYY�����(+�}z�}"""�Jq�o>�y�������6���~}1���@��Җ��	HDD1�gDM:�v�]�R@��Di	*::��� �(ְ�����LA�z�YȒ6�p8����p��Ͱ�lX__Ǌ��M�EE��faU��NDD�ǯ���_���z�{��QaS��f�F���bff&lΓ���tJzy�]qa���ܻWq���
�
�cD7C�Á��9x���'1VY���^���	HDD1�������Qqnǎ��ɉr"Jt/�����wݭx�$a���]��_��!"�����N�CKKψ�����X,���
�[7����@YWXIE���DD��RSq�/)�隚��={�@�p�ѭ�p8���~-���@q_R��$"�$"�}�)L���MI��={� ---��()��fh�Z�^���Άѳ��
Ɉ�(�L����O 
�
QUU�B*J�$!++333���ZL�����%v#"�k��T���+�]���Q��Ct+h48LMM!x��$��a���/��<""��-Έ���yFD�MJJ
�f�b#���LH����Q�m܉�(��$	�����p���F^�D��f;B&KJPu�W;%�Kw܁�;�B���v�]�T�L�V+�~?��ɞ(-E���H]^V!łU�o��%�O�v;oţ�N��"33S��l�Ʉ�Lʺ{TJGDD�f�a�/��E��ڰ���\��֪����N���f���dY�fn-5k�T�������bψHm��� ��������"8�&a��#�,p'"�����cXa�R�Ѡ��f�Y�T�l$I�������A�͆��%���b���S���*++QXX�B*JFv�]��Y�0^Q���|~���ZZ-����X���3��hii�$I*$�d��둖����鰹E�Z����*$#"�X�3�Ƌ/��q��'Y,�ڵ�/�QT�F�L&�n�s�90������!"���3"�6�n�����N���r�uwð��N8�Mpg�����HU:[�����x�EUJJ
v�ܩ�y~��ݻw�����Դ������,B
EaYYY(--U!%��n0)))as��T�)ū݉�(��z�~��䄍k�Z�ڵ�F�T���v;����N�f�r�����b�����l��q�^���&��GQ���q�G�����DD�<xFD�����j7�O�n�w�Hm�[IDDqi�l��{Tq���yyyQNDdff���Bq�Ç�<73������~F����dB}}=;�Q��t��Ŋ��e���(%���2t5+��������*��ˑ��6�$���3�*�""�X0\[�����q!`4UHEɮ��v�=l<����<��V�B*""�<#�X��h�k�.h�'��|�߿O�TD�c�;�!��SOaM�ˀ�jEMM�
���(++CVVV�xP�ŻO?���%��]M���膪��THE������Vq����yDDIb�lƻO>�x{GYY�b�1Q�Dz�b%#>��
���Hm��{�qŹ��*�c�h����,N�{P�TDD�6�Q�2�LhhhP�;�?f
���hs,p'"����Ҍ��q�N��;w�MWR]}}��f�\NN�wo�QT-�l��窫���#����|���Z-�fw1"��'�{��"�LF-Z�6�_oS.�T������"K�y�)�n���())�~(�O���hllT\�t�q&JKUHEDDj�ź��,��o��&R܉�(�,�l8}���suuu���b�N�CCC��f�;��LA�
���(d!��O��ׇ�egg���#jkk���6�����{�Q!EK�Ν���j���E[ZZ*����{�&S��Z:���tQQظ^���}�(�222PVޜKǟ|~�%�Q����BZZZ���ՊS��<�,p'"��!N<�(
%��򐓓�B("e6��
]9663���(1u77+^�g0�c�)۬3�;kk"���I5��(�����Ģa�!%%%���_7��![���ªՊ��P�۱c�
�cDj)//��jw������F?Eψ(^H���;wB�ф��4��oI��w""�=��Q)))����~ �-TTT�b���/ef���w�����n'wz:>��`ظ��t*�"��b����<l<$I���!$qۈ�(�|��#�*�~������<E��:z��c��]R��(���L�jQQ���TE���E�P��yo�%"Jp<#�xc6�QUU>�q�Q6m�X��J""���T�z@��X}}=�\XQB���^�3��}��ఫ����n��{T����B�ΓD�������a��\t�ݫB"""�]F��0�� @�׳q �,�����Ź�}T�葈�C_C&nI5�L���T!��L&�b����!��w""J<#�xTTT��6�d���囔����DD>x�a��(.��bEjj*���;��4���c�B�;ş��VT���F�RLB`ǎ�/�=x�
��Q���t8��g�jkk�E�bZ^^���&�V+����V"�D����S=�8W[[˦G�
o�]t8p��;UHDDD�ψ(����AR����]w�i#���DD�f
1�Щ�`0(_�Cc��ˑ��6>]X���:ѭ�jq�A�fx�J� ==���a��'�_�DDDt�]�w7�iia��999*$"�1uuu�(t<�hi��_%����zJJ�x����b���b��c3"��3"�wf�Y�i�$�GQ!������b�,N<�b�kv�x�Ygԓ�߇ �ŵ�w܁U�5l<''YYY*$"�qHQ(���ta�
����VY�XpI�S�V�Ŏ;THDt�RRRP��/���d��DD�v���6���Q���(��f�����t:|t�
����v�%���2�)4ǘ,)�(�����Ŵ����S�$f�ۑ���B�������x�v�����@  �ߏ`0x��F���K��A���`0 55f��/|
V�����f�m���]wa���*%#"���IM��}w��k4���`n��kkk���W�0�@ �$A��@��B��^]ǘ�f��f��1b�F�Amm-Ξ={�������}B��	GDD7���#��-����������:�n7�n7�^/B����_�,_�_�����a4��Q�:|ҵ���199����k�G++1^V���!��ѭt�R�\������- ��յ�����C @(���i풒�����ĵ�6���arrkkk׌4ԣ��idMN�����n��z�,_�g�X�|�����Cq��V��N����b4�RdB�����ɓas>� 
!�*$�d�w""�Y>���!�e`��� ���1??���e����������� ==6�6����PYY���i�k�/�u'�ϝ���Z""�}��z}�xyy9�nR(���\.������w�4�f3��Ү�c�F�-H��v;\.�5��\��܉���UJFDD��ta!�jk���f3���TH�<��籰����U��no�Oq��=##6���������裏��>|�A<�7)R!�*/-]�b� 77W�D���vcaa���W�.�����X�����j�r��$I�����s箝>�0��� �L��(����Ȳ������,E��M~>
!`2�������dff�l6ߢԉ�j�"77SSS׌/�l�hiA�����܉�(fu�݋��԰���b.>7����Ӊ��y,--���_������"1::
!��"���,X�Vnd*���(++C__�5�����c�TJFDD�ƂÎ�������(���n���`~~���7],�$byy��˘�� ���d��#��1��՘��[C��� �/]��:�������>�jjj����F�A�����ra~~>�� �2��ְ��v�E3�V�Պ��Ldgg#%%�����f�!;;333׌/:��G�ŋ*%#"��%qe�k���p:�W�.��Y��>�v���pe�Q@���â��eee�f�a~~��qg~>F��P�ӫR2""�Y<#�t|>���177������[�gȲ|�����i ��`��f��ϢU�퐀��*8�ΰ���F͹s�{�*%�d��Oi�G�ADDt=���w�}���:�MMM�h4*%�M^�������n˦�V111���	����h4r�:V����a_�泳Q��C���ѧ����b��ohh@��Kz����cjj
������Z8v;^��,���2���1::
���N���dz�>�KKK׌��<8x}6Q�//��}���333QQQ�B��������!ttt`rr+++a7��N�P�sss���,B��fs���c||<l�8����3g �	��(.�؁�={��sssY$�Y�������!\�t	��Ӫ�]\.FFF���g6�!IR�r�"�Պ�������gς�n�'�m_(���,��ى���[r�̍�X]]��������� ���l拔���j!�r��yA��@ ���*%�d�w""�I����5���հ�l*$�M������BOO\.|>�ڑ  �@ KKK���4RSS�� W��2W�� �ш�޾?IDD�d.;>�PXGԌ�TUU��*�,..������p:�Q9/�P(t�����ujjjR�n�^��<�����g Eqә��>%!��g?OZ�u��v�^��l���122���cii)�����z�p�\���*L&S�6��t�X\\�f�g4¼��uWiQ�%	�}�xM�k�%I��ݻ�a3�ߏ˗/�ҥK���rTlf}}�������lN�5�^����:����_7���r!��.�DD?xF�=�������VWWՎ��ˁ�333���GZZZ�7�`�X011��}.75g�Bŗ(��M���bΚɄν-a�F�*$�-�,cffCCCXYY������, �ǿ�dY^B�HB�AKo;    IDAT�Ȓe���F����E,..b`` ������O�B���l����mf���c��އ康a��(����`��% vC݆��y�u�A~ �B�iY�� V,!ܲ,� 0˲�*�HB�>^�Xo�q�������� JJJPXX���:�%%%�fܓ���={�p�JɈ�h�F+*0��6����.b
6��65o��0�% ˸�ײ
�+�0˲l��+�+y J ���i0������������RX�7�̉{���;l=�*/\��q""�m;v`�n/((��hT!Ql�z�W�.�� '��]Vpe��*�p�˲l`��+k� E n�@0���&''������R����L�T^^���ɰ�'��s �==1�R%mψ6������aLMM���w2�1 㸲��Q��eYH����z%C�e��@΍�!>����E~~>JKK�~���hPVV����k�}:�{�~G�`���T����Nǝw¯�š��<�:g*������ �n����4��dY>%IRO 蛛�9z���}���.
�U�,W	!��`[w�z<tvvbpp���(,,L�B���
�={��1Y�pn�~��ӟ������Õ����ʰ���L�4����9�u�܆E �eY~_��^I�z4���Ço�����fV0��$�J��B���m�g}>���0<<���"���$|�{qq1FFF�.�}jϜa�"�w��=acB�^���chh�����g[�% o�������/���o�ꫯ$I�BT!�eY�/��W�l��t��t"33IU��B����5���t�55�����э�%	��96��hPZZ�B�����088�����e&(��9!�;�,_�e�����~��_��M��~��Ƶ��*Y��$I��B�� ���YY�1==���i8TVV"�ۆ�F����k��v�֢��S�dDDt�xF���F?�N����P��w%I�
�B}Z�����Þ�M^}��t�FS-IRU(�pPтm���A���bllyyy���Lڛ�+/��ݾ��܌�>�!Fne��'|y��qG �����x�[(������I[�v����u#�N} ~	���$�}�ȑ�ە���_/ÕB�<�mld@ZZ������z'O�+�B!|���|s�����6z���bpǎ��;��E�D�m}}�������p����F��f;w�С�҂���F��� x��v�SRRPSS�����+f���/l|��7Ps݋zDD;&KJp�������Q__�B��499���^�|����4��e�-�V���Ç]�#�ѣG��c/�� <.��k;?'�@AA*++���nG�����q������׿	���Q]���o�{.l������*$�=�,cbb}}}۾mF1
���,�o���wo��}�~���N�B��%IzR����̇��"TTT$|����x���^N�OO���Rэ�Q�`0���!�Ha{��'�`�m��w������nG��|�;i^��Y��B<�l;?��hPQQ���⤭SG��Kx�o����O����܉�(�tܱ>�P�x}}=���UH��@ ���!\�|y�_N�~(���v���來��?'��2�����d<|�$�˅3
�?� {��
���h+n���ކ�u����v�ٳG�T�I�e���b```�Q{eY��V����ÇG�~��������{\��/x@��B�q8����ɴ����N0�����
�,ss�ܷ�͢1"���/~c�ujB���HIIQ)U��&k ~"I�����u��Ѩ_a�o}�2�$�x��mlu:����fmppa����(��U!ݨ���`����1�V�@�p�o�Y^^FWW������*��
���r�޾�[|o��^{m�$I/	!^�e�`��F#�������x�������H��c��OȻ|9�������(���DOO�ֶ�O�eyF�?��kmm=�x������_�'IҗeY�<�-�1&s�FY����ϵ��M�����_�&x[zS]��DD3B����b�����`�����ȥ�%\�pa;_| ���h���Ç{�m[���o�W������z����p8QJ;N�8��뺵�^|�կC�������"9�Ѓ�t�a�{��EFF�
�b���Ο?�����q�h�9r�(Dۖ�^{-S����,�_�i�v�F���jF)]tE*{�?B�Bww""RעÁ��\��������F�R�Y�1<<����-�|����j�ڿ?|���n��a�B�{ �l�|FFa4��N=���g���ɿ��R�v9
��?����"��֪�(vȲ�����vBB�������׾�F��=zT���z��Ǖ�H�r8hhhH�fH���8~�xؿ�<�V)mψ~/���s����B��333?S�y���~��F��sH� l��,**Buu5$i��	gtt���a����稺pA�D�lX�NDD1c��o=�L�xUUJK�lP�P._������6-=B��������W^�V���k�e
!�T�l�lII	�����e���)\�x1l��_�'O�����"���+_��`�f<==w�u�J�b���4:;;����e��eY���_~9�~���o�
���,�`�
����ر#����|8~�8��u������J���(���������.�����(6�|>\�t	.�k�G �?v��{��m��Z���o5���B<�Mn����hhh��n�b�������h�@O��? {<f�̈��o�{�kk�B`���	{[�v�����ŋXXX���. �t:+�bJ��o�B�%�G7{�h4���1�/^�����ke�������-׫DD������2Ο?��f��H��9r�����i=zT���~�_ʲ�{�g�����ԔT7$?~~�����,����x�/�f,p'"����?�2���|��hp�����ذ����ҥK�����1��	!������h7��W_M�j������/�b����)�;�m�eǏ����5�i��8��!����(ft�4�Ge666"77W�D�%
���ccc�>'��1�F�gG��R�����P?;;�.��� �"=g2��s�΄+ ���R������-2gfTHDDDJ�F#���)׽le����ҢR*�����ҥKa߻�3�?����:t(n�W~����_�e��H�!PZZ�����m(������{/�QDyg'���S)mŝ������.����hj
a/Y�\.\�x1���:S �����P��ݴo~�{eY~@�ũ(--Mص���2>� �"��3g��7UHDDD��3�+FGG��ۋP(�DqI�寴����h7����3�,�5��H�h�Z�ر999QL����~��?�����˗���Jrݙ@DD1k�n+n�����)n_]]ŉ'�*n� IҾ���O�� ��+�,������Ph��x�疖�p��	,..F3�j�(.�~�b�b��$����(�����FcRmbE���p�ԩ���Ǆ϶��?O�� p��!_{{�_�� ��x<8y��v��%%%���J���H=�a������'���1�>}z��v�wB�Pu[[���Sq; ���]<r�Ƚ�,� �}"Y�144�3g�lu�N�JIIAVVV����j�'QW5"�x���V�$��exxgΜ٬�=(���������Sq; ����r:�w
!� (���e���8�|�mr�"==���a���$ə(Q<J�3"Y�q��%twwoVܾ*��I���[q; �����F���W o��p�����NEEEE���I�R*E܉�(&��ޥ8�T���q�ԩ�\�eY�s���|�ȑ�q��_������3~��O�ު�?a@�ф��h��(v8��1�p��%l7��Z[[éS������\)��nwmkk�F1�-���|e���틒$=`D�P(��/btt4��n����U����������b2��PX�$���tuu�u�� �r�F��_~y.��n!�����= 5 �6�ssss�裏��)��ƽ������V���z��VdIB��ư���tX�V����g�B�sB�����?=|�p�M�Xw���Pkk�7�5 ~�9�ӹU�\SZ���֪�������gD�@ gϞ����f��<Զ����Ç����Ç=mmm��hv8���atttD�wJ$�A�E��5�� �f,p'""Յ4ԇ6eff"%	Csss8}��f�t}�,������G�M�V[������J��A�;w���QN}Z����a�#UU�4FD#z^�B //O�4���v�ԩSp�ݑqI��D[[���}-�C��ȑ#��h4;�?V��e���	���P�%�ш˵5*�!"��9
��~�ZPP�B����bppp�G��%ޛ|R[[�B[[۟!��x-���2N�<	���t���fCjjj�x�.�DD���2�-���d\�Ȳ�����(�G����fkk�h��Z[[�mmm��Iq�haa'O�ܬ9T�r80a�M;UHCDD[I�3"�ߏ3g���rEz$ ��v:�O���+	S�q�����yP���@�e���Ν;����|R~~~�P4�����T7\S�5�)l<62���q�̙����`04�����f�h9|���n?(������,���s��݄�T4�j��РB""�$���Ẻ��,Ń�d�����!����ȑ#Ǣ-*>�t�ȑC�,�9"\U9<<����('�="��
�������G�0!���S"�e.\��˗#=�𿵵�}���}5zɢ����_eYn�X ��xp��)��&�?�Ra���g�1����F�I�"�O
�B8{�,&&&"=��P[[ۗ>�xo�hoo���N �J����֢���B(��Nb�nW!E��gD^�'O����{� 0,�����~��ѣ�E����ѣ����� � �X�?;;�U�OB��l0��a�J7J�J,p'""�)�ѧ��;Z'�˅�/F��($��Ӷ������x%�٢�СC����?�e�y ^�gzzz6��MV�U�A��5�DD]#����ta���2^$n�gϞ�������<��ښ���J�ײ,�`N陱������Hr�� +Iz}<Q�j��	�Q#;;z�^�D���������b<������(Ǌ���������eY�'�y�׋ӧO'\�X~~������l@DK�F#�**��sss��hTH�Y�q���ͺ�Ȳ������h�RCkkk���n�S����5|��G���ĭ����l|DDc���(�̙3�����������z*�������F �%���4����s��E��IJgDY�rsUHCɂ�Dq&���o Rr�`��4l\qS'�,..���>Y������j�s��������XV�������l�SE�җ���l,�[�����V�v�[f��6l,%%���*�Q���:N�>��]��������ѣGQ�������, 0�4?<<�Y'ٸ��a/���G���`@0�
i(�W�ï�_�l�����"�/�r�$I���(D&�?��?Zokk{	���4��zq�̙�^X�;�f\��AH�q�/��� �Y(���� ���N�"��uwwcffFqNqV���ooo�r,�|�k_s;���dY�;����5�>}�@�l7�L&�l���: ��H)�$	^���)a$�Q(¹s簲���G��կFl�h^y�����{ ��4?77�Y�˄���0ψ�6�nQ�b�n�rf&33����UK:�:|�O|P�^h�~h�~��W`�����u~ֹ9�..A$�'%���Պ��|�����s�"m¹eY�\{{����Z[[���׿�_�Ѽ	���׌�ٳ*%��rss�����g����S��DU�$a�fÒ=�6ە���	Oj*�:=�:�5�5"�������C���.,ss���>7�OBެK	�k4*�������/�E���q������yt�u'�ﯪ�� h4��b!� IpߴY+)j�i�v�ĊE@fƞ8s�Λ��s�e�L��-Q��O^��S&/NB-�-��%J�$R"EI\�$@����"9`�-� U]���s�ϯɓ�6�������MNNR/'�����+tvv~�{���d�e �+X�9M��l����ב�hi��}o�c�R����/�+���H��	��iӭ�T
����Ih�����C��/�,�}}�I6���s�l��+�Fk�3g���ɓf/��L&������<A���3�<sJ� �I`�����`ժU�L�-++3L�pa�T�8aST��t!0\P����/��"F0�����!�i�<��žP,-G���}��Β���訍�E�]�&���|��Ǳc�p��Y���*���w��!+c�;w�L��;�v�:+��?�_�����r�J(�^+++C_ߵ����[V���6EŘ��χ�h�j?�`$����S��5횽O<-�'6��8����t��r	y�P�I��������2���O�.���===�qӐ�+������G?�[Ӵ��u���wwwC�4��:\�7��@t���^{�E6���1M�B讪BWm-��*1����O]nz��\�������qwu���YT�<���n�1aY�d������kC4�/�����7�Fq�ݝ���XVV��w�{�瞻=�J�@��ג�$8��k�"�����|(((0<,�li�wf���0�jk�U[��_LݸN��)W��`4�3i������/�S�0���-̦����Zn��c����&RB�on߾�﬎+�l۶��O~�;���^��~��a��~r:�S�����JK1� Ϥ�͘Ut!0XT��˵��uu����TZ�2-��?s%w�8y�Nq�;�]B�p6-�����u�5�ŋ�駟�������}?��L��v����?{�g�B�g�_������nGhWTT��c,q����YV�^g��`&��������Y��p����?�;0���gQz�,��G��,,�L��8�`�a�����`l��Յ�I/'��;::bVƔM.�۹k׮�?J}`` �F[[���̓��b!��N��p�;�
qM���J���EW����^3�q6W�!�HAӆ�y	^��ҳ�P~�$�Μ���,��q���>3�e��o��o��'��ر#�s��ǋ��� ����ٳg���yePVVfhp���Ų2�?oSTLfb����]��D ��[p�m	.�[[�	���a4<���K�����d ���7�k�"���.�)��u��\�x�ziJ��:;;_�:�l��϶뺾@^�k���X�f����gΜ!7�۽����e�JJp���[[1
Y��X�Q|�<}��Ç��c,����8W_w�Z �-��bSD�9r�N�:E���zggg�.k#�^�w�.K&�o0�v�����u���65�I&''��_�Ұ����h�-��bn�[^��mm��u��n�H�Pr�:��O>�7��f��MMx�ˏ�W�^-��g�MLL���F<�^������v��� �C���F�S��СC8���ꛘ�7���@I�l����@������6�[9�E��Ѝ������|��
��/Û��oX_�~������;＃$ݼ�����]n?�7ݳ�>�C]׿G��x�bTVVZҼؿ?z{��l(84�ǟ~���1[$<�ilı%m誫3���'o,��#G���!��>��f3�������?4{�/�o��ۗ�����?�����#��;�5!V�^�p8lGh�*�c�޽H��W��}k~���b2S�}n�N��`Lv)E���f�w痰o�&�]���"�eq�=UU�t�J�ilD��A��>x�,�ɩ�&�lj2�777�7�){Nq��)�9s�zI�u�������꘲�/�нe˖w |i���b1$	��<���8}:}N$A�����ݴ�P��Z��6m[o���J$�n�cyy8�%t��    IDATЀ�׬ƥ�Rx	���C��,�	�^/�m�=��_UU���B���ǥK�L'�
!vvtt�g�C�j{��}����R��
!�9)�H$0::��+L=.]�����k֓>/0-|3�qc���x����~|�~=z+ʿ�f%!0���3���x�j�35���[�Om؀���k�|>����;3���>�8ݰyV��;;;;MG���/��Ɩ-[
 �M������șí]�J����k֒���S��;4dST�m&�~|�b�m��~;������-�ssq���׬Aoy9�T�:7�1���6��j�z4]2������ӗB�����01͞={^���j ,K����hT��D]�ñ�99Xp��c|ށY�BM5�v+~�e���b8�Ӵ�LHz<�/)��%Kpt�RL������dl^�}>���>��MNNb��������\�x�w�q�������=��?�R�/	!��_���CEET� 'SU���K�Qb� ���MQ1�q�;c�(��8�ڊ׾�>[ގ! ̌�B8W_�OW��D0�hSSv��\�u�1P|�&l ���988����������V��/��©͛7B|���uhhyyy�6E7?TUE__��ȭ+*��1v������m�����zLf�gJW����8��O2�H�Eހe�:�Ѐ㭭�uY㙙�����oV����guLN�gϞ�-[���� ����(����L&WP��Bh��x�	��e�H8���ފ7z��j�pb�LtE�@4����p��	��)D.]�܅�+]��t��`jyy9���-2:z��ٕ���T궧�z��19��U�^	�� Z�_���Gyy��7_�~?Μ9c�_c�8��,���qh�Z���#8��h��x3Ѕ�Pa!N���x[ ���"�j�,�TU�ۼ	���Y���}��'�g����~kGG��c�v���|�E]�� ������@yy9�K���Oޚ��G�]�����C��[�WR���3�_�@��COu>Y���ː�ׇ���a19�Ѐ�]�G4��wTU}��~�����4{���w�}��(�# �9řH$066���2���?�Ἐߏ��>�I,��Ty�0�a	���\��׮��/5MC0D0D ��녪�W�O�T*�D"q�����166���1�n�JlO<��bɾ���l��B�o��o0\�^]]���f����d���3{�;::�fuLN�k׮?`h��47n���)���ԩS8r��5kJ*�o��ὁ�x�(#aذ����J����#\�WTU����な�H�RH&�W�/�]�U��ǑH$���3wpK���E~���onڄ�V,�f������o�' ����{���'_***ڸu�V>);�]�v�6����.��ڵk���gCT7g||��կ�w��g����17,*�q���05i6BC�(ʌ�����ռell���.����ڇ�C��ѝ͋K�e�ٷ�mX_�|9�ѨY����ON��u]����_���I��/�"7���1����R,]�Ԇ�2������HO�����X^>ܰG�.�������k��E��i�x<P��_��LMM]������P�%84��＋�����M��]uux���׬Y�p8lCD�����G}D��pgGG���(�w�.J�Rt]�L����/�#����oe������+�"b�'��p`���������z5o	���Wk-��BQ�R)�������FGG1>>���	�s���:j���7�DaڍM�͇77o�g�ۯY�u���ѣ8I��u�����O\���g�m�u} õx�/Fe�!�q���)�ݻ��=���E]�c�eǱ;�$rf�B�}�=�C!&"� �����O�%�I��������� �i�x�*]�+�x-� ��cl�����H�{��	���㪪n�:'�x����a�z<Ǒ#G�vy�,�i5)E�������/06I��_��֯��W!����|%??��'�MNN^�U̾'�1�͛�骕X���(=s�b`l6��kEEE6Db���ϛ5��7�Ϯ��㧻v�����뺎Çc�ڵYr�����i511q��ٺznpg�zq����x�����]Q��a"� //�'����cpp}}}���7ܸD*,�>�OV�Ć�_B�y��2�l}�aMQD"�O�C�u|��f�����g��O����?�������*���nTTT8>�F�����b��B<��eTJQph�|x�-�k��_�Y���PTT�������Y000�K�.ru�X~>��{�X�/���ӧo*�fC�Y4MC~~��X'�L��>3{y'7��n۶m�v��� �D�-y]]]���t�����"C���S>>b7Pž�6�Bu�u���w�����b�.t]�����}������	��M�p�q!����^��?l���3�9�Y�266F�$@O�RO<��S��>��۷x�g����׎=���b��6z�^���bxx���s�u���2N���y;��1���㍇���n�T��@�Ann.jkk��ڊ��:D�Q�B!x2pݓ�((,,Dee%jjj
��N �I�����z�Y��=��x�ioǅ��k�TUEss���nll�^��R�M�,ɑ��ݛڴiӫB�o!m�udd�H~���o;���CWW����M���1��b28[_���Wq��i�ɧBc�hmmEUU���Z&��=rssQ\\���TTT@�4�b1�����D0��K�`� ��s]�f��݈�hn�`X���C(K���o�x �!���ѱφ�i��Ϳ ���w,���s�&���8����Y�����pV�>�f��ᕯ~���rDQ��������T������d���i���EII	,X���2h�����Y7`�ssqd�RL�B(>{���2��/݁���@"��tS�ҝ8q===�K�z<�o�ٳ��v\��^z��-[�ܟ�������wo:�׋��ͺB���
�?��م���խ8��:��xB]��TWW#�\��~���Y����:�������u�X �cK�`(R��s�M�9f6?޹�n����b�����5�;���>ú��?���ݶw�^���:��������;�_Bee��s�ǃ�g��ԅ@��_2��a�FĽ^|p����\��Ɯ�TUU����-BII	���]硾�!�������������pBLLL 5�0F!�[^�cK� 0>���ޛ���t�"|�=��>����tvv���x���_|����_���eR����Pr�ed�+�����C�;�@��LYq�;cpt�R�򵯢��x�?��xP]]���444 g��}6�� 77��娬������������.[��?�N�U�,���zF��QQQaSD���a@��?xꩧ������_ڼy�i!ė�_v��k���1É�)�����l�⚆7�܏_�u�f9
�P__���6TTT 
Yr�H�4D"TWW�����`ll��!�WR��˖"<��E~�q'��qv�SQ�hii���zNq��Qrz��������?��c���S<��> O ��Kupp��wu�µӨ^/�>����o�`l&1�{~�o��Yn����CCCZ[[Q^^�`0h�s���E$AMM���Fg�<m�5r�yi���*�ix��{�?�����͒N311��R�	� �ھ};?��/�����߿@���x<UUQPP`Sd7��񠧧Si��ީ�����Iz<x��{���{1��g�~?������RPP���j_����,6P\�#���BA/7��̚��ޗ�dX_�`����ddd�1�� ��~���'����U���B�; \3Akjj
^�ב���|8w�aЄtU�nSTL&+*��o|gg" �@YY�����Ԅ��"�f��d��@ %%%���A0D,Cl�	�	��-BOe*N��6�ÐX�li�����Ο?o<���TU���|�]�@�����J5�QUUtuu]��RUT�<�P�p$�n7�3v�^/~u��8p�-3N��4���X�d	���-y 0��x�5�~?���̧w��8W_���'Ỏ��)E����k��TUUI�	���M^�$�8t����޻w/?�ы/�xx������e:55��#տ�T*e�H��A���<����@q/}��8_[;����Css3���2r5�����A4�:ugddĴ�=�i8�҂�?��S��D8˘�W��@ɵX��0���m��Z###8|�0�R�����⋳�wϮ��/to޼�H�f�z*�B"�@�,�����#s��(Jk|gl.z����7���U3O���W'����ٚ���~_=�=::j��$�^|~y�k�3<P�ݰ��*]�԰�h�"[k���СC�a]������m����wE��k�0]��©�g�^/Z�{Ϧ���#����p����9,
���	�/FAA�%Î��|>D�QTUUAQ����6�'=�ln�x0��S���4=��9誫ŉ��zss�����6������|݆�m�޽��-[�� �<�����M�###I�]]W48`SDL
B��ڵ���È��X�(
***�l�2TVV"�6X�� ���JD"LNN�M� ����6D���78ha�Lf�^��b�����$���O��R�'�|��|g����ۼy�y!�c�;�ƙ�|>N�>mx����Giڭ4�݌�����KJ�'���K�L����hllĭ�ފ�����B���6l��%K���c�g{�����N7-�0B&���R$�σ��BQ>�'*躮w�Ν3�a�L���	�p���ɓ�×c���B�����t��/�?}��,*2�3�P+V���u�PRR�U�^�������PWW7ㄳëV�_~�71R �Af���*ÚL�fs��q�9S����SO�d��L&�=����]]]w��s��CN���\�� !ph��/~�g�����ŪU��f�D�Q�]NN���p뭷����4�҅��7��o~㹹�al6=U�\E�4�ɞndd��D�c�d�?[�,������ד�$N�<iCD�C��#��s���筋�O|}���������6l@YYYV�Y4MCCCn��6����Xg�l�r��o��"#d2�r��?�������a����h4���xd�}����Y�z"�0�@��>i_Iɬ7�1ff2�+_݊_�u'R&��BTUU��[o��ŋ�n�p$�Z��>?
��o|�o����0�u{����9s�p� !���'�|ۆ������?�������:���^��="�a����8�Ѐ������+�)%%%ظq#jkk�z���+�6l؀��Z�bk����{mXoq�LF=�À��R]C���cv=����x��xd��OB�I���Ԕ�
$'���!�H�4Ʈ�.޾��y��H��!W�_�E34�gMӰp�B�_��3�_����O��6.^���؍���(q��[�GGG��1]�������!Icǎ� ~����#Ȩ�>մ��lR��7؂w���<�ǃ��f�[��,o��z�hjjºu�f��议�Ϟ�6���Q�9�E��0???�)3�����z*�ھc��{�٬��8����ՅI��i�|��؍��������6*����zlذ!�og�x<hhh�ƍg�	�������6.��+��E�:�����(OnݺU�i=6�u�����Ϝ9c~s�P�	]Qp��̆h�Ӎ��~��p��������b���hii������0֬Y���V������-��c�"��=:,����bL�=�d2I��
�/�L����HGQ�� N8qh&���'������9:��?��r�4�EC�+�l�2GM�x<hllĆ̓2!��w�����?F�&PM/�m8q�Z��u��:)��G .���<y��6�T�7��Y�T{~�W�2�3EEE�n�F�`+W��ҥKM��~?^��7p�����L̦�T��ɉ'��S!��w�����ߤ�����n������9�7���橨lN~�/�ؒ%������jG�.���W7_͆��Bx�~�]o��nr��̹��< ���SO�b��ٱcG,�J����T*��I�>����6����͛q`��?SPP�6�����a�l�����gy�^���|>������"��ݸ�ǃK��2�.���f�����'�|��xd���9�������H$p��;BʈP(Dֽ{�y��Q_I��o����^���lTQQ�[n�3::�h^���1��M�,{]4yft��e&]]]��v ��o�y۶m�L����ׇ����[�D}&b~����36W����Z�{x����h4�)�3	�X�z5jkkM���kVc�C���ͦ��4 ����K�0<<lX�u�/:;;�mI:۶m������I�;g��X�u������L�5�l݊�/&_B`ѢEX�bE�]39���X�~��oG\���[q����Ș,zˍ������)6�011��nc�"�x����B�����W�Z*�r�����^�I�]�XN^���qf�B�uEQ��҂e˖9�;����֭Cnn.���c��Lc�ő1��D#>�]�=�����Xd�����B�C���Ν3��v�s�SP��J�*^}�Q|���|]���z�Z�
�@���2����֭3�Iz<��c��H�2�#c��/)!oj�i_(���������Xd����0RN�>�dҹ���KD��13jj�·~� �z0Ě5kPSS�!�i����V,Y���p��*���o� vC�=�@ `z(�if�Q�WU��ju<�J&�b��I��H�p��-��$�b�:}�~޽�N�!�|�r�i�Nr=�=��.�k�>
��,�M�|��3��W<9��d�����c�c�Y"�x�a��'���>IU�PQ�Ѱl��x����\}�zNNV�^�X�<���cv(/�(����8��fqdL��%�5�7]�;}�47�Y���c����]]]�ڄ��|��e}��6DÜ&���o|�t�n ��5kP%ɔ�@ ��kע�d�^���/��Ns�;��ѨaM!Ume���I\�p�z�5>��9BDΗH$p��Y"��s1P\��e�Y���ʗq���\����b�
4448�9l����Z�
uuu���(�����l�r�cN�_l�]TU5= �tcccf�9�����S��նm�� ����x<���."�*w�:�^j����_3�\^^^>�|�)++�񿧿�/|�70���������L5���nLNNR/��˃Y�ر��/��188hGH��*B�A���]X�pg*c���ex�;��TUŊ+f�x�T�h�֭3�<r�i޺�^��bN�WBo QI�MNN���xc����m�6�ދ��v��1����ccc�!����R�صtE�k�<��tX^^�#���͕CyK�.�7����؂��������.K�&���5���}��׬�GfB]�u�����ǎ�n����%�MRU�|�L&�D"�]�y��h'S���hii!s�����GA7_?�f�_j�U�~���:����&�	!7���SXX�� ����?ކh2��U�|>�JԜ�����zB(�ڵkQX(�
!.\�e˖A��	���״�13T�%
Iq8�2����27H$?`�fwr�B헎��!��Y�5�KJ��[��x�����&�s㕉�Q� 8 E"�ׯ}q�ȬG,�i���wr8��:�]��'����\%��P�D�Q����,�,\�77o"r5M�ʕ+�+bN����f��M��V,���n�8*�dDc������u�.��������HOU����I���� ?�����6��"zs1�`ժU�\�G)--�ʕ+�!
�)E��_~�t:,c�&��V���fz{{15e�Y�?�:7�F���� �Ӧ�Q�.^���B`�C���V���bin�3SUU�e˖���	��|u+��<�    IDAT��& Ʈ��ge@1y����e�֭[����Y�����c���}68_a3y��/���F���|�^����H���X�j��}1d�t��72F nʓ5w�u�,w��������nǎ1 �f���!������3�D-�8�$#���v!/^,���+TUE{{;*++��/����[���d��l~L�� �Y��b�9��O����9��?�utt� �O�����H�R6D�y��ɡ#�n7�36��x�G�"&U\�ZZ�I��׋իW#�����|־�⨘S�>�d��۷o���X�`۶m��/���4p"򁀧��i��z������bŊd�lfj�Ox<��֯`����Ș�P�
 W�b�$�����cu,n�u��$��I_0�4+QM	��Kܜ�n�;wߍ�--�k��߲���O�iS>���a��=��P��d����������u]7\��2�����X��I���4M��h��>G���5kph�Z򵢢"��oل�a�Z�����T�>�(�i�]!�z�����3=�.�G� bN�]�~?��8PRjC4�	b~?^���'jt��bٲe���2����|M~�e��Q1'2�#��p������(8W�?�O�B<Goo��d�:
�E���Θ��ߏW}	����a�ʕ�L����b����o�{/�J����n��0 �����0��
௭��MR�����c��'u�/���Á��ע�(�,YB_)-���<�X��l������c��6+*W1k��I<�ŋ뺮������	BrUUy���ڄ�������3v�N�����U�keeeX�x1q���"�����|m<��?�E��>qM�h~�a]��J:�	�	 ���P\�w~�w�u]1}����|���멪�{w~�|��� ���8�wEnn.V�\I6�O�|x��G�pA�?�9�bDM�e��xNN�?X�[l߾����34�e�`�x��@�YA����
�X�d	�]v��������k��Z����GĜ����4M��L�>���8hu,n���K �+&y�����G�2�wH��_>�c�f�����+���m�^W�ܩ��ǃW{�����醉C�2��0 	!��Z��$�� �������8T!s,/��]���D(�_=� t�	,cɒ%�j�"//˗/'�.����w�eCT�IF򍹊������!*��W6��۶m��{��N�c�� �{3Z �mglnF

��7�����Օ�K$�ҥK���5�8p}����h8 ���R[I���cX�u�����n�q!9L���P~q��1B�����rr����5���\�Ci��B���D������sjO���N�����|�'��H,3t]7�.fC�����5K��Z�3���k---�kn��������k��s7nd3o��%o1�mB�>�<ڶm[�ߥ�_�t	�d҆�2+''�<>�7��q_%���ph�j�&EA{{;9��-4MÊ+�Ӊ�xk�&�bN�TU�Y��l��|�����Pr�;v� ���u�n����*S��qI�pe�GW���#*3m<�E$A[[�(vx�
�nZdCT�)F��F74���n�|��'�Y����7�kCCCH$v�3gB���7^�4IUū�>B����wm�����hii!_;�a�/X`m@,�Q�� Hy����&&��!��,����^0��>00`C47��=RM�ń�=Hސ����b�
r��[��a�:ˑe��y[�Q1�%�,��H����� ��9w��'�O�������ͣj���g��[oy���3.Dee��e���VӃ�^{�!�]�۱�Q{D���芢���y�J��`*��ࠡ��HT�2���,,3ܻsĘ��h��A����z'������e��b�筋q|I�Q1'��''��@�L&͒�W��ōt]�y���F�Ә}>�yҘ�\�j�W,z<����z�����R���_�|��K:�ݼQb����l.]�dX�u�!�3�rvUUy���j ���8Wa����nå�2ú��E{{;9��m*++�+�uE�އBL� vc��G^�W��f����ju,n�u��) {�ם�$F����s�ņ˗���uUU���.e#�\����|��M�����q�H�:�I�2566�K�cq����I_w� $*w�ɛ��;%<���#H����R����UvB`�ҥ�o�PQ޹�o�a4�/Y� �<�ܶm��cq�����6}������k͆t06W����tB����#��,--u�)������hr�ջwމ���؈�U�23��d��kV��F��� ���ԍ��4M��t2�<1�����Í��ZZZ�)�dBCCy81���ݻ�!"���+��$���I�Ca�[�=�䓟 8����&��ι
��`4�Ckא�-^��ƦY�h򈛚�C!|p���Ĳ5�H�g ���C���wz��ō��\�I��LG~F���+�D0��M~g-Z��}���֢��Ȱ�z����$�hT�"Þ�$wy�?���ձ��!w�a�.�Q���ǃ�y?����c�8�����x�b"�N��a�ҥ&��,E��0��{DT�"��~lݺ5	���u'�̈́>�Ǉ�Yfp�;c�]�����A��`��'�A�xe�Q���i�S�L���۷�:7zꩧ� L_�偀ڈ���w�=�ՉUUU(#&���K�,!'�޺�,�>(�զ|>rB��McW�MG�z�{������/8���ʷͰ+��{9H�����)���(X�t)�����-/�!*�md�hMG�RM�l~$�Iä|]�y}���x|]6~}=����UUU6D���hkk#wN76�S��ɘ����ƹ�u���%�LbhhȎpn�Y-r�'�2 ��h�:ú�(X�l������T�"޺3Y�b���0E��p8oll�X̰�J�8W���0����ɤ�d������K��e1��}�����(~��������?moǥrn�cךk�2�����B獆p.�@�Tˉ�����w����T� -ZdCD����T�w߽��̽̾[e�.l�{y���ZG�uC3::�T�pAMV�r�I�U���Z�eyyy��"3��t!��{����7)qme�X,Fn�&�I�x�Hgg�'���A'�ZTU%>OC6DòIwu5����g�%����5}o޾�$x/���j-24��'o9���:����h����]V�z���i�b ��}�!I��644��±/�,P���G��d�
"b�j2D?#�Pw1y�Oz<�_Z�[�R)�>����U�Q��	ɇ�1�p�;c����˵���<yΔ�ih$�tE��w�mCD,�ňϘ,�G�ƌ7L��kBq-!Ļ�k��~2u�h�\GW�s�������M����Wh���m��e+*W��a�pc?EQy����#�9��b~?7�\����w�iXB����ܬg_���D��t�[^��یMx�]&��0�{���~5M��"B]ax����	�w	,���� r���&i��󡨨�������0>^�Ɔ�X6sK�b����4�}�cq�m۶�H_wb�"��k-�/�zgp��ΰ��o��Qss3Y���m�m>̝̞e�#2�=<�m�6�bw����O@�sb����[R����Ę5���1|�$x�}�a����D��PQQA�x����"bيjȕa"j"����$���cq3!���vRc�L���oºΉ�f�����d�6�VKK�Ƀ��!ɇ�eT��lCI&f�M��p�x<~��J��1T����C.wd�R�S�***x��u0;p`�z><�r�W7�o۶�ձ��!'t�ƫف<�^g���G4i����Z�-"�-|�f�4 ��qy���m۶9��^��.T�e�s��p�zr�	�.
�� �|>|�j����D$BHq���k�u���,ty����u�����`����r��(�,Z�H�"�|hjj"�>�e�ѰlEm��3K8���Z���G��םZ����2Ɠ:�E|�~�a���`ѢE6�<~��������\[�Ć�X6��[=�ԛ�d�X̰�y��v��p&}�)y�YNϓ��+�(8�n�a��8f������*��PQN55��
B�����xYC�&1����G�u!���m��yrrr���`X����Y{��l4��!E��܅�����܅��L�]�{���AQ'(++#�2���:�9�^�� ���8W���*ә�q��n7�3כ�������@ ���2"r���\���ֻ, ��;QS�$��)�i�I�cq���� Υ���@@n��iWW9�؈��a����,�1Zmm-���Ѻ�H�ݙ��zo&ccc�uݰNM�`��P�5�V��L�spӘkom�h8lX_�`��߫�T__ONF=�q ������K�2LK��Y��'�I����V�t�kj�SYiX���@0�!"g���&��[����Ml��n��܅�#�{>99�D"aG,7�|Ĺ���Σ�1���A]]�a}���g˗��6�Ğ��,3�zϹ���lp7����3,����ާ+W F����8�g%�a  �]cq$,[MI�Y�4&�z'�m��:C3�7]�Q�$�.PEAMM��8������6���q�'�1 q��U�FL���d4���X�N�uC311aG(sf֜0E|��;P��=9����z����0�����\��f&����V�*G�x��4�|ϩ��Y[�\ŵ�_oXB�7�1s��`�����P��Z��e��ɤv�]�|1{ϝ�ODNp���v}.�����SJKK�sRQQA�:�vBb�3����8��$��*K�R�������$|<���<�uf�wt��ZNN���m���rssQ\\lX?�p!O�c ������n�0p��8 �/}���9�)DA%)��4�>CEE�h2U����]MM��s��͆hX�I���V�;X&&y��֭[������<����#� �����l�.VT`0j�y���J�F��V[[K~���,&��I^"c�b�,ϵ�uuu����q��>')�.��x(�s��� vc*++���ҥ6DòMR����8�NUU2wqJ}e:�90)��*�1G��5 >�7wfã�C!t�td��~�ι���J*�"oZv:w�/�g��E��.VT`��аn�y�fG=D�'x**]x���i��7bu �����R��\�X�q�O�q����c��j1
��&)����LL~'9�������I�t��s��K���̦{�ٙa8��ȷ:�P��U z�����d�k�Ν	 ���N����x�Օ���A'�=p���x<򶼞�
���6DĲ	5H �3w���9w�^,#�sYr��3��RU�hi1�G�Q�������;N��1wI[d�[��k�ƹ��TU�&WIG�]8wa7��w�ըMW!���l�F�p!�9���d���dx �
�B~��p������>&!p�u�a9������*���)E��>��v�a<r���4Psc*tRC�8���6lnR�Jp�F��r3����0��5����S�dSH�y�o`*����Z���]�SP���Byyy� v�\勚���'ȗ�$	r�&�.�۱cG��VB'�.��`����نL��P���x<����O/jD��!"�-��Y���~��*3; 餽 3�$�����鑱90;�Z\\�Wf�$j��Ŋ
G"6Dò	���P������O͘6��TT靯��(1��ݜ`0���<���V�&7sj:���L�&��!�pt�����K�1�t��������~��̾We�.{:���ͦ\�y'E���$&�g���Ri)��Q�:�*7���#B��ok�(]άW�Z���"�.�q� �+8waWP�������Ȇh�A�KhN56��n�g�����:�SŰ8�Β�� ����oa�nPwe%&��A.d޼��2�)F!p�'��^�Hhd=�*���!�B�����0`�9���;��XHSU���6D#����2�@s]5�*2/gB5��<����'m��SQ�C#Ln��4MC�h$csCի�/X�XN��0��&y����̞��b)j-�A�����a�o���=*,$0���'$[�J��uEQ8w����9Iq��uR����z�zii��u����a'��_W��Yd����3�v��I'1l>��
��d����|q��0c7��o�fFNN�Ds؅��e��tnC$�E=��n|"f�Na)�$;��*�����c��F��wm7��k�=g�č߫f���0�T�<��<���Z�ϊǁ���P������5�؁�]tEA7�.��&�g@�������F�Z�ئ&8Wq���faa!�^����,�;O��1�0��a_h:�ƷT*Ź�=��]���y���by9�fX硍�A�����d�3s�Q�����o�Ν���b�D����d��#�܅�<��b�u�h�.((�M�),,4�uWU��i.G5�:qjB:�d3duH�R��kN,\�3��x��]j�~?����|�df�|>���2�����Ur��p�=���cȦ�x܆H�]F
��M(��dF0D1��sw1�^�a�u:EQ�Oɤ1�g�N�uG�(WP��'����$4++뜫d���A~~�a���[r��$�]lcxߝ�4F�.\gq��EUU�7����2��oQv-j�H����^�F��Cal~��J�N����="6_����RB��K�ƤXvc��pB��[a, 3�����pi�1̉��t��DI&!$��0s�j�M�HĆh�D����jm��eY��3�<&{8��o���5kBX���܅��\�쐳��gyUU���~�
r�q��WOe%9���,�C��jj��T�rK*y8���p�b�ݻwk |��N�]��g8wq��M(�H��6fH8&���.�<��~��%8W�X"� ��d�i�8wa��J=��H�*o�fN^^�0p��چhX��6�$~ ��0���N}N�a@~����~�~?�l�)���x(�a��v-Yo��	�1���y�����.�5��%77q�6�1�`��h&<l�-T�f\���HMg����WB���LǇ�Xwu�aM�4�B�ӑ)�SPKJl��e�4�_�@��'�[O�����<�]�$���H��y�#�@������o�s+Y��̞��~7��QE�w����7�3W,2�4MCn.�vg�ٔ���ѰlA]�+����|%���݉��t�0�NT���*(( '�D9_q+j�H�\e&&E���;w:���<�/~�5�n:0kf`r,4��ƃ2�|?��`���39�=�x��Z�Cwww���)9�t���� �oV`7&�M�č���rk-&{9w�X"� �s'�&s�r���|$�����2����s�ŵ�="j.3�K�?v�Q�-EQ�\��:�]ؼ�w�JCD1���3�zO����ը	�2<�|��!����0[,L_��ɱ#���B�;�
O�,M����A�W\��n��R���w�STTTgu,̹y�YsOs!0Th����%��~?�Tʵ�p�T�7P�hC(��i��;%G��������s��R�f�ab�s�zȱ/���mT�s��R)�=�j��.A��<H�]��!����ȋ�i��E��!f7�{V�����5�mư'���:�ƒ�t�]Xp�;s�A�D���n�p5\X8���q�>���ht�š��O�� �;�d(���hs!SfqM�QT���s���S�A������L̾W��,����)�������� �����v�~5DԹ���d��0��I̤V�Mb�3�'�Ǒ��T��q����`��Y����=9�f5l��.��s�b1�=��|��>�Mb�2@�~���Hqsu6!kWB`�o%t%��-C�"� s��^*�r�>�L�ܹ��n7�3W�&�����m��Ԭa����4��%(�pcXv]"����}jjʰ杊�	�ʐɁ0�=g���7^��K�*SSSROqWU���p#    IDATl��1�я~�P���f9�6i�L19Qu�s�����χ�3�ә|p~b=�{��$��h\[q���|$�f0�U2�lp'��3w���P�fs��G�]�'M�B}N�)�全�G���%�� �ǵw�y���,YC�w����c26W���\'��`��q��#ۘ��|�սB�Æ�I	�^<7�e��c��av�ib1�k`dĆH�UF��J!�~��ȍ�W����Cp��ݪ뺔��Q��F�Z^������)ϩTN/R)���l���a� lX�4^��9�I��a����$j+�3�ә�<���V��r�4�Q�J������L����9��u�U�JI��5�˰/��$w��|�,�5x�)��tT��}!W)06�s�yf{�Ü��R`�Xs�e���=B�>�Ũ�ܩ��tf�=���L�w�:S9>r"�Is*�	����]��^���Ȳ	k�t��:7K�R+��rrr�(�Ow��?Hm����z���*�9T���3w�� 97^���]���l�$�I���z�g�?6FN�cr��{6��2?4M3�M�pό�P�&&&l�d~�p[�(�2Զ����:�V\.N<���
��cC4r�r���!%A�����"c����Q��b�V��V�?��
`Y��s�d2I�>0�]29M�S��2?��5NԺ��̞e�i1�jz�g��4ؼx��䥯;eh&T~�ŠI��a��js���N���9?��5��	nn$N�NLLHq�S^�!�;t]�nT�!������oG(GNp'>OLS��+�*�z_t�xu%��8ِ+C�r&�����ҧ�~��a����A��a�{V�1�������i��O�wjj��Mb999�a�T*u����O?ݨ�ze��I,��])�Mb�'�q�2?��W�s��K&��B!�ΘL&��l~���.`������3µw�}"�P����S���r�} Mq�ձ���(��P��\%y�ߚ�2��6��Ѹ�9?��uJ���
����S�����l׮]MV��F�w��1U,1^��D�4�>	bZ�*�,�8�<��'R)����2/gRXH��+B�۬���nO_pRC}F�nD`r�nj�M��An�z��m�LN2ߎ��䷐�-����kB�XV3m�|�5��x�������u1w�[d�]����B�n}4�(�!wQU���%ۙ�.\kq�0;���iaW(�r$�#���%	p�b)C�{^^�Ϧ��\sa����u��B&����BOp�B�[�^dx (,,� 
�i�,���m �'5����bH'�yʘ���j�,�ҹ����� �~?�7�Y��[�&}���AV"�s�m3�'6�x�u~P�.�+���r���v�e���r���<�&�lG�*"������D5(q�e~���f{sL~T�j����~�Ɵ����k$X�Q�K8����:����A��p3G�Qp�e~P�8<�ݽ�!s��]�\%�Jq?�t]p����P��ga��l����4)�;���	����ƅc��BHz�������7�!�!7�+}���!�KF�M��	�r��8W���Ÿ�ݵ�/gBф����$�IC���Ts5a��+A�Zx�u~p�#�͡x<�d2iC4��d�OB�!�y�s�N�ÎN�x��y��8y�<�S�h��:��0�<յ�:�����ɜ���V��6?��� 6��;5w�>#�$�>	���k-���������Y���AB��ݻw���<��3� ���N�UґC��&c7��7�ut�pj�5s/%��|ܰ>N�9�|�~�O~�9��,�s�N���[�ם4�t&��C�:��4����Ƶ���e�,6�I���[iu,n#�x<}-77�1�Qu]'�|�1�q���a<@�|% '�x�u�cq����{ 6����J}>�n�d��ޛs/��s*������!�.����= ����܅��:��7�������s���.2�� P���W���m�|�i��fB}F�j���7�3��T~_�amD�Ħ���Z�MMM��Y攖��#�(I_�F`i��.;wp���1��<1�Ut]�vQQY�O&��aC8��k׮: �In&yeV%?�g�1����� oǓ�����MB����O�q�=K�R)C�i�c�Ć�f��K��0Ƙ����us!���P�_޽{����e���|>��e'�>�}�g�1�XfQum����A�oY��<���*��^XX(���͒���L�w�c�*�hX�x�(??�쁀��Q*�2<py<iܩM�"a�1w�߱�dRʩ��y�^�S���ݻ�1J܁t]� �ɂ��r��1Ԧ��J!��kC4�1&?O"A6���$ eeeԲW����ɏ~��< �����BQ���D}>���c����"0:fX�5w1y��K$Y�[����y	�������9�Z�urߔs��F�Ec?�L{D&���ݻw7Y�[�����Pન��!�̣�Y���~+c7�H�c�E%1��xL�=��s���v�ޝ���w��q_��g
ڠ���b��bUw;�]g�8v\r7��or��^�nVY���� ���b*V�z#%Q"	��D!  0�e ����?H0��΀E��7���y��y�3��'�3��}��t-,,��kW@}П�x(BDD�#kxP�K�4��,7~��\⁔R!~7<�j�*$''���MQ�U2GF`Wt� "��:[�j�Xff�������V��n�� t]f#�������.��(Z "��O{���l$&&��ܻ��@ � ��Xݻ��� ��ؔ5�"1""#�R�Ye�����դ+5lT��H��@���	ِ�������<
�B�����LH)��ѹăP(�� t`�zp.`nnN�4!"�����G���.n��˥������7kB��	�X����5 k�㱶�Q>��+�JRu��^%�ߍ����ۍ���.=�ӝa���`ժUf���E���NbDD��V�Z���"����������.M�vx<--iii&d��E��7�IyDDFH��G���.n��KRRR�������;�G�v�K�Fx<??��y�Bˇ�DDd�U�ð):X�"699YYY�������b�Z)���եH)uw���1{�.��U1-�lŤ�<�[��fC~~�j�^�-?���_1���MS���he��z���caa��lV^��bB���y��/ ����ɕTg+)��H��5!"���j|4;;͢��"L���B��1:��4�w ���#�oT�,�##p�&dCD�T��V�#���dNJJʟ���	!����xqq�	٬չK6�h�����e�12��[�� ���T�$MӾct.V�
 /<�z�j�Y���Ĺ9�&��Ɖ�h�����p�W�f��n�' ��)��G���y]���VV�K"��W���#�m������|�LJ�|�WZZjF:�By���xDD�R��H)133cB6+/---R���x<�F�cU���v �G�#���T�<g!"2��'� !AWs!�_�۷/ф�,�?�A>�?����[�ac ����Źw���w""2��0s�B�yyyp��ӛ����l��}��%�l���'$$���Č�V;��Cu����-��J���, 3��{�f�s�"��_!"ZY)SSHRt����J���*UX���q�ݟB�
�#))Ɍ����lE5����VN�ovE��8ܻ8 ����X����o X/--���W�R*_d򜅈�H�C�?w�tGd��Q^^�Z*r:����l�+~@rx<��:sxGDˋ�DDd�E����	ˌ�B��Rل#UQcp:��t:�\J��d///��n7#�1:��v�30`B&DD�%ҟ��?��(R��f�g�s�"����Rʏ�����bFJ7mddDsMN"٢]������l��{���t��䨖�X[[���|�����!����x,>�����Ǭ�1H6�V��e���x\d�Kvv6222TK_�z�����j~��'	!�_�`/&LMM)'���DD�rr��Zi�RVV�|&���}�������<���R�o��SSS���oFJ+B�{"��Gڸu���X�NDD�+<wN�B7!���@I��׻Ǆ�,��v�J)�6<�p8bzdv�����������?DD��\��H��UżV��LJy����-R����� ��c�xLuxY�����+P�y;66�P(dB6ƈ�w�MJYWSS�0:+����3 [��EEEHN�5�����(��1>"�8Wt�[����d��SJ�R
����ٿ���PRR���2Z�s��!��τl���kbic��+���v�����
�?������A���BXg�ڻ��,��'������=8�D�_�ҋ�%��ۤ��������$��������a��l�d[(���^�!"�?ŊEVګ\˚5k�q)�C��q�����U� 55Մ�n������u�n�!"�CŊ?oC�&&��!)++YYY���rKnn�7MH��^o1����g[1C��B���;����n],(�WZE^^�ӕG(wz<��7:�����B�Ux��p�d�+��.�}��Ttu'"��U�ػX�h����.� ��v�o1:�ؿ� |><�r�PXXhBF+#*�!��w�>
��ᄔ_텱����"dff����������X����,�_�'''���IU�{�� ]݉�h�uu�b������3!�edd���H�Th�������ڍB����v;֭[gFJI��;/����38�D��C��gB6�ٸq��ӕ�~�a�慖
��///WN'�%��J1������6M�ŭ�	U���:���A�ǳʄ�b��iH
�WVV"11ф����R���,DD�P�s[���tb�ڵ�% �6޸|�e���E�i_���ƔӘxGDˍ�)��I�&d�2�/^����6:�X��z� �@�V]]��:�)%���tq�Kq""Z���)G�Y���J6lPv�B|���~҄�b֏��P(�( ݜ�5k� )Iw/�T��飣pMN��Q��
g+Vk��rEz��n�������RLs�ݿ-��Rx<)))滷���`^����f��L���_���%33%%%��< ?�RZ��� �� >w�\X�z�	-���	h�G ,#"2Gaww\����(�6
!����}ׄ�b���r�mJ


���mBF+G��O��F��~����S	FDD1E�5Rw�X������RՒK��z(��bQMM�MJ� �̦��|��暐�ʙ��B@1r����DD�I��A�����*KY�{�MJ�SvI�~~��� ������b�V�!��{""C��]"�XIeee��a���������*��]-���H��p�ҲR�B!��J�1T��GGG���d�ڵ� >W[[�m��U�������6n��M�Tg�΅�����ʋ�;"!�R��k<��F���n���q�ݎ6��
S��vu+�}���'"�����!ezZ��(�k�F�xݚ���ODW����� �[�ˀ���=D~_�	��/U�������JJJ����Z�c����v�����ט��fff���u�bE'a""Z9��X�l�J����xRʿs����R̩��KB�p�����!//τ�����.�30�EWw""2�j�i�r���8�N�_�^�&�������N)��۷/�f��@b�Zaa!���L�jy�b�}�Y��*Q4��;����HM� �z��H��jkk7
!���֮]��D�&����ajjJ����i�:���.\���Á-[�(����_����"p�ݟ�R��jm�ƍ�Ĵ��]����`Єl�����uaa�r:�"��֭[#u����}��b����7	!�U�VQQ��u1!%
86���P�|#���?��&//%%%�%��1�ۭ��%@J)4M��9|-11�6m2!����Ċ�W!"2U^?���F�w)..F~~�j)1
�b߾}�S��jjjl��� �	_KNN���1����abbB/T�M�q��hݺuHMMU-I)���S��!����~f(z�&999(++3!��i���=C�Q�����LSq�M�����,TVV*ׄ�Z[[��S�	�����O�������Ȅ�V���4�
�[ZMȆ�(�wu);<����RRR�*t�+����F�+���Wb��~ =|-++k���ec��1^O/�ggMȆ�(�I��6�����0�q�@���iii��B!��0�V[[�? �~x\�-[� !!������࠲�F9�V��Le�4��=��[��ʦM�����Z�����я~���Ļ���� |1<�ؔ���z�Hg���>'���v;�m��]9���P(����֙�y衇���1|-!!�7o��)�ע�=�30�TŃ=�����iJ�v�� ���Bvv�j�
���z�w�S4s��k4M{��pjj�%�r��
�D��""ZY�`�g�u�x�x�RAAA�.�B�/�������ߟ�p8^�k͑����[������4ffft��f�!"���]L�4�|>�1��f[��u���y�ۭl?�<�7���Z[��*�\�pAKC�E���bIe�~�b��G�N'n���y�b����3���K4!����z�NJ���֭[���©�r��>6fB6DD�(����R�v~~��������III� �+|m�!^b���v�����3�3J���w""2M�/CCC��Bp�NX�R�gkkku/;���-B�*����t8��["]`�<�%laO�r�<��*��k ����pKtI ����~�������N��l/Н/�c�PS�/B��� ��E�wK+r�\ظ1�Q� ������������� �etvvv�Ƀ�&R�dU�E�xk|.==6l��|��������ּ��A��O����Z���Cyy����ߏ��I]�Bq&IDDƋ�;���b)פ���x<cpJQIJ)|>_-Sf k5�<s�R���h9�����L��B`�n���صkW���١P����輢��㩔R��"|M�m۶��r������Q+��LȆ�� ��#�/^�d�ٰcǎH����y��/�W4����U ���7l؀��c�ZfCCC�XQO�����BJT��������4̈́��WTT���*��3>��}����VT�x<_�c\|�x���Tl۶-f�˄��I�g+DD���,�:�����a��Ց�kdd䩇zHy�/�^��B�wIOO�֭[�Oj�(�Y$FD5��h���K�c�7���?���8D�	555���C �Z_��
T?�yH7!�,p'""S�������.����k����] > �F�~�/S1O�so����Q���b�4���������JIIIعsg��z	R��=�׍�+x��򅅅CB������*����ֲ���´����'��̥��i���M��k֬AIII���������52�h�v�k � G�Zrr�R{���:[����G������p7`ddĄḻ~�z(פ�_HJJ�U]]]��i�NJ)�^�?I)��Z�˅�;wZj¯jR^^?RY$FD��h��`zz�^U[[[�Sg|�AW^^��B�?T����b���F�e���Y����
b�;�*�����A22Fvv6�n����%�|�����v�?
����p^�~}�qXV �����u���n$�Κ�-�t���q�h�u��5������v���} �T륥�X�F�~/�����b��;�q�{{�25����ܶ��7"???��n�����?��gU�:�y��ZOHH�Ν;���dtj+fvvccc��j�$�'R�#���U	!�u�VdggG��=���]WWWhd^f���O�z�?�R��j}��BBB�ѩ����IL)��M�&dCDD�������Ν;����\�R~���=OSg��ۗ�r�� �)�zff��&�(��<C+��DDd��f�A��i���7!�`�ƍ��At    IDAT6�N ������ۗhpj�����y<��[�+ ���TUU������v���+���ڕ��t%��H����{{{M�&:ddd��[n��1K��^������Y�f8���G�P�} �K���BTWW���?/��c<""�	)Q٢l422���22�u�����������y�a߾}%yyyoPN�q:�عs'\.�������^e�J��E��a�u'T��U	!�}�vddDl�~K0<��x02/3x��r��w����c�$'[�����G,#"�:�zG����]�v-�0�ד��?t�ݱr��.����V�zZZv��a�)3�B����F~_\&dD��DDd���N���_ ���[�l���S�-���^]]]����?�A~~~�� �;��_��O�Eu��8?���&�!"�+�4kO���GGG�]��ENNv�����#����p���v��y��v�z<�G�?�lcRVV��^/����+',Uk4!""
�>Ǫ�Vf�ٰs�ND��*���K������z���Bmm�g�1 w�֓���gϞ�F��$MӔ��
zz�9<lBFDD�����t1)e\�]�n�c������Q�!���v�����ޒS^����R6أZOII���ފ��4�3[Y�@ ����x�ٳp��y#Q4��;���d�z�HMU�)��r���������R���xSJY��LVV��ٳ�]�%baaA�>���-'���l��r�3==���Q22Vaa�^s��4���vYJ��Q�x�����R��U닝׬޹��������I82""�p���d������Ğ={��q�LY(z���|����2�{��6!�Q ��3k֬Auu�%���Ϻkr�g�MȆ��­����9]��������y����"~���|����n40������n�?�B� (��RSS����e(�P6m0!""����^d]������)�qX��nǎ;PTT�#6!���|�7���G?�Q����/�|
�*�g��Ұg���(�
Ĵ���+���5!""��x�#Z|(����#.!�O<�O�4�w�������^�= �g


�s�N8�eKQ=DM��EES�	�P<a�;E��ǎî8ȉ�/����w�FBB��a�B��x�޷��߿��ܖ����W{��g���P�T[<�-,,48;s(��H�jdE���Q�tu��ʮ��$55��v\.W��8|OӴ�^���2[~�����z��
�= �U�B`ӦM���̝3FGG1==��W76�
���l<�����oB6�B���k׮]�c�C��q���O>�`čL,�x<��r����.��,>L\b�xLS�!�LO���Մl���z�
y���qAQ�nuBlٲ�Z��4��������1���������V �D���b7�%�*�,)�r�>:��N��#�/�N'v�څ��ܥ>�充�V���Xn�X__���z��f�5�D�ϕ��a�֭�٬_~;99���q]<R��r���0""�	�33(on�Ň��077gBF�����޽{�z�
 w�l�c����G?��y����K�x<ߵ�l�R�/D�\jj*���q$���A���.d��"�X����iZ\��KJJ�m�݆��۵E��oz<�G���b�ۥ1�l��ڤ�_E����D�޽%%�I�1K�ϮiX�	�Q$�ϜA�b4��Qu�������ۗ�R����j�z�_42���v�׸���@Ė�eeeؽ{�e�e���+��o�c<"��Vu�	���x�4>RY�~=�nݺ���$)e���?��x>mdnˡ��n���yM�s [֗��c׮]��:22�߯�o������C����vl߾UUUKM���o^��������������>!��� �#d�v;6m�d�	�עڟ�PՍ�&dC�ƚ���(&mjh@ǖ�W���[�Τ���8ީ��]���8�����?�x<���o|�c�eyc���R4M� �x�����z��[�����J"�Qz�,R��1��ܹs(--����H�mۆ��,���"�.& ~OӴ/z<�J)��7��UwuuuNM�~�� B��E999غu��
�fgg���*�[�<3cBFDD�-Bu�14�����SSSAvv�I��+//{���ɓ'�ݦ.)�R>��zC�������������h�ǳ�'����DJ��6m��#Ęw��9]�
aC�1�!"������	�ڳ����&''���nRf�*,,Dzz:N�8�|�u� ��x<��l��}�k_{I�������d�پ�i�o�x�t:�y�f�����񺻻u1g ���O�]7�]�:�f�dee��ɓ�W<V��!D���y���7��E<� �+�{��\jj*�mۆ��TC���������ᚘ0!#�7��NDDQ#��9��QOO��	�C�u��a�ΝHHHX�Y �@�����n�;�n+����gz<���4����Dq��nǖ-[�y��*n�4My��:>�Ҏ�""�%E�F0;;���2�N������[�r���X2�o!�z<��߿?�^3>��C���뚦���X���ʽ�Պ����R�=��񈈢��c��)Qw��w���d�ٳ���K~NJ�C�T^^�I�������K���v���x~��`�����t�~��/n���R>�+omE���	э�>� ����{�˅�n��z&��
�^�z�^������Qu��v�w���m6�I\|�1���L�~��/n��Ȉ.^u�r�E�����,�~���j�`� �x<��x<w�����������{<� ��k���[o���v����acT�Y aw""�*��;����b�����+n��/�����wމ3g������¢K҅�/<�+B�G�~�����w��WX]]�3~J�� > �Z�&??6l@R�5?j9����W�!8B��(*�?~����B掎�E��둞���{����]]]���@�?��l��x�B<"��7c:MMM�-//�.\,�"�k�����Buu�e4�~?Ο?���� O'""�LϠ��E7!oll,�����_�hnn����R�$�|����n���6��?��?=lT�W��~�~��l����v;֬Y�իW��޴��C���ł��Q�vt�g͚��CCCq�� l66mڄ��B477cf�)jۥ�O�|�A����f��׿�uSځ?���E6��wl6ۗ��[��y�Ӊ5k��M�۳g��Rb�#�'CDD7�wD�.!!�v�B?��ڰ�����?����MJ�����o}�[�qlؿ�&���e)��b�&������q�F����]t���Co�~s�χbE#G���w""�*U�O��;1�j�U���^���_����8�Nlڴ	���hnn^j%p����J)?���4��x�B��p8���W��oe�L<�* w!>�i�B�^ϯKIIAuuu\~ �`0���.]<iv�|�JD��fgQ}�(N��{U|vv���(.��YX�X,�***BKK|>�R �R��_<�RʗB�Л�����a.�|Е��z���~ _��z~]BB֯_�����J-*D*���&dCDD�k�{�s�FH��\Ϟ=��222p�m��������K}<G�-)��nw��I)�)))���̭T�uuu���} >>���)((����㦉@���E�Ρ@qKDD��u��Žˎ;L�(�dee�;�@WW:;;�4�P �;�P�;^����B����ï}�k+6*y����l6�} >�~ �%�6]VTT����������p�ϜA��	э��^QQrss��ގ����7�z!��+��G��sPJ�,�����O��ԬH���GAA�nM���l�AJ��z�)6�����-�-^Dj`���w����!�r`�;E[(���Ł�.����ׯ7)3seffb�޽���EWW��y���+Rʯx<�& o
!>B�-,,���?��%[����ե��u���c'��p�{��z� ��W�^������"  }}}�W�[>� Υ_7�ɶ|�!Zv�Rv�(**���#%%;w���� :::0==}�_���B�/��vx<�n)� ޷�l�6���k_�ڒ��*���	���U6�m���\���*�t^��.���(--Eee%����e1i�@>\�� ���MȈ���W�χ��tl�tU|||>�/n�_I���2��磽����׺��b��B�����{���C��[ NJ)ۜNg���y��<)e5�� �p��iE7��LOOǺu�����*���cp&DD�Q������Y��cbb&e=����Daa!���188xͽ˥��[�5���x<�w�o!Nj�v&77��K_�Ғ��*�:����l �%���[FF֭[������ǴH��w8h|2DDt�xG��t:�q�F�����������%6\l�x7 �����^��R��P�Yq�����\����egg�v8�B��!�= >
�҄��?�]���X�v-RRRn4˘��G__�.�x�Hd�Q�Ys�4��y&�����PQQ7��-^��������������_�	�k[J	����3 ��!)��i!�4�I �W�� �M�J�M~#KHH@yy9���`��o�_a��)��'��r�6QH���ƣGq"�C����ף�� ����p����09y�o�ʅ����4�gDJy�f��0
��qq/3 ���Y ���W.�p\+��v�����D����dg"����Atn�Vvqg���KLL��͛QUU���n���);S)$K)�B�\<��4-��x:�0`��bZJ����+� R���B�b 뤔�7���U�PYY���NNNbhhH/��Fa��Ś�
܁�{��;w��QtJNN�֭[�f�tvv^�#�K\ >)����B�|���s@ǥ��ԥs�i)�����\:c�R�!���9���w���������+l���Qe�_yk�i��(z�(���t�޽���������O(ɑR���Xl���xf�mR�\<g��Ŏ���L!Dڥs�r)�: ����!�@aa!***���zC�֊:;;�gd;�q}ggD˂�DDu����_�*��ى6��Yt��l(--EII	��ݍ�����W^�gE_'''������q_ؾ�ܹs���>�3�bSB��hm9��w�D �ع�����q=�d)B��� �����N*�B�����+��ILLDii)���,߱�J333��s�ٽ��(Vd�����g�l�*>11�.�
��ɨ��Fee%Ν;���>n�����_5~PU��Q�.Bdgg���".��utt(���9`p&DD��o��]{U���a||��7�̒RRR�y�f�Y�]]]���G0��M�� 6.�W�*Z������������n����BJ�8��Q,���233�c�LMM���CCC��P�J.)� ;��ܳ\�>f)v�������Drr�M�;����+�������ل�(�������Қ�&��L��V���Aqq1���L�,z!PTT���"LOO���������7;58��塨�(��c_�����{{��,�LȈ��nFҥ�'������,���QYYiRf�#77��������� Ο?����ӂ�fC^^
�����D[[[#toǄl���f�8p ��6"v���҂;�#�/[U�n�:�]���øp�.\� M��N.�(..��ב�u���N��{;Q������Y�}oii�m����ϯ%))	���X�~=|>p��.�ZN.����(**Bbb���jppccc�xyk+����-E�]���4l۶�@ ��������Ȉ�iA��������ô�����8 �L�/,p'"��$B!l�]���/\�R����v�2)�蔚�z�vdd.\���(fgg�!))	YYY���Cnn./�#hkkSvR���!8]݉�(zm��4�ډ@�%]WW������dRf�%))	������122���i�.d��������a���|>�.��ߏҳ�N�DD����P�Ԅ�-[������ܹs���0)��'�@^^���a����all�f:��t������FAA�=\"�DKK�rmǁ�gCDD�)gpeg�꺸ONN����())1)���X?//���0���{�w�ޥ�������w���ihkk�Ņ��q�{"�X�;���t:/7o����|�2>>n�=���@ff��s�Xo.kx孭&dD��DD����q��[1RPpU|dd���(���Ĝ��ˣ����0::���LNNbfffY� !���|��2++)))��ku��������Q}��	�G���c����p�=WŃ� ��ڰm�6s�a��U���`tt���Y�KY!���������,dee�`�H���{^������#���tUW#��*�����4����Dii)JKK!����$FGG1::���i���-���p %%�V���Gq8x����[9��������DD[v��&���thΜ9���|8�N�2�			(++CYY�����������0==�lS�\.�U{�xnIGG�r����	�b�v"�X�;��������JTVVB�4���attccc���Y��			HMM��O����D�k�R�5B��7�`�v2OG��(j�P���
���/�FR���!77��eא��t�%,pqC���1;;���i��~h�M�!���N�v�v�IIIp�\p�\HII���-�e��^�C�՝�����>@�-�0�j�U���A���"++ˤ�b���DAA�U����033��������=��f����v8��v$&&^�Ǹ\.N�����[9��t
zzLȈ��>���ql}�}4����⋏��n�jRf�iq�uFF�����aff���������<4M��?Y��]<_q8��\RRR.���a�6??���DG ��^{̈́���h���a㑣8}랫�@ gϞEuu�I��&!233���y9/�[�ܻ\yW\,`��l����J^���p��������'DDDˎwD��n���# ,,,\u���p��e����GY<oIHH����#oܹs�0==���>s�~�4,p'"����ׇ��O��i��͡��k�FU�҄�/N���@+���SSS�xqg'V�9cBFDD�욆�_~/��o�֚��q�w�Q�2JJJBRR����N�r�����ե�;��q�o��-�mￏ�[6c2�Ru`` ���Xv	K7�n�#==���f�bymmmʉ>[�?�ԉ	2""�����tnڈ��ԫ⽽�(..�߹������ ---�B���w�A�b"��-���$$$��`ʦ�`�M�TlYFDDQo�o A121�Hb�h377��g���6M��/�bBFDD��J::Q�ޮ����(�4E���e���w�C��������P�577Cr�0ŀ����ic��v�	�JI����7��ť�ܻP̸p�|>�.�5<��&dDDD+�wDd---����C��66nBFD������^���8���B!�<y�������.�����>D��	�r���k�+~��ە<��I__���t���Ql:|؄���h���9�R�����i�+.a��I0DSS�rm�k�}8Ŷ��N���G���@ww��	݀��477+����
l���DD�xGD����]��>�
��X�NDD1aӑ#���'''���iBFDק��G٥�55�m�gBFDD���ư��u�P(�ӧO�AE���Y���)����
슮�DD���������n���5E�����~]���egΘ��8)���� ��,�h��Ԅ��]��t
�ɗ�ȒxGD�jnn.bS��_{NE#G"#�����b�-�ޗ_�Pl�;::099iBVDK�����	o�+���8�$"�ص����66��ONN���Ä���&���ӧ�c'+��Q����DDV�>6��￯�U�i�    IDAT/�}��QE�.���_w����MȈ����=8��]\J�S�N!�.��"M�K��í��nBFDDd�Q,jjjB@Q�^v�,V���#��DD3
��`�#���'O��E,E��CvU���S�P�/DD��pϳ�)��uvvbLq�Id���n��e��4ƈ�,j��w��?������=�̲�����f�ڞ��@:��DD���ͷ�12��OMM��ٳ&dD���,Z[[�k���2R��Έ����p/�(���������I����MȈH��DDSv��&���u񙙙�������ى��q]�55��^yՄ�����}}�z�]|���Q����VH��^xI~��Iъ��B�����P<����Ű�̅�,�O�Ƃb�]qg'�MȈ����p�3�¦(������	Y�I)��Ԥ<�+omCUS�	Y���xGD1����̙3ʵ;�0��܉�(��5{�9�af�ׅDFS�R��g�C�ܜ	Y�Qv8��tq�ߏ��2"���i8q�r�{uc#J�����2}>�|�-���ӧ1��Ν;�|p�������4!+""2C�� ����..���ӧLȊ�j�)SS��Ev@%"�';@v�;�HSʈ�
�p��q僋5'O��w�EX�NDD1'gp��ť�8q�����L4??��'OB*.Z7>���n�"""C�4�=�,�Ψ�ϟGOO�	Y��ӧO+��icc��ƛ&dDDDF�|�������Q�L5>>���6����"FD��|����������Ǖ��DFBgg�~AJ���H�<"��b�4�Ꭸ���wDd���fLNN�⮩)�}�U2"���DD����>�Ο�Ń� �?�����J[|d��v���a�[o��"sx;�9�\kmm�m2Mgg'uq[(�{��&dEDDF[j����;��i���p��1e��S�QɟM"��d�p�s�á��E{{�	Y3338u�r��hJ�����ec���(�xGDf����yE���w?���L,p'"��d�p�3�"q~^�633���&��x��܌��1]���_>�<|'""����(VtF�R��ɓ�QD+�����ٳʵ�"O������55��_zY���ߏ��^�3�x�8"{A��.ml{_V��Q|�����וk]]]08#�w��El��5<��orJQ<���(���ŗj�G�������ڪ\�z��;gpFD��w""�Y�cc���g!]ѥ��@�Rz{{��ק\����}���ل����_"ubB�6??��d(�ߏ�'O*�V��a�{����	[V����`||���(�577cB�wv�x��FDD_664`�ɓʵ��&LMM�ų�'ObzzZO�����'�LȊ���������*�Vp��	�B!2�x4??�'N(�J:;���O��:�����bZY{;�8�\koo���38#�G���_�n9|U�N�E���Y<�ē�)hnn6!+�7���رc(.V3}>���� [ŭݯ����$������Q�iD6��ǞY���'EDDQ�_���~}���ﾪI D˭��CCC���p�3� M1허��O��,>��S�;���q��!���+�����_>���X�NDD1oǻE_\�x�nc�������ب|]]�ۋݯ�aBVDDMrq׋/*����p��Y�3�x��'Vu�s��で�F���5[(���|
i����y9r��b�����"6���!T����`��'�D�̌n����������ŋ�����y��~%�gDDD�,{pw���r����hoo78#�'RJ�<yRY7���'�@��oBfDׇ�DD����/��LE''M���بH�Q��͡��A�5ub�?�$l|�JDD �N����G�k8��J�Q-\*�I���^��&"�����_�:��~;;;���F�ъ�8"�����yǄ���(ڹ&'���O��؟LNNFlJC�Q��i�����6l;��Q,�:݄-�+�:;;���mlB7����Sg ��_���kDт�DDd	��'��@ �M�jaaG�U�\9�A<�ēH��5!3""�V{^��z�kmmm48#�����?W;Dyk��Q4˾pw��%�����?�,B&�Y���qGd��{{������Q�:u�{ZVccc����>�g���"���(����̙308#����6�?^����!�=u����n܉��22}>����ʎsss8z����6э�4�Q�@��~�9�H�����B!���S�Pt�^�=22bBfdE������S�U55a����ł��NE�;���P�����L�� �~?>Q���&"�k�|�6=�\DKK���UMMME|��2=�O����;H""Z�-�}O>���*�ĩS���X�nBWWW�� �Ϝ���64���w""����N������֥.Έ���i8v�&''�뷿�
*xhNDD$���3?�9\SS�5)%�;���q2#+9w�:;;�kK헉�� `���`CC�rm`` ���gDV377���,,,��� >��z��>]�������f�Zoo/���Έ�fffG�E0ԭ%���S��i<�#"�����ӏ���	ݚ�'N��}d}}}8s�r����>�KṆ��w""����&�}�����8>�N�tS�� �;����w��Q]@DD��51��>�(��@4M�ѣG1::jBfd]]]s��q�SO)']鎗_��x���MMM��N7��������+��_�x�4�"L�!""RR�g�Ei���wggg��k����ѣG��A|���2!3""�U��)|��ǐ<=�[�hhh�_�i}}}h���3kx��áx�G�X�NDD�����T�MNNF<�"��Z_&���#""
�>:�O��N�~D�4466r%ݰ������K���R��g�EI�B���>�:u�E�tCfff"�CJ��(={��Ĉ�(��B!���ȏ�H������ܻ������Ç177�[��y�����ź��1|����y�Z0Dcc#����n�RM)�����G�b_C�X�NDD����t��rm�C)�p�@ G��8�r��DDD������'`Wt�^,r�p�	�Q,joo�X��g{\95���(������F���r}`` ǏG�#��:LOO�ȑ#��n}��;y�ଈ��J� >��zdFh��ۋӧO�ȝ�����=��-%���K(om3>1""����|��'�wD�PǏ�]���.�D�Ƙ<;�O��gHQL �v,p'""K����Q�Ԥ\[�k�%���8|�0&&&��e����!x(NDD7���w?�l��0)%N�8���A2�X��҂�Nu�ݔ�i|�Ǒa/CDD���<>��_`հ�Plhh�E�tM8|�0��� `ǁ����gEDDV����ӏ�ic�f5����BC�4::�#G�D,n��װ��q�#""�)���=�|f�;�����9s&b���Y|��Ǒ1:jpVD˃�DDdi"�=�>�������Ø�KER���8r�Hğ���<�ē�)^U]���f�����.RJ�<y}FlS|�R�ԩS�0;ub���O��{��H���gy$b'���a444��(�D�~
`��obǁgEDDV暜���ӈ�����A�3�X044���Fh�s:!%�|�el�0=����fT���'��]�7�� �7)%�����ե\O���gyY�@1��DDdy"��^�6xX�>77�>� CCCgF�l|||�fff��U��po���DDD7ju[>����\XЭI)��Ԅ��&v��� �=���~�z��8>��H383""����Y|��ǐ�۫\]�;4ŧ��^444�/u?���!�#""�K�����S����q�/�;wǏW��B������ф̈��������N��3)%ZZZxGDW�4ǎCo��:��>��G"Ne$�,p'"��p��,RG(M�p���/)��������XP���F���,n'"�eUt�>��_ Aq�	\�������Q	333���1a�d�χ���G�݌��y|�񟡸�S�>;;�?�###gF�FJ�3gΠ��Yy�.B!ܵD3
""�����S�=��S񦦦p��!��ax��B8}�4Z[[�{��ᾧ�u'O��ŋ�s���Cb�x}}}��G  �ߏC�axxX��6>��=�(�#�!��Q\�q� v���rm������|���z����Q�����!"�P�Ӄ�<��"`�|>vG�s>�~�ağ���A| ej��̈�(8|��X�֦\hhh���8��A,R	
�cϿ��Ǐ�ţ��y|���Q��kMG#�[ܿ�?^�n�4���/Q��jpfDD���w��U�gÇO&���A�¤hpDQԪ8?�?����S֢ۧE���`3fd�L��@BƝ�~��ivb��\�������b'��>����ֶx����K�������3�i���g� q��0��]R�E�ȱ}���%��˽�:͌����Çso��f�=_�#�"B�����-v��~�@��vTƦ����	���hj���r�� ~�2�x�?G��������UUUL3�.]�p�؜��x��E'N�y2 ��9##������~>66'N����z�]���[�sݐ7wp0���Ü/w�����=^xｸ�q?w���u���(//����q?_��b��; �����?�!���yOOO|����ٙ�ɘ
.\���Ҝ߳FG�ɝ;���<O�t���#^}���9�����(//��u��cǎEMMMο��G���|���- ��f��œ;w�C_~�����ؿ丙�kK{{����_�/��^���y2 ��=:���?Ž{��<s���8x�`�q2�Jkkk8p �w�E==��[o�ʦ�<O �8{.^��뱢����_������3�i ��ĉ'���2�����J��&	���n9y*^y���1Ǜ����q��!ǮqMMMQVV�r|џ��/��N~W��� �����ŋo�k'؎z���(//�!Q�5����QRR����~>cl,������33�<O�tw��x���r|��퍒��hkk��d�K&�����8v�X�[f���ī��K�; `*e�q��}�������q�twwOx	W��KN�8�9��jh�W^#n��)t��K�����-��FCCÄ/lq��p�B���Dk��X���;�w\��	���uw�˓l`�q��t�����/0,io�W�x3nn� ��1+��'>�$��ޝs;jOOO���:e��hjj���s�����S�]R��� ��+����~'�������h?~<N�8/c]S.߈��ܜ�̚�����{1�o��� �ok**b�{�Ǽ��q?�ÇGEE��.טɖDDl8|$����1�& 0+��m;?������Y.p�lY㜑�x棏�޽�",��%p`ڛ;0�}�a�?r4����(--�]#:;;���8:'ؾ���"^z���<N ��f������cv���###q�ر�������<��mpp0<8�x{z�7ߊ���<O �j�ٳ��oƲ\ۤ"���5JKKゟ��	��������?\���Ɩ={l I�Μ�W�|+�=��̙3g���9�����f�ԩS.�96�|�����g1��� H̝���>�99�]^.��kÏY�xCoo����q[uM�����=� @
ff2�خ]���%�~���3�_�\�:::bÆ1w��)������H���DKKK�3�2����Wqg�Ao����UUqcWW�~��8���inn����شiS,^�8���f�������1����W��c��mb $e~_��λ����Qy��3f�˙���(++�իWGaaa̜i�զ��?*++���;�y}}���O㖓��8 �{���Ko���=�w�5�˷��Y�&V�^3��~C�.^�ћ㶡���'��3��>��� ��s[uM���F�~�g��ψΜ9��ݱiӦX�dI�'��������>#���>��Ә�c�;\K� ����ͧc�k�F����ioo����X�vm���U���=���bxx8�;;c�_v���H��g��߈۷G�[�=������|��ظqc\w�uy������b�FGc���q��<N ?ެ��x�/���>���r\Zpÿ���A���-6m�K�.��I�we��hll����	oZ���v~����8 �4s����O>�������1t���r&��D]]]���Z(p�d2����N�ʹ�4��X��]�bn��� ��_��W���gD[�_.p�ҥ8x�gDW������������gfe2q�7��]�e1òF�	�; �/7vu��o���m��?�q~(����hmm�;�#-Z4��cDeeetvvNxn������� R1kt4���X��{_|!����\{{{tuuźu��[n���Xcccq�ԩhhh�0��ܹ���c�sy� ~�[N���~�����Kq�p͸g�СC�^zzz���"���s������Uձ��-�~��h���q�\^(�r��ذaC��&`�������~w�=:�[" �U�ψc�K/��$ψ
-nL؏](���|<��Ǳ��5������8fe2�e�����ӱ�c`��q�]�p!������o���5kV�'%����hll�S�NE&��yn��`l��X]]��� �?w[MM�W{{������HTTTD[[[lܸ1,X��)�HgggTUUť����f㎃�⁯��Y��� �C����׿�}{��8�m[�͜9����j�*\2<<������2����ɏ�K݈�UlAoo�x��8���q��G�]~���]]]�~��X�bE��d"���QSS�|'Y���?�K�4�b$ H�m����7���_}%�n�m�3###Q]]�q��X�pa��d"?楼���G���_~�-kd��
�����6�}aG4�{&��FCCC���Daaa�z��N�l6---q���������x���b���y� ~^7����G~8�>�52���1���;JJJbժU�v�ژ;wn�'�Ο?uuu���=��}}���ϣ��6O���kF6�*.�U�����g��㞻�R^SSSŲe��<)?4::������8�Ҁ�fc��c����s���7  \!3�������U��qa��q����ǣ��1֭[K�,������H444Dss��]f����c˞=� pM�������q������h�fzzz���4V�Xk׮�y9���/^������e�y����_����<M���$���ů���h.*��矋�E��=7<<UUU��������M���������/Nxn��`lٽ;69��l �r3�����X[Y��?g֬�\6��3g�DKKK�Z�*��������[���O�I,��X{�x����� ���[[���.*�/=�D������G���n�)���bq���+��Ҁ����$X_��[?�<V66�g8 ȣMM�~��8���q��G#����.���cɒ%�nݺX���WF&�����hhh��I6�.���v}7���i: ȏccqwii�����瞋�k�=��f���5���<#�"q�ԩhii��D���<#z����'���; �Huu���1�>�X����Z{pp�[�
c���y�t���鉺�������ꪪx���<? p�Y���}�a4l�%�=7�0�ˡ{GGG�^�:


bV���<��ɓ���2"�;[w}�Μ��t �3�����q[m]�<�|�.�����o;)//��I6����������I^��96���ǽ�|�&�� W�Y��q��}����(��|��~{γ]]]QZZ˗/�����?~���.��W__CCC��=2�������̱�<M ����/��K    IDAT�x����~q����q�]~F����f͚���v`~������MMM16���E==���b��w ����-�w�m����;�����y���/�;��ͱq��X��~�����������I��,�t���*V46Ɓg���͛#r�(322������k֬�[o�5ϓ^����?��'���쑑���ocsi�� \��?�~�a���({��X� �ٮ��(++��˗ǆl�zzz���2���&=���)��Y��ݝ��  ������?��_��o��y�r�moo����X�re�_�>�̙��I����Ψ��������W=�/bAoo&�4���/�os�o�5���ψ2�L444DKKKFAAA�'���ꢩ�)2�,	������%qwq���w �	���ƫ��U��G�n͹!5����Ν�_===�����]����l���d 0����?�4�=�~*ή\�����`�>}Z�~�4N�r]6k��b˞=���|^f�~W�ԟ���m����L�e���?��^�dI�������O�/8>�|�uVTFLr \���X�h�������{��^�.^PP p�Z[['��o����۪k�4 �e��Pl���Xw�xx��h��������+���aқ}o�����m� �C� ?�̱����`�;~"N<�@�x��I,�2��t�P��mq\��T� Sbyss���[Ѹ~]�?�D�.]:�#�+�ݻcik�T� Sb��`<��ĝ���ǣ��;#�##���t)~U\�����@���G?�[l� ʟ�7�9���������u; DĲ��x��w���(ʟ|2z��<�#��O��-_�_�93գ@�� ��34����#[����˹��<�fc�wq�7�Ă�@d�q{uM��E��w��m��҂S=մ���#ؽ;n9yj�G�$����>�4�*+��'��梢�iZ�=2���%�q���T� �Y��O����\��w��ի�z�i���\Rw8sFF�z HNA]]�Z_��7��m�G��7N�H��M���{����ک�����ɼ��x�/c�ٳS=ʴ6wp0�عS� ��̱��p�h�Q^>գL{��+q; ��g��S�h�ǘ�V65�}{���$���Ŷ�;�z�i���.�).��fd�Qt�x�]��G���|���~$�;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�          ��;           I�         ��c׎    �[OcGq,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�!K�    IDAT�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�     �v,    0��z;�#     `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap�صc   �A����Q          �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           _�3    IDAT�;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;       �k�    ������8   X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X� �];    �o=��        ���          ���          ���          ���          ���          ���          %%K�    IDAT���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���        �v,    0��z;�#  w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           R�;;    IDATw           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w   �صc   �A����Q      � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          �k�    ������8��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ���    IDAT��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     �];    �o=��     ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�@�ڱ    � �i�(�          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap         G���    IDAT `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap      �صc   �A����Q   �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;          4A�_    IDAT �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;           �;  Į    �Ǝ�        X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�        �];    �o=�� ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���         ��Y    IDAT ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���          ���   @�ڱ    � �i�(�       w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w          �صc   �A����Q� �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �        �P:.    IDAT  � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �     Į    �Ǝ�    ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��         j��    IDAT ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          �� ��v)n#ð�0	8��V��=��J��*130�� �UU��u]?�K%����-	         �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w           "�          � p           ��          �w��q[��~�3Y���ǝc[ך�nwǙmq�����b܁���m��Lch|6�в�����\e�c�f�3�inw�s�i�����m�YͦW�)4��MS�18W��aC���L��/Իִ����T��܅�U�'��������I��⼺�/�W!6Ϸ��N�N��{8�O5�c�Q�1��p&0����������]��� Z���\e.Cc�ɽ�
myU���]�1t]_��А��ߺqe��ʺ�C����\e6�k s���ʹ��C{�o�O9������|�L2���'pgqN�G��Ө&An�к*�� �F=�����n�G�1t]Ol,аj>n=4!*K��|��z��x�ͩ�VW�Q���x ^�j�oL���u�RZv��X���83��b<1w�E��/���/K��|�yK׹G������#a10�)KdA0��+n����:�j9�n�#�6��G��R_j��F�rӕ�T+�W��%,��b�bL����}!W�XM�g|��U;�BI��W<8C˪h���F�����	�Y��u�YLahtl1@��1f�'�ld��U�c7D��ӓ,Q����83o�`)��L�)Ө����9�S]W��z!I��{8��Uc��v���8��|��\�D�s���X�4Cp�w��5j�]w�d�.7�noo�p6m���{y��M}Zqz}�s�3�j�9�v��3�q�+l,L�GN��#��l�7n�2����^w��sS��\�V�v���ٴ�W�n�]h�ٍ��9�}�����mMDcN�����j���ٴ��O��:и�b�1w���c�.�Sk"ZtZ������Z�iZh�POa�2��=>v?�P��8}ߝ��s���U�����=������α��;q������P�#]g�r
�|��E}��o����b^bM4�r����������E�<O5����A՚�zh|�ժ|�К^���B����k���
p�y�wn����m��������W�w_�\�.-;���;)s�h|�5=����C�	�Y$��yT����_}���U޾�-F6���w6x�^�ֽ*6��W�WFb6.i��v۽)�5ƌO��R�_^vEd`\_���������b蚾�믙��u�^{�L<��R��<��n���Ѡj��E�)�]g���}w^��Գ���Gti|�B��"U���ĕ���1�i��c6h��Ƃqd\C�KP�έ��W�1�t��t��~�9n\�f��V���q�Ѣj���l��y�j�rzs���:Ӡ���*���M���"TZ�V��;�j����;*�H/]u�sh_����.'�uw�~����>����	�Y�j3������Owuu�s��l9�f(��O�t��<�l���~��������qd\777�cq�ÍW���Ab��j�*o���&�QU4��X�t߾�ksZ4��6_ח�>�.w�A�q�\e\www�����q_�a	�1��{s��Us�!ZeM4�j>���늗�AK��C�~��yxx(���?#pg�>��q�X��墘�Y���h�?�^{hч?��9vi�:��z���Sw��(4�������Ud�4�����c��?�������]�U��l�fh}��X�B>|��@n���Z��Zu���h���M�S�[Wu=��9�����y���ud�4�>�A�w�|�����y��|ѝ_@1w�н�_>chӏ��ݛ�7_���鬉X�����Cw}}���iӗ/_ʽ� �	�Y�����u�G�b`<C��?��6��~���������/E�dh#���:���D�q�[�U�W>��{w����l�?{���u���� 9D$"�����m9ɒ眩;s^ϭ�/flɖ���
�$[�#�sj��� �"{5����T�T�wX�W����y�k���r���R%��S��~"��Xu{�2��m��3��@>0�X��@ `�m�ly�cf����Ӄc�]6���<��h��U�J�m~>�9�����3�`�<�a8ka^98�pXa�:Ŵ�M�����?:8��ee @w`�pG�2mv�����~��s��t�̦=�S�����0&�D�|Ҹ��rC%e:F�9�y��,V��j�s�D����r�,S����H&��d���٣pDL��`PQCuT�i~��[��h��W���P4����a�Bg:W�z�t�< �sq{<n���Ӟ?*��`�P��3m�� ���:a���v`�    IDAT�����G���k �����n>
ɰ7�e��t�=� ����U�!�`�H��3�K	�6a�qe�,�ͥW�Y[[��h����
���w�˥T*u��3~�߸�4%A��8�T��b�s�.cmm��Җ����Vb^9(����˲����ԡ��t�����|>cR���G���eY�NL�;��u~AE$ ����I�u
{��a�=6���}#Sa����-�o( �Y.�w��`u��[8/��o.���޶�L4�SS�i���ֱ֨O�eiee%�y�ܼ��l!Ϝ��J{����0��bZ�F�T�AA9iX�$	.H�i�)J��N�/�\�a^Y__W0��h�i^����ࢻ�W�߯���"���_86v��������H$B���d(<R�L�}��(�kk���}X��_04v��a��V��pVk�'���b1cR�t����LwD�d�������Yk�	���U�������g��E":99��� ��?0��,�H�!�'��kl��?<��� �����1q����$�Ic o��PP:fgUe� ��?���NNMQ�y�pP6C���F�ƶ�����Jn@>9c8[Y__��>-//�W��,�q����5>�2C�q�*�cY�G��	��o _�,K���k�өx<���LAb}��Yp���=����������1��p�,-�ΐ�kJ^�ޘ�Gm���;9 �#��߰8�T�����c�TL�
L��j��Ӟsa�?�ߟ=W��XF��hT]i�����p�i����fY�31e�Ȅ�q�݊�8�0��W۬���{�.]���@��6v��uL�x-�˪��5�\q"��##i�WWW��3���k
����9S"<vǲ,�P��*	C�6`^�Ӽ��t��Bu(0}�{���u�)���<��0wD��!���ؘJ�n���YM~X\\Tʰ�:C�"�ڬ����-?�nO$�l�GFe'y�ٍ߰�b^�i�W��}���(<�.^�=�YCpoi4������y%
�ᱳLsr�ꪱM9�o*�~��ͥ=_\\4&�bg.��X푤
�9K2��(�>����P���(H���jXs�=����`�Z]]5w�e�Q���o���{�'��z������y����PZ�H��Ǵ?*ɐl`g����3TE]]]���H&��`��W���G?  �2^%iff�G�fggI�A�955�2C����4�"O��t.M8@!h\]U��|�Jý[__���N{��`D��>Q ���Tb��}zz:�9�VVV�����BbJ���bTqBSSSiϊ�I�>x��� G�m~^U�s����Y��������wxXE�s\����Ճ��V�
�DL�i�x\�����a�ofO��LgT�T�.�(H5^�Zs��⢱K���^���Tj��`g������V�3˲�x}KKK�*(_�u��1�z�K���7��alK�����2N�:H@+J&���{iϹy2�5^Q2��n���h��p���Ҟ��q-,��`��I�������4U�����>�Ϙ ��2�O�c1��?#��wxX�3�Q����h}}=�y���i?�a�,=}�v��H$B��0�Y�.p΂v��}cq��.c��{��ꋂ�;2�
C�F�D{���!�˕���ؘ*�,�Ⱦ���D"a,p��eZ�]��;"�I���׶�������L�`�J�������s7#rǕk�Ӟ�H�w����J�Wo\���之�}g�����޸�nc0Ǚ�Ac�6�P�T�ߟ�<ӿ�0������j4<�ٕon+v�ڛL��}�@T��x\��6�y$1&�#���ɴg�TJWo���h��9����8g���gU��9P(*�A�3,�tn��2+�r�,�Ȟ�x\EJ�흩��,KW��@��Q�כ�|aa�*�{�p8Ҟw������IW�_K{fY�FGG�0��izzZ�H$����3V) 
I�ܜZP������H���5^�z�i���W���􄱍����eY3����R�r�`��dR��I���b��A����k��M ��x��kX�{<�!?�%�IMLL�=/N$t���Km �e
F����u������#��x�0" {J�Q���^�0
inn.#:~,���Ȉ酮\�q�r��7U�L�=Sʐ�t����R��=����nc�Q�䤚蘌fK�t�F�>��a6::jL���5wD�~�H:95��+i����Ȥ߅p8l��^���[�>�Bd:�ߺ�*��<x`<��z���2$������x)2>>��Xw477'��Bu���9 IOݹ��P(���쬱z0���$�a.99m�k���us����1%k<jzzZ!ü|��]Zf� �F�:�}z;�X,�e�.$�Ic¯,KWoP����7��n8O���4���������ҞwMN���F@U~���=�B�b>xT"����x�s[*��+A�ʔ�Ǟhw2&��|��Lݮ�Abَ���U���I��� w�����磣�\�� S��k�Uj�"
Q�Ԕ���Ӟollh�P�����j�Ի\:30���Q����o�I{�Ǎ�=�/�H�x�[�L�ٯ����S����eY���x<n�t�,=�a�	�z�K�CCi�#���4
�Ơ{4��7�@���wƄ<.[w655e��RÚ3#��<��o�M{�1!e��Rz�_faD@nz��uc��Lɬ����	Ew���ݧX	
��o�U9{�'233c,��5>����,��-Eɤ����e���m��vE��⋣�gp~przZ=����p���m,//g<��-���,K�~����������b1����~�@>{��/UH?�[ZZ��������ac���7�~���;j2T��z�Z�?���c'����Q3��Q�^��c����Yc�O�+��TH�ٯ���Б(e�^�<�bв,��@Z__7&͔E�z��V�+�o�f}=��ᠻ�6<x��!h���;jZ]���T���+��;�$�IŶ��z����C!=��daD@�(�����m/hzz:�yI"�W���,��Mg�j�7���i�*����f,*�>O�K`�p~�O>5V����0� 
����w�~򩊨|<����C;�D"���3��������au��B*�F��知=�,Kƪ6�nvv֘�W���2m'�G�R)���G��$###�T�fqqQ++�A���0�I����eY�w�10��MNN����=op�t�B���}.�C���7'��x<���A��s��R�@F䎒DB�~������EI�0$FWz�V@�+�|�:�٤��6[�x<���/���p8�r˹�����~?]h���ݻg,�t��k�dG�`Y�^��cc����q���%���0�*�F�"E�A�;�#����~}��nhhHa6��R)ݿ߸�R��* �ٯ�6V���|:<fffƘ\T���?���П���X,����,�#>���2[�^��S�	�ҜX^��{�Ӟo��/T�@ c ݋��KW�Oߺ���i�#���0����x433��²��'t�$I��W>����aaa�tY�2�6;z���,��=����e8;�.ȲPm�z��ύ�{�BW�L��O�f|755%�%144d,ztbyEg履Wɲ��_?2����J7�G���(L�\�����faD@nkXs����Ҟo[�`ɿ�B!�=��/UIQ�@�<��w�3^�3i�������H{^�eO���Ѩ~�+����q��ǣ��	㻗��w6(x����������TF�{b���ݻg���RW�9���矫�P�#jhh(#�=�x<c����I�%hx�fY��_?RI"����tj�yI�����߹�v:X5������w���
pf )s��DB?��/�q�<��ǟ�ܐBQ������vML�o��@ꜙ�Sw�=�+磦���k��x\?����j@�jt:u�z�=�)��-..j�Pt�(��O��WΪ H�}���M8���I���ɤ�ݻ��ai���� p���ߚ��/ۃ r�ͲtrfV��/)a�?�.�(���M6�-K#̾��I�.Vm��~�ޟ�h8| �/u^��%%Z�:����t���AYYn����}��1��`P�}�UF䖲pX5>�f�~*���Uyy�jkk�0�ܐL&u��-�!n�ǣ7�{O�T�2*I$Բ���+Wd=��	J&�jnn���/�J��ݻ��|i��~��λ*��	���`Pe��ΜI{��xTUU����,�,7��qݺu��9����/��>�ہǴ-,h��)���y�J��t:��֦���,�.�VVV422b|��#�xLi,��KS.H��|>�JJJT��|SH��@��GU쁀]蘙���s
WU=�<�L��v���]EE�[�pyy9c���?�D'���xD@�k_X���[���G��R)�\����\.�=������Iq2���M\���c�`0�h4����,�.�,��ݻw�n(U�����X���!�0(�FU�t3�����Z[[�4��Z\\�X��ٯ�����M�G���k��i�=t�,Kkkk:q���ʲ4��	�B�u떱�U�ǣ7��A���N�jj�joK{�r�
6Pl�P�����+N$��;���
�QU~��I-����[__Wqq��0��ڪ��2T/)J����S�� ��ʊ|�M�.?���TWW����,�,��ɤn߾m��bz��wUA5j �ͲtrzFS/)^Z�ȻD"!�˥��vgi����x2v��ы���Q����Q��T�'O��s�ݪ��(�b;���Gջ�Yp��Rj���ĕ�J=�>��b�x<��r�t��}���a=��퀀cbsO4�ɋ�xlO��zO���t��c1���Y����t� vP�,���w[瘍��G=��044���մ�6��/����dx���dP��(^Q���δw~�_�TJMMMYY�8�3Y;�����~�F �%�e���&._R�n�T�a�{�c�,�����ƪ�%�����Um� 
Y�̌�ΞS��?Rav�غt5����W?��J���.-���.����v\�˲�������?���?�~	��ΙM�?�XEyڻ��5555��<�]�J�R�w�<������� l��bjp�i��Ŵ"%�x\^�Wmmm(�����+^�׫߼�
 �h���R_��55i�N�jjjTe8��W;큞��?�?<|ģ���PH�~��ΝK{�F�������޽k\�Թ\����	l�����6n��b��|jmm-�=Q Э[��H$��Uz�w��=��Ȁ���ʊ���Z?q"����n/�NW###Z\\4��z����{��G�?܁mt����n�X__W<WsssA4,..jhh�X�����o�yWvZP{R��uiI�.��vJ&�r8jjj*�J��`P�n�R(J{W�J�~_mY�ۊR)�������iU-˒��(���d2�{��en����z�ڵ#p�����b��N�S%%%q��J�488���e���z�j�����I������J<��kY�VVV
��{"�Н;w��P��ٯ���[��xT��S���,�bzE�H$"�˥��ւ�Z�r�t��%A`��~�_�S!�m�,K�&&5��S���VWWUQQ�C |��*"�8XM��J��Z=u*�]0,�`T�ө�w��.��~��߫2��Ȁ���=�Rooڻp8,��S0{��������Ѩ���;�3t��٩�)���V�P�h��S!Tr�,KCCC��{<�k�|������6l����19����K{��������ښ�A�3335�����o��;Ur9<�j�O��k�9����摭 ���ڼ����Э[��F�_Z�^��c�Q	Ȩ,���iM_��dI�#�,����JKKUgX��x<�m�X��^��#�'P�L����ϝS����v�}��N	4]��z���f�Ry(�����D��.W���+++�:p,���ￗ��3���]����G<*��jY^�U\,GWWڻX,��K���Ě|������������z��?�"�%{,��IM�Z	Cw͵�5���!�;�D�=p�:gg�����-�](*����e�.[A�?��Y��b��h4*�á�����m%͘*�%���{����S)u��i�L������U$щ'���h5ùJ�ܜ~���V�a]`�pvP�J�{|\g�(R�`��zu�ĉ�;hH�Rz���fff���"�����<d��Q������3i��R��G��:�������_��w���"R��f!�̓=˲��ؘw�[ 666��;gf����3�
�>��quMNe���|
�:q�D�U�ú}���*��,.��?��v��U��jZ]����i���f�XQQQ^���~ݺuK���G��Ƈ0�Q�ܜB55r�����q9��թ�w�Y�������I�R)�����>7w�#���HDs�p^�Ǌ	H����u���@�!;59���x4���TSS�J�0ǙeY���μvI&������Qd�9;+}�<��i�������Un�Rs����khhȘ4c�,��������,��%���'&4��ӊ����������jnnλ��H$��w�����79z�we7t� p0pv�$��!Ƚ_QC�H$��������%I(��۷�t:���"���?���8�����Pi4���޴ wi385
���9/�R��FGG5>>.+C����7��W_�Ȁ�Ʒ�FǪ�z����z��x��Ԥ���q����;w�;@Hj��כ��I%* �V���̬fϝ5�������Ae�����p�Ν;
����'�W�ֻPi�9���<չ=�;w���v���������ݻgl�-m����Vc�955%}�<�-i�ɤVVVd��T__���XL�����Ғ�}q2������'&�xd@~�Ժ��٧���}>��n��������ڶ{�f�@���Y�����<�)}}��x<���e������6#<x�Y������59u�#�G�Ĥ֛��~�Dڻd2���e��0�G�DB������5���Rz�Otf`�h��hT]SӚ;w������W�4N�S�o�V(2�o\[��Ｋ��' � w`�Jc1�=x���n�m��.I$����X_�l�E"��J�_���ߩy��v� �,-�nݫ��g�[�c����:pl+�&S�[�e���>��k׏xd��W��mn^sO�S�p����WSS�JC��q�L&5::�����I2�cc��{"c8@��z��5�_1Cbo<���ұ�|�q"���$����o�@`�_N�N,/k��9�A�PH+++Ǿ�r"���А���3�]����ߧ*�6����q��˴��i������;�U��n�n߾-��o|o�F��?�Q]��G<2 ���|:93�����HD��˪��RUUUFx0R�����4::�q�9=Mp;p��R)�?������J�����p8����c]�����֭[�.�Ѩ���u��v`_l����1E�*���0~��v�E�卍}���Z__7�/N&��>P�����_塐zGG��׫��y뎨���X'�X����	���d���/�����v���AI<���ay�۵�hn���x�������c��
�v�p�s�����w���~��4���eaq3�����)��bjll<V��ei~~^� �R��G��۷�xt@����Щ�I͝;k̠�J���jhh8v�kkk�w��nw�Ϝ�{Oo�χ���,Q�ȈVN�V��:�eYr:��z����;v���n��޽+�˕�3}C�����$�8����U�̬�ΝS�P�4�HhyyY�hT����n��"Ӆ�$]��[���'�e8��7'��U�h)C��P(���%����X*�������"���~�]�-.���T�������(V�~�J��p8���p��m�2u���a���쁀�P��ZR�I�  2IDATQ.g�=��/�á���c�L��522���Q%3��V����Q+k�@�$����,i�t��3�`�a��Cq�\�H$411�����J�Q���H�Ai4���a��:�`]��3.�KN�S����.n�����ݻ�5JR���~���TJ�5�H��Qq*����������X,v�._S��fff400�@ ��s�s�z��wU��g �_���:gg���gN�6[�.//���\Ն�\�r�t�����d�r-���������#�*B!���j�t������0����6�:�ᰆ��455����fYz��� "{,�������h�L8��⢒ɤ���r>)/�hppP�Y��޸�W?�TE�3 �L�߯��	-��(������Ʊ�|����L�@��TJ/}������#��Z��U���b_��CD*������Rmmm�wʳ,K�w^o��5�9����Q�6�� ��,V�ȈV��̰	ZXX86�3�HD����vt�o��ǟ��Mҩ�)'Z��6&�%	9mll���^vCrp.�,KKKK�{��ɾkN����~�B �L����6�Z��e8�M&�Z[[���96�Jǎ�I�����;�ui�G��DB���Ԥ����D�Q---)�����X�m�b���C����}�����Y��-��I���&/_����R|�ž�nשS�t���;lH�RZZZ���L�j��f���k�����d�82��J}���[����~���^===jii9�������Ԕ<;t}h�_���_��Sx2ɒ����5�ܳ�~���Z���jkk˹�H$���---e���@P?��u�����Bg����/����Pj�����R�>}Z]]]9���5�,..fL6�~���NMM���/-յ���ԥ��~���F}}}jiiɹ�K8�������2vǓ�j�O�x��P�8T����?�S�'Nd���fSKK�z{{U[[{��ۙeYZYY���̶�I��NV�|�)��C�**�����_|������R������ȹ�J4����=g)�����P]G8: +�]�����kޖ��"uvv���GG8��Y����UMOO˿�}Ϲ{��ʧS	�O�C�jk���?��А�36�M���������jN�S����&�H���1���U��� ���կ�����n�����:u�T���E"���iqq1c�<i���O?����Ǝpt $܁}�57�����lsI"I������RWWW�[�$�I-..jffF���Yf�i��uk��1i3ȣ��W���Y�8�,K.�kW6���7�̗_Q8D�.��o�Vl���/`��I
��o&I���z�>T]f��X=yR_�������ݮ��n�:u*�����fggw5Ǵ����|@"p�ƞ������%%�~���J���joo�z�X ��̌VVVv�W��������m� 88q�]7�~K�/�����f����a�����L&����caI�G�z���74|D�0������K�K�����ӣ��ά'���a�����+I�����jc�F���UU����]�}��~�f����C===���:�љ�R)9MOO+n�Y{4��?�D}�CG4: ��2]���j���m?g����ڪ����'�n%����hc�5Iq2�?�L��uD��c��v}���!�g)%%%���Io/����%���T�C���A�;p %%����4��;��l6555���C---Gv�iY��n�VVV����m�ٖ��Q���'�l��9;�u������m�ϖ�����M��!�� -//kyyy��I�s���ǟ���H�t�ok��g����v�������H;��VWW���,�׻������k]��[�v$p����ؕ+�V2�6�D'N�P{{�ZZZ�,�&�keeE+++;&�I�=��k�t��7$�Y�=Ѭ����N��Y�ݮ��v�������F�ik^Y^^������eѨ���:���8r3���替޶"���Juvv���M���G0���[�׫��e�������svV�}��jw���kku��4�̎�-..~x^���pd�y�D�s����J	]�~CW�_gd�e�i���u�g?۱h�$���=\�eeT�ϧ��%9�wQ��}nN������#��M\���~�K�w�ǩ��}x�r����pws�ܼ��������#�Lbee���74�쳲r4nn���ŉ��ܸ��?ڦ���E�;p��'�u㭷��ݵ�����E���jjj:�6r�XL�G�GN�S�HdW_W����O>���������4��s������ABUU������ب��F��Pq/�������x�r�vl7��$����u��7l�,�>^���W
������+=�H�U��n��n�\.׎Y�[zFG��S����v򤮿��ܭ�����nd�r�d�e)<�c�n��[�G�������]�8D6��/]����|�6�@[k����� ����@��W,K��Cz�/�8dY��Lw�S?����J����=\�t`ꓞ�Vz�w���@�͟9��yS�]&ٕ�����EMMMjhh8�@�`0�ȼ����k��^��S�x�J�Pu�����4u�®>�UT���I�����Eb�^$	y�^y<���)
���*A���g�&�ȲhE����=���]�m�Q�bZjjjtO�L&�+N�S�]��lx��]�H�r���]��~KΎ�]}���D���癃.2�u��uG��{�S��z�ӿ�f�� ��A��4y颾����e�ؖ��
544��������+Z��H$�`0��������M��F��t�]�yS��9+\]���sM^����Xi� ���N��ժ��z�����m"~<ǄB!�A��~����:HL�l��ӣ�z��/h�dY��Lw~�<���{X��l���U]]�#k��$�%�ɇ�H(������U�kp���g��)�\e��������: uKEE������D;����G�C�`P^�wW��~���ҋ��S��{�: �+Z^��?C�W�*�����=��ڥ����h'�D��%(���*��i���^����>����p�<--���_k���=}]qq������l�-;�+�e=<S���|�=�ߖ$z��-=��5��q/��$�v��5����{X��l���yxf[YY��e���T*���x<{>g��x���_�{llO_�h-�>�o~�<'N���JKK�o�]***vU���獍�|�=�'�z��=�嗬]������߼����=}��nWCC�����_���v5�D��G�E>�o���E�����?���`pOcp4,�Mc�<�;?��B�U{�����;����]�m�1�@@���{>˭�x��_�{���+pI��X�/������а��e��U\\��OQQ���R�����Ğ��+�u��u��T��pl��u���4~�Ҟ�<L���T\\������(�H(�L>���TJ��t��u58]��^ V��Z�/���g�U��􉿏�fSII�#k�T*�d2�p>I$�k�ág�]S�ظlT����ݮ�g����/�kD&[���#�=�~5;���`]���Ʈ^�S���攭??^�l�[��viY\��k��55E�B ���<�{�����>i�UKJJ9_ٚK�{v+I�hT�����o�����~�E=x�y�vف���k��9��k�d2��}P�ӥ�ׯ���UO���f��ٳ���kru���[m�-[�-**zd/���KI<������7U���iK�����kZ�������|b��UTT�H<K2��u�d��dRgu��u:� �D��DcW�j��������ۺ�.))�eY�7��F�SW�]W��# ���TQ��/����/��ښ��<�����[�u���	l��`M�_yE�/)��J�G������.߸�ZZ79-RY��_��3�(\��L�CeYj�_Х�7	��dq�Ư\���/h��9��y�fYj��ӥo��)��X	UWi��5v劢��$sTl����]�qS�����=p������h��9%�YD� U��z��]]������l�.E�����4��s
UWg{8�hY\��o�!�8��z5��Z���w��A��t��=]��[U�B��=p�:��W_�B_��=t?leѨ����7ߨjc#���REE��|YC/� OKK���/����]��;u��sG�(܁#�ii���K��x1k��e��zFF�74���0�<�,.���3��tI}}����$�R)���R�а���T�Ϫ� �V��H�}}��tQ�g��2�~Ի\�R�а�ש��WG�&.^���YK�it:�70���a.E�c.Y\��3��tI��Y�IR�����?<�J�?+c p0���>^��/i��3+c�ѨN���o`Pss��ǘUT���Ӛ�xIsO�S�n��8j�^��hX�OV� �p��5q�&/_���1+c(���=>���!���VUO�c-T]���5q�R�Q��I���T����&'U�}3�7<����|IS.d-n���R����s�Y`i��i-��i��[��Y�xYR�����Y���V������C�Y rC��R�g�j��[+=�usP
�mnN3�:=6��`��~��++�ܹsZ���r���#E���WV�13���1�X^9�� 7�����ۣ��^-uw�{�{��dR-�Kj��S�����C�9 �+RQ����i��i�tw+|�k���%u�����WW�gȞ��͝9����rtu)VVvh?�ƻ���Yu�̪k|\%�^@n���j��-��
���ϲ�Rjr��snV]�j]X8�� w�uth��-ww��٩�!V`��>;���i����)�S��͝;����Z��<ԢH塐����1=�ޑ:Xyn+nn��G���r���я�rOML����� �� w D**�8ݭ�S��kl���I���'j�T���V�ǣ��%��Ϊ��3�����H�9!_S�֛������)�T�v���V�ө��Y5:��k
���I˧O���&_S�|��
WV����R����#��j���(p��J�tu��١��&�76��ظ����DBu���P�˥օE�.,$�M��͵���M��͵K��b�ߪ(�R����].58]j��S�����+@A����lk���[��M�V�O0�T�|��xT�v�yš��9*���Р���r�w�״9������ʖJ�ڷ�z�[�.����67�2�Y��/-���VOu����e�	�Y$�,V�ǣ�������C5�\�()��ɓrtwi���}���Q�'�W��ν�'jZYQ�ܜ���^�hy���Z�ؼ#�55n�]�8�'����̥��R��g��1G�;������56*P_��ݮXy�b�eJ��e�$UY$*{<��hL����n-�Z��L�����+VV�xi������U������4�=U�׫r���H��B��&���/-U�^�XY��e�*J$d��d��T��$SͺO�^���&`REE�74(PS��k�xi����*JY��6�D%�����P���E��"���k��J��뗲R���U�H�$�yβ9�DU�]W����R�l@�
WVj���uJ�b�e���J���4��*��d��T
����R@FѲ�͵JM��b/ݜWJ�T�Jm���hT��S��C�^ ��**���^�J�K�(Wܾy/�,)�=yd�R���VE(���QVQ�uu�54(^��~臻�Di�J#����xL���j=U�:�c UT�@}���J���r�e�*�6�J���1Uol�z�;" ��                �	{�A                �! �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��                9� w                @N �                �p                ��              ��v�X    `���4vG ,�           ,�           ,�           ,��z�{>
=    IEND�B`�PK
     �9s[T��T$  T$  /   images/8ade0660-1c92-4b58-a3e7-adda420d3982.png�PNG

   IHDR   d  6   ��7   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #�IDATx��	|U՝���-�CBB$� [E(T�E֪�uԪm�Ng\:U�^�m�ڙV������� (*����,��@BHH ��{�����}/yyy{xd���9�r߹�����}{����&N�:<�����@Z�W������@�p&�i���4-��e�xd�=���4-��v���3	ߗ*�P ڔ�Я�
槟���#=�ȑ0w��Ćb@N�!C`n�����π6b8���- �W ��/g���sxg��eX�����d�&]6�;����}�2�~�+�K�v�z�r�n���~>�7��φ}����g07m���a�t���8�O���ۣ�B�:_�N�N�l6�Ax�8����>���؂�5G$�������6��5+u%���u�jBn�1�OF<�������:�s�(G�����������c���|�& �:�@DB��6Rc�l,�9��
D��y}���,�iM������gb�r���h���r�w��5�1��-!aY6��5������r�YGZ0��0h�ՊSʊ(3ه��ro�[M� 9*+PDn<��h���iN,��*�?���>��z?����]��n�ױ����no� k*
�t�Dx�-v��AzN��a�~ݴS/`0���$"�����I����#)g�^�p�15�˼{��o�𿗡�r��^�
�}���K�����F����d�j��r���^"���d��)=p���;qJ'C�2���<8ݞ�)�����8�^cߐ�[�J����e*��e\%<NG���}Q����]5��R��q����G�?���8��r�������݇�w��tת�c+ҧ,h�$�J�r�E�)�����3�=LTE��ܥ��_��>��jP�ź`��۰R�r#qi,��O�Tپg�2|�C�&��z,7%�V 䣺�h~����d��YM�pST]Q��zI[f�D��W�\��5� ���8�ꊢ�M_6�g��	�O���օ~�<dKk�7�j����=4���f��$4PVP���]F��}�D6�<�Ο�(w�J��>���8�f3����;�wj�"�+b�E�2���>8�v��\Q�q�=��;M�u�M��3]���zA��P��P)�*ˠ0�ĳG��hc��ѭX�B�3���M�"
�Ѐ��p�	�O��Cqj/�q}�ZВ��$ퟨ	��r�42���U�QT� _Eng$9�|�/-%?�:�����#�1��*���a�܄�<�Fw56�1�g��>�,}�O9�1\0t�^�BO����#�>���*z9�L"��p��yVq3�`?AP����D�{8���"g������	�9��*�␙����H�f��"��&,݌��G^�NsrN�P�Ɔ�����%�2q�&����J�1�vN�.�M��e�Q��F<7� �B�ǒ�:���e�vD.񒻗��p~��k"����2����E�����ĝ=g1�-Esvz&�'ʷDz�[*4�r��b�!�*�mT�؊���w�(z`�=��j����W�PC!��!e;kE'A���㨮
��{�>��
�P ;�m@�
�­3.�΍uC�<چS�n�.hVN��i����{��e�k6��F|�{�\tUl���9'	ܪZ�$d.ڗ  �ȵn��g[��^��5��zmZw?�
���)��c�X��+i��w|�
�0�6cV��j�C
�9��P G�:5����Āa`�$�<���p�˺���&���ߛA�y���Y#�ћ�\�u�W��ć�� ���)�Ǖ�h���}�������De�ڟz
��"�r� 	���a2�8G����7F�ũ�m�C��Kf�oC���N�x��P� z�a=�� ^]�����H��"�7�	�+Qo^���/~c�<�;���G9�����BT��k`��
̚+W���\4;��7����⺠��ְpC�%7��&CO��nEp�j|dL�� ���Ϯ:Dӡ�v����=B}�����- ÇC��zo�s���EV0Ԁ(i�'C���0^x�?�G���
���	�lX��*$�����p~B�p���ܯ�7t���9�\IO_�5�����5a��o�$��g���_��w�����Hu���������q.�C�������ʏɽa�sҹ�Ƕ��0����_��7P/uz��T�e�cF�[5yy�&L��⋩9a�'�����J���^/M9�Њ��gq�������y��qC	�T������D�|X�ʨ��wF��"�n��C6ޱc0����;0-� ���\��J�F�~��|�CЇا�?��9��v�i�z*��
�C����xtw2�Z�#�}J����_a��U���o��m_E�-(+̠b�x�䧈GlJپ�o��'`��u�>�U)��~>���S
��}�����r*�2a+)0�����w��K���+���u��mj���v7�X���#'��>\���ד{<ڃ��_B���M�>\� ��AFD�a�ou�~�s�.�E*���^�n���n���o���wÍd�v�W\m`9|>d�6xh��i]�ǘ�|��H��$[���Jr�$�z�b�0��`�FU�	*n)�P��k8��.�3.�N��J."��DE�**�9�S�r�b������E�9�!ٱ!���οC����wo�8�B�E�?�V�*Q�乨���z!�i��x�.��L��Z��=�N�FTd�?�!̃a.[.���x�m۬�:��4k����/�c�R���q�$��ĭ�S:�H��.r��E�D9����9B;�\�������*x#�L7}o._ai�N9q�T�ӛ0^��\x�e�[<��'U�[o�J�\���p.�z����}ݞ���ˁ{��3|)\x���0nQ�����3tf��+�g$�G8�jQ���ʋ���)��h�GA@����j�����1�J�+��8�P�XC���dq�����o��gx��=�g��=��X�z��0�A} ��LW�ܶ>��I���0�y'~#$�OY�fZ)=�{�^�;�kz?���?��e��+)x�W��rG�����վڂ:���'#�R�F�ܑ=d.�'M��\ı�+a����.�.�@�F�Ӏ�-�$F�c��p���9)�,�AP���rEsN����i�=-v:��Hw�C�R	�}X�������=�B��Y���g���xQ�E碽��m��pa��k����� y֊ǖ�����n��(�)��@bcT_gqg��z^�2���`�mx)���#l\%��@��7�Z�Wac'����'�ieC�Ŧ��HOG^j!܂�1����pC�a{L!Pxl�]�V%tR��o�m-p��'�]���I��F�`�蜬�4���X���q2�W��& �e%��hkA/Ž`�]L��c
a��|;��-��*M�����}��I����7W�寄U�Ś�9������Wp������\�?G�Ԣ�t l�I�[l��?�{�k�=
�%<9���-�ݼJ���;<(��~x	@��de�@?\Ӟ�L��w&�xW��J�'�{ �����
aA�[����3,i�౭x���ԓ��,Jv�"X��zS�<�;��~��g#ѫ�L`Q27&$(���
�_����0KaU��g�9X<����9��l��:хt�٧έ�� �����%�@ �+����+ZQ���0׭������"I��N�N�3R?�*��m�t��71O���0x%��w�E�Qh�Ӿ�
<�g�̇k���-�0��w��w$݄�[G�u����%�L��Ze�8hF��q��u+��ˡ�v��,���ef¬?���eg�1�k�Y���
���R,��"�7�Y�ۛ"�,S�İ��Z�J�^;��V�v�b?��i�X�h�m�Ǎ�Ͽ���y~^�ޱƎ��f̀>s�8���Zo�G���Mo�|�$)6��J�}�Z2Ĺ�O��΃���k�_���^7�E�O��F���/1���:>������֥�m��1jo�k��X뽸��U����3���쯂>v,������:*���ll9H۵�r�*��7���F�FP���Ӯ�)�����n��\�%`�(�?	ۏ��\�&���L*���β�����#���~��3a,]B��50֮=.K�N ���U�gn�w'��f�
�{pN�����R8gk`(�(#�*��	��е$�sU��/�8��~�[���YsK�V��[t�L��g9NKi��9W���:�W�l���k))��	?FKNr��PXUm���A���J)],X�Z����3lZ
���3��/G��7V������� 	�Ny����ϥ\�S���/��.)��v�,���oʹ�>�}�|j�D��c2��P鿎��Q��K}�(#�ňǡy�)h�N���p44 Y�Jt�MHq����/e@�`�E�+#]��z�ɔymj��V璡^Jw!M�d��/��{�>lmj�k9ٝ�4����lw�]���T�QN�\\�UcO��r.NSL��K	��L^�Ά���x�D?�ad�Y�����JX)	�_M�|��?a���y���\��Q�?�v�j��+σ��Bk<"@}�N�'�47��4��|�ƻ�����_�6�¸�o��1(�{p�;/'�yy*'���\�B�p"IO)r�b��*m�������d�w�1��);�������1�������fvՅ}�0��XKR��R%���b��Q$�"a��'����R��:�R
���|"�?%��)P�Ǜ������D��3�7��R %��(�58���(u�3 o�����V����CƢ�f��<aR�ߨ"T��Q��gN�]����dV*� �Ann��&������7�R-��6|/�q��_s���h��s���1L^�L��
�VQ�ӁӦ�C��d	���(�H5]g_�='g���B���B?�/�"��	�A��5^ܜe�'l�a�r��G<���jP����:b�;�<���>�;t(����}��β�����q8����.'f~��m�с��k֠��ݝ�c��Z{>;�DCĎ�����Q�6(��/����9�N�H�V`Z�?
_��Tx�8魭��;қ[�A9-�6#Swl��,P�k�e�p]��]��1��}	n P8����?!Y�y9��/�~�-�I�7ˆˢ�Y��`l��,R7��{_���s�ަ����[Hi��=��	>�+��⎌�#zO�8T
�I�~@o��	�H�s``�"���JH���"(E�	OkUorH�"�2�{�4(ERҶIHPq��G���O��#������������<95�i,,�$zri�9�Ϯ�:��#�������\�u�������1�K�`�hI�7�$�,�Hg�o�w�� qk��x9��gށŇ���Ň�
 �䒸�����i.�����~l��+�ˑz��{�n�=Ԁw�r�-��H�A�C����ᩨ?|��O2������m4�6�=|!(Q�����k|4D�M�Kfq׀��֯�ńH�R��GB)Q�)�(b�t4(a���(��3N�R�ˆ||����HPz 	��C �}Y�V��MlC�%C���t���|0f��QJVܙf�v�hg(�N !0��dn����C�^�mʶe(b/b0{�B��Wd� ̳�t��ǒ���hXq�b �=�����@�x�m̶���ً�"���2|����;�ۚm��񑊝@���g+��-�9۞�Rlg <6�����m��%�=3�����P������@y��z���Q�ٰc�q-\����<���^�x��������y�_۾4�J���)�B�*w�wT%a��ŉW�{<"N��%H&N���wc��6�%:�i�s�@L
�f�7�<k���N��/Q����޻W3^i�������r�N?hkGڢE(^� �DS9�i�4���C߾�/���ݻ�%wFj����&	 �+P�ƛp��	-+�@ða8r��0++�C����(\�&���p��:�_q6BV}���/�����.#����ƍ�՜q&p��޷�[�d���>h�&�¶�\T?�\'Bkmk�ݓ�FUY���=~�(�C�I�"N�g������6v��v����{D�	6:K��.V�;���a�y>ũ��d��I���d؁�?�#�������9�a�H�����,.��>�i�ٚ�9޻�A�{�Y?�G����>Z���Vu�ٲ[)E�]{/���߻������C��/�b����ҳ��n/~���ƞ��k�U}�
���f�9a�����ٳ����<x�п8��ӎ���|��`��^Ɨ�������Z6� K����kŞ�����O�z������A����+��o�w�S�q�$dnڄ�;:�$R4���<����ݻ�������C�<�1s�#���zIa;��OqJ㟓�C��W]gQ�����Ν;PVvq�A�4��:�Mvuq��>�Pj;x����0��o�%�/r������VX���G�N�>������MvA�eڰa:��T�`۲�Q��Cp�����8yo �>Bl�nll�[�~�>hooG}]�J�s;�����֙�tO�7���O@w�p��Q>g�8�����`�okn�?eʔ{��׽s�̹��[n��>tX���9�;�xg큻�}�t4o��O���z�~��a�Q�75��������&���myA�K�À?��䷞r���q�ŗ0衇D�%6�9ZC���u���[^^^;���|l�ƍפ���tS�Nۿ�[�S�w���cp%�E��0}o�!�9��?���C�����/����ԍ�a`6"�����������#+κ:�W>yCe�a��?==��.��E�ͽvݺ����G�v����T�:�+�_��uޮp�F[.W�ܹsϞ1c�2��5��t��o��8L�\)��q���A��Cq������V��'>��C����j��ի��^��lq���/����N)�M��}$.��k�s����3G�1���k��6��1c��dC?�>�\�3�����2�TU��������M?~ŧ�~����|"o�ɚ;O���!6��7|���i����������-,�ֻ���#��t������ys��]JiX�hB�y� tj�W\�6l�[[�l�H���d<[�ܹ���@����{ZM[?\
/w�rTSC {���������_�\PZ:���v�P.��@0��E��3:���K@2(����1pР�6n��/�F��Ȧb㕿#�seHŞT+K'����=�]N�͜Y�a��������!��[��6�pݐGEFU���e��ӱr%J��uD�{58N��|
UT49g��NKO?�C�����(^�,F�йT��=��;�@�}�!����5��Z�}��T�l���J���Q���Ʌ����������ʞyF$�Н�Ia�ePV�y�M4�>��`_U5�����w���,�t�e��|��T�sE��`!�)�����N�@.5MgRC���;p }翝T�
>ۀ������Ta�o���T������;o�~p�ee�얂�߀��y�H��p�gwXE��%p��$��K���l�O���ԫ.Kb[�(*��&�8�(�8�s~�^w���('ѝ�cY�	z=�qb8��|ͤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�ɤ�H&D2) �I�L
�dR@$�"�RDK�Ǹ��B���Y��_���|��@t���`����h�_���;Df��-�{�6q�f��L'�Ό'�[x,kw��ķ[���̦w>3rx���?~����n��la�PX �ݱ�K�sD<do�!^�[ �`������@۾��vq����jh�Q]�10֯���Ѯ���0`۶�����v����v�܁&�zZ�۶A3��qb?55���A�� (ގ�6+Qt��GKL
�[Y	�}p���x۠�χ��_��׵?���`A'�v���p�o�.+��[Æ��t�߼y�?t���>�A׺��f���o���+��j5l0�@iǎ��׷�������'p�A{D�^�����~�8	p�ƍ0�_���R�7��+�0q�C@�o�%Z�E�j��v���?� -B��-ȠD'�߂8|���@��5=l`��ȡ8'wY�?�ZH)�ރ�{��>���Y��׋~�wF.���y�R�(NᲵ G�(�R�I/."iU�λ"'��芖��U��{8�pE$=?�rk�Ĉq�k>s�[�?�+�tʹ��.�j�%���aC���)�����W�o(B#$N%�Go�HDH�~8w�\�Ë#N|�8q�+�xm!%�� ��?��A�    IEND�B`�PK
     �9s[��r�  �  /   images/022fab5a-d187-48c2-96d7-20ad2a5d1671.png�PNG

   IHDR  �   �   
VS
   	pHYs  \F  \F�CA  cIDATx���ylTe��񧥅��E��Ũ�W��+"����K��Ƹ�5�ܪx}��z�AM4z5��B"�DAcQ$���EEJY
]�=�c��t�zf�s�sf��$��az�<g&�g/3���m�q����S (o~(o2Q��P�dJry#	`  �9  `   � p�  �  `   � p�  �  `   � p�  ��D�y��)))�WSS��$Pmm턖��;l��&���&�M�D���N�~L�.�Z������{a֬YM.��̙3K���/�~��w;�{^֎My)o�(/��WW+o�iFx�d��ի�޷�'�����1c��8��w�*�ż���ƻ��(/���-��ZS(�r�w��֭�yߺ���s��_�<����nhh��w�[��7񢼔�*�+�[���l���-ee�����������y�i�̆��ݻ������:��۷�xo(�奼aQ^w(oq����n�y�������{��޽{�BTZZj?�p3d��e��z�j+�9r�8p�IZ�奼����@y����җ�2}�(� N�1h� kǳy�(P�p(o�P�p(oaڵk�)S5����y�  ]ASS��|^������6u  �={�e�?�����   �Ai~ ��4.�Nm  �LY����DWTT  5?+s�u��#�
��~��q48̅7�|3����Fy�Ay;Gy�Cy�᪼��ωn`�ۢ&�B����㓆��}|�P^��O�k��Qk7��m����t���   �T9M�B���j�0  �i�t�~�>}�  `W����V�(��  H2�f��JZՂ+++�Z� �bSWW�u_V k0V��b  I��Uښ p�  �  `   � p�  �  `   � p�  �  `   � p�  �  `   � p�  �  `   � p�  �  `   � p�  �  
2�{��m�8��k�.�z�js��g���#�4Ç7��S__o6n�h֭[gZZZr����sꩧ�ϧ���ذ{�n��n߾=���ٳ�5j�0`@��777�m۶��>���ٳ'�c8п.zN�ijj2[�l1�6m�@�
.����o}�Qs�A��^�b�y���<�1cƘ3f�nݺY;�����ܹs�o������z���s�5��ݻ��y���� t���7����O=��Y�lYNw�'�9s��ݻ��wk֬1�?��ٰa���\ O�8�5|e�ر~��~���\v�eV�W�?�x?�o��6����>}�D��@�2e�����x})��RUUen��v��\Bx���9���v�ifĈ��3˗/7 ���}�f�ׯ_?'U��!�b������z|{��&]ߠ�l�n���\�2pst��R^^n�O�n���̧�~j ����$y���=��c���_F��p�|��G���/7Gq��c�&|�)���A,]�Ԍ9�TVV�}�iӦ���o4 t� aժU��o4Æ�W]uUƠ%4�158(�Kε�T���͵�^k��~?�|*C���ǏϸOc ��5�馛�Ar=z����r�-�ٱc�Y�h�ߕp��G�	&dbSw���� �� I#fm���袋�F+0�y�f��[o��w|p� ����&���6�s�Q���^�߶`�lӯ�֭[�ԩS3� ~���Q� `KV �����d�s�f�{��[!�p�B �d��j����4�TMwQ�qI���臰�}ӥj��{ 6d%kj� U릦;-4���E��z�7��W�]�����` ��� N�fi-Ƞ�BXF1��j������3��K���Ԃؐs�}����� 3PH*�R-��Cm�O��K/��,X�� @Xyu��i�v�ի}�	���c�����W��4�K�ඣ�'M�d^}�Uj� B���k�D-t���HmV����;��ˍv�a�����|�� �a��ڰ�X�.��aK{�8�0I>t�_|�_�;��_쯂��= �+#���/E��;w��W?b�V��u���j�z��I�x\y����)��=�u� ȇ��[�4�X��tŚ���w��v$L?������/���J�5��P��y�gN>����~�q�{Z�]-��N+t� °>z*ª	w�>����W\�1b6,�4�t����~��6Asݵ���c}1�={v^���i�^--�?��_SZ�&E{����� �+���
���>�b�����m�ڵ9=^s�/^��Z�v k S�������~ڸ�k��?�c�=��>M������ @>"�?���T�U�:묳"	_}�)���amذ����O��p[���2XM��Ԉ�0�RT��u��ĉ�S������3��O>1�ƍu�#F��$����ƅA�e��\` ad$�6`H��X5��a��۷�)F������݆O}�6m2˗/���-&���m�Gp�Z�9���c:홬�����СC�j�ڶ��Z1 �a�T��ԇ�>�4�(� V�h��F�����y衇�}���-(r�3gNF`+��;�8���_�8]p�Y�}��� ��6��Q_��4���)�MJJX��|��W��DZ{9ݐ!Cb`�lo���)H �
�9��Ԡ*M�� �\�֎�w�,��͛7g��{H��m�0���o�5 FΣ�R�aM�E��Z0���կ��d���/ +��ɪkQ�\jª+���/ũ�����oV�Ze  ����&�2��� F!д#-7ٖj�6��@�	��9�A��h�F
�Y��ꫯ��ib�~`K�240K��V�s1���§���sN���-b�g ք`�fUS�O+���:ujV+�ւ^�r� [�������<b .Gy�;vl�������&+��BЭ��T�>��k�k��H�����j�+V ���.	
Ԡ5�<}���i�_~1.4�|�M��P��y�P�C�F+==�����qҨ_�)֘1c��ɓM�~�B���*�\^g��h*љg��a�����5�����q��y���6��y���Y�z��������>}��8ai������{���E���Ԅ^�⨣�2w�}wd#�7n���Z�R�ng�ٺu�rZ� ����|p'�6Q]]�o��f��OŜt�I�5�k��a�:|��硫U�j}�\Z(��|�n�G1�~D�I 'u!��5�3	��p�ש���j�6�Ɩ-[�ܹss�&Z����O��|z<���y 
�8I�Q���~_���۝>��_�ޯy�I�~�s�4i��ի��v���%K�>�j�꿞2eJ�}��z=�����s��K/���5�_:�3zOn۶�����fٲe���q�;�k�`}H����Aj�:G�ӑ�x�	���]w�)&
`��R`��Q���~� @Ym�f�#  ��  �p{�';B  �:��"� ]�� ���A� ����fAk�
_ ��Y	������%| �������~<�  `!�{����	`  B��7���� ��w k�sG{�v��/  �+���m���"� �S������τ/  	�
\mX�K�o
�_  2�m +xU��\�|w;R�2� ����
Z��U�7�6�����d  �_2X���]--iko���F  2e�B7�>ގ(|iz  [F �\(C��� �}l+0�4= �1�5`����  ��Y`j�  c-��|M� L�>`�r�<_\ \�B
Ԡs�S�l��   ��
`����LjmgV�  ?�ր;�jnf�  ��n��T��� ��vk���W�g誆��}����'��� (Y���D郰����ҥ״������iLZ�Z;4�]5  I�����U�TM���>��a=N7m�� .--5  "g��ٳ'�)LZ�R_���a @Ar�
�ݻw��[N���� ��X������]�c)���  *��}�����ci WEE� �P��QmU� ��,�� �"� �r�`�Z0 �P��QnW�c� �B[ ��9�]�R+v1 Pb�8����  Ik8�s� �B[ �4 �_�*��� (�p�H  
E�5`�Ϧ���M;8�� (���jU�~0
qm� ���Vyy��l���jzV� P(b`5����z-X+`�� ($��۪��~`[�B�x�Y PH�t�VVV���MMM���~_ �B�l�RUU��7����/� (TN���VS��Af���G�� PȜ��Q���hm)��m�X�R�c� �$&����
aV� ��p[/ ��%6� (f0  �  8@  �  �0  �  8@  �  �0  d�m��݉  ���O���
��;w�;  ;��A�~�2������  ˴ß�5}׿� ���7  �>Ur;�{�  `��gϞ��n���f�? �}j�VStj��� �Y��ݻ���466��x[M蕕�9=�����y)o�(o~(o�(o~�Zy���G݊�
��� ���{�}�jjj�g��٦P��P�d���������������  DL-�ܒ��?X�_�  ���U-�G�0�� �GF 3� �x�f���Wâ @�����b���0_|��]��>��$O"��M��-L��X������矛w�}�lݺ��q,X�/�=n�83j�(k��¢�vP^���#��͕�^58������Q�y�~����.^���(αc��t�R3~�����O�\�xw�7P^�(/���Qy�f�V�,3�{a�~<�=�'g̘�3�sN�6m����y�E��{�����8�My�Gy)oT(o�\�׆�`�~^ZZ�?�v�za֬YN�K��;�x?��9s��VWW_���/�>#�sQ��Q^�k�_��)�콰˼�8ϻ��LBxo0�?�jkk'x���9N�ql��奼����EY�($:��v�I�����y/��>oʛ,�7ʛ,�7y�  +  `   � p�  �  `   � p�  �  `   � p�  ���i��x+��    IEND�B`�PK
     �9s[6ah    /   images/39d025b2-988a-45cd-b457-87e73cc458ec.png�PNG

   IHDR   d   )   �$��   	pHYs  \F  \F�CA  �IDATx��[hG�Ǹ&�x��FATP�H�T�R��iT��!�>zA��ڂ�WERP�S
���/�A!Ѩ�&^� jLLb���g;ߗ|I^�����Μ��=g�3gv=������ͷ)��7�4æ{[�n5���L��ܦ>~�6�J&�Mr����L�h�݁8U�U3���7۷o�������+�&�c��7�|���bΞ=k�N�j&O�����K�)�Lyy��7o��ݻ�inn���3g�>��3��}����|��Y�`����A��B�}hǰ|o����{���	�=;�2%(--m3fL���2,z���M�oig<��Gj����O��ɦ3�AN�T9�6�j̰��6��Їr�?|��<���;M˼ϟ?���E������oߚ!C��d}dZI�1b����3)@X#G�4���.�"�v�mgPvFF��0@�YŬ��"tc���z���FCC����������!���ӧ"Gm�4�p���2�޽k�3#hC�����6��#d��{���"u�ŋ���:���m����MG�^�@�>�>lc�t����x,#�'�$zh����.��I�Ĩ�$�)$�K�θ���Ϻ���,;ϓ+�
��w��s=��>�~(s�d"�S����cǊ+k�a>�ĉ�p�Ǐe�	����gf͚e���������1c��}����Ҽz�J��2e���L���
�@� ���y�f	�\�zU68
�5i�$�z��`F�7������B���ev��!n"u�F�2�?6;w�W{Ŋf�С����Č�J���6o޼�q׮]2F�{��b��h��
UA��Nf��k�DP�ӧOf۶mf���" Vƽ{�̖-[��˗/7K�.�jۻw�����Ǐ7�w�6}����8qBVбc�̆��ŋ͹s��D���!��e�c���x�X�C00�v��P=�
V�NUoz&�\�u$��������K�.��y�x��0�p8p`�c'�̙c6n�(�H���G��p�ܹ#�k-��Ø0!���I쌄jS[�L��͛7ͦM�Ė=x�@Vl����a�f5�q�m<���O�<1�O�!��O�t������e�e_��0���� �ANN��K
�i	�Ǟ$�a���C��.�\U
���!�Fʸ�
�~�C� �� ���X�v��0�QM��n�:�S�_�N|ucg0�'�1S�j�*3}���K��7��hs��EqU]��̞6m��!T\bM(�6Lht߲r�J�DD>�>|8�U��sg-�A������Em�����`Piii������,�G�LYYYT�SW�l�Cm^4x\555��zK*5��G�� T�֭[�ƍQu��<���S=1l�ɓ'����K�V���x�����2���	Pu�Uf��0^G� ޘ�OcE&��v�3��!x�}��EԳI���S;��p���}I�g�i��UU* �B�ӓ�~xz��2aF�ՂZ#���3���6��aW��X9��l��{Ѯ���5x�D���@to��rVO����
Az��;��@zq��rl�"��z^G�lR=WAD��P�N=�v?щGw�B��B�������o����r���Dm���Lǥ�86����������2~Z�G�1�{��e�8T�?��;w�|���t�A/))�j<{�l�hѢ6��^�O~�E8?_�f��Pl(?�c�8�v��g�~p�k�D"yuuuK�Qii�WTT{ߒ���Mt�h�������TMMM��ͷVUUe���۾��ȍ��nԞ�����}P�Q�[�ϱ�]Z�8�^29��7؅�O���{{���;�[��������ۺBۦ�����U�Z��p�8]v��������4拐�ׯ������]�~b�gϞ���}��G�~�Џ�Qe$��b:�,����B�bl�1�v�����;�"�u�6�=B�4��r    IEND�B`�PK
     �9s[��9PN  PN  /   images/779eddd4-9cc6-4216-b155-89a4f50be07b.png�PNG

   IHDR  �  �   ����   	pHYs  �X  �X{�M   tEXtSoftware www.inkscape.org��<  M�IDATx���	�dw}��_��Φ��h$��.�B6a�x6/Jl�l�<�^�B�q|��>I�N��<'��/f�el���ZG�A#�H��=�=�{��FHH����u���Wսu������o�[�Z��j    s�%   �9'�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   ���Bqqy1~�7��b,*Fg1:��Z.P��`ԟ���6G1�F}ZU��h��q*�ϲ8�^
��Z��b�����b<^�����bl���U4���?-��qQ1�@�U�W\taԙ��ǣo��(�,]л敫��ؽ-���F�p���v-�z3���8u�^��ʝ:���h�m�tq��b�A���$$�I�x�,��|��.�ҀԳ���5?�����
��e�b����h���aC���=�.�z����4��{^����6�@q��b��"�w$!�I�x������b\�r�t.]=k.���E���ѱxE4�wFKGW�t�D45�WG��?��_�F���7�+��KQo�w=������&s�?�X���$�Ͷ?�X��o�Q\��_�ś�����c�T�����S1xt��{wL�6�:����Ew1�U�b;����E��0�:s�xA|Cq�_��]et/����n�%�o(}U@�*7 I����e��q�с��h:/��uY>FI�¥u��2Џ<~o~��8��!?����,�׋��'������sD�3'�������/��K�zm�~�ۊ8}4��  �Dy$������|%v��q��oF�:~f��p��۩����Q�z_�,�̺�E�W��ߊ�g^?=��9V��ָ�m?=�7  �Bs[G�z�['F������-����Q;�Hy���b���E�<`	tfM�"�V\������_q�b�{?���  ̖��FW�⿍K��x�ӿ��wgn*w$}��~�����E����ά(^���-/O���̼����ҟ�����  ̕r���_��8��]��+N�}�ro��b[�5E�o�1�N�/h7_-�s(_�ڷ���ˉ�� @ˮ�5n��x���]��3���b���E��PC��*^��/s�_�h.�� ����ƚ���y�����hk�DKS%�|����x�U� 4��$�W�ܯ��W\[��oN�T.N���b��]E�>�F:5S���Xq��j9�ֻ8���'b�E�O��-�h��;b�X��K�Z���w�S[cE�������G�����@�(��޳�x�?~0�O+g�;�>[n���5 Щ�����s��8/�������^�aJ?ga�W��)F�D��lk.���v��ŝ��폝� h7^7}����<���Un�~��ֽ���o�g��x�*�C�����W����OEǒ��3V��ŭ���+�Á�dP~�❗/��}sW��;� E�����~2��_��G����=���H�p	tΫⅪ<��k�(�R-Z{����s������K��U+�9�,ho��˺��� 4�r�Sy4�=����H�����ɏ�)�}W�>p�tη/cey���=����=�7��?�fUO��K������keO�@�Գfc\���{��1>:\�Z^����@缩T*?[\�ؙ�K���Xt�g�w��o۴t�s搝���q-������Ŗ?��3��^l��Z��π�@�s^/L��~�������������C������-`>x��I� ��]������<{������Ŷ�g�H�u/̘@�|��bL�o_�l�#�fA{K�����μ���p<y�T  ���?G�/�����6�/��̐@g��3X��.���GKgϤ����)~�q��q��h��#�� @kWolzϯ�ÿ�/����b��_U���3 �9�[|��Ηl�>V��Ó.�\��O]�"�u��8���ظ���&N���C'�v��Q'i N[��Ʈ��0�'=No���?0��T*늋Ww"6��#��y�+Ǻ��Ӻ���'1�~�T<�7�N��Ș0 `�ۼ��������3sn-���T����$Й����/��X�~�oZ�7�]0�;�؃y�10<  0�^ty,���q��o��g���9`�:�V�T����Lo|��O�|�uj?�邘|���=�o ���#� �t6����z释m��j�jÕi���/����`å�����t�[7,��������ϔ����}�  ��`Zp�8���r���?L�@g&~�̕5���I,����u�~h��X5������  �կyۙ@/}0:�$Й�J��Y\\<q��9V���I�/㼵��n/�����9  �êW�5�~�w�:6qd��b[��Z�L�@g�~:�|�ڦ�m���]��Z��������9O�  �틖��W�*�<q9Yn#���#`�:���3W�\z�nZ��-M��C��{v  �O�m��z��!Й��t]w����0�W��9�8^��Ҷ�  ����O~�w�LN�^�@g���knk���xم��{.Z�qN?��q��H@����O�eԛ����H*����z,��[#iz���okԛ�8�m���*'�L�@g�*��%���1�]+�G���F+{������v;�&�F��ãIODC���Xk���E��G�u�8��ZZ�k���߽}b��f^_�VwL�@g:^�J����.�fA�9������l�P  �|Un7�Ko(�'�@�3ן��u�@_��zN?�#�� ��ֽj��'�5	t�D�3K�\i_�t��bI����� 0�}߶�)�Lǂ3WZ:�&]����>~���  ��;��?� `�:�����5�%�ۚ�-�G���;  4���y�0E���<s��m�Pkm���)�  �����ON�'^�@gf*���  ���/3$�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�$s���طo_ԛ���h$���u�K�� � �������V���  �J�  @   �   ��@H���������z��֭���[�(�������@ԣ?���ŷ�7 ��K�$���]=�Qo::;��4����z,�� p�y�  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @ �{��F<�ukԛ���h$�=�P��G~5��������ܹ3����� �t�dN��M淓�����`�l�?.0w:   $ �Xz���C���hM�mQ�z/��P������ҟ�c�{>����+ �{ �JsK�v/�JS��X'��:& �&�   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@�����  @���T��X\p��Y���r   �L�SSO>��O�̮��  �F&Щ�{w�������旼}����G  ��	tjjpt<���}�VĒ�>܆Ǫ��O��  ��	tj���H|��q���X��#Z�*q``8��'�|�  �$Й��Չ /   /&�   �   	t   H@�  @   �   ��@gF=��<�/`�V���h��	N+�G��S��^�!�l�>����c���/G#Yq���wQԛ#O��vD�Xv�-ѱdep����{�_LU��'fB�3#;��t�t\p��yNo�}�7�Q���'�2��i��XZ�Ჺ�=w����b4��>�	��<�Ǐ4�s�A�  @��x������W�aV�ҷ;*��;v,������T*�~_�Gw��b��=��.޼)�����.� ��o�F�v�����[��s��c�Ν�(�-[���Qo��������K�.�j��.\3��y࡯�����S$Й�g��;c�5o��;m�uT4E�yQ����?�ѶǶ�s�a��y��'�m���֮���Xz橧*З,Y���Qo����9(�8�r������Kc|�������,�ـ)�   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   ��t,�cO=8�wZ9�3*ǏF�|�t�Z����͘��m��7���x2{w�Fr���\���wk$'N����Ѩ7CCC�ٍ���Q�_�ZulgT�g7{�m�²�)�Lǥ#�N��_�d0��@�/��?���o?81�߶?�ub0��ٳ'h\'O���۷�Y��;�4`�:   $ Й��7�)����������ϣ�?�s�(\tYԣ��Kj=��߹-��h�]��{���Q��\��8ypW��o�K�3#k^�㱬؈f�{Նx�~)��:/����n�4���E��L����.Й�   	t   H@�  @   �   ��@  �:��R�K.���:������c���14:   tf��xϕ�cuo���������ç  2�VǣR�f�Tf�@��Z�+�׬��]�/����)�{Պ����Ğ�  s�:6cÃ�^jjj�����ӛjM�SSׯ�}�8?�����%�o�  �K���"�Oq^}n���XT�NEKGw@�	tjj�Ү�.s��h+J}x�  0W�GG^�g��^�Y�47Ԓ@��z���"V~����%��	  �3՗?�q�ZztjK�SSM�xR��   �@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �NM�����  �f*��n�5�NM�>>�z�&]�oh,��  �R�����ȋ��^in�5�NMݳ�x�juo4O��o<��  �������}a�7����Pk��:00w<q(~l��hz�Hx�@����  ���:����щ�J���"Щ�o���[7,���:��R���q���Pq���  dR��v�@gV��E���  ��&�   �   	t   H@�  @   �   ��@gFN<�5��=���E��&��:��F����OD�h_�<z�l�z3zj ��z$�WFKgwԛ��O�б��z��7GkϢറ��8�����6��PV�ȶ�|<`:n�wwD׊�ӎ=�h<���F��֟�+~�ףޜܿ3��w���5���X�Შ7;��S��/F���C��eW��6t�@�=��:   $ Й�}�mW/���ٽׁ�Q9u,M�:u��J����b>z�[ߎ#��[�n]\r馨7}G��C�=�b��q�UWF=z��G����(-Z���Qo��������.�j碈�e�z�G����ľ�)�LǶ���^��w��6�?*�F��Ͼ(������>��S���K��"����fۖ�*�7\|�}�������4T��X�"z{{��<��3�tvv���������_{�������@�0E   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ Й����h�<���iS�᨜<�fdd�E�vn*棓����x_߼]ǓٿgO4�����\���wk$CCC����ftt48���1�_�\�؆����r[��0E��vx�Xl��f���x��G~5�_��������塇'�ߎ;�����[�l	�r���\��S$�   �Ό,�tm�/\0U��]���/Z+o|S4�]���{AC��R�;ף�1�r�qk._����=�ў˜C}����oL�@gF6���c�U�03.��|���[ײ��c����4��EK=����=�̀@  �:   $ �   �   	t   H@�  @�Y��T�=m�\�����qjd<   8M�Ss�b�nâx����ib^����/m;'G�  ��	tj��-��Wv�`^�W��U����=���t  r�Vcld8���6k�_Kk4f�@��6-�zQ�?�]-�ƍ�㎭�  �T�C'�8?��<�3�Ǌ�hn��5�NM]����\��'�rۑ�V  �����sq���#�������Z���Ү���\�����  �+/�߻mL�Ss��*��~>� ���hOjO�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@���ƫ�u9  ���Z����S#���u�e�Ǫqbh,  `.U��"�^��Z���C{�c�ҮI�y��@�U�A `n5�����hT���7��t�C�	tj��''����/y��������  s�R��������Ĭ2��p�� Щ�r���;GN�ƫ�-�֦�s�:wl=�o  �"қ�ڋ+��M�Ss��j������buo{4�~``���  �G�3kʓ��86   ��@  �:   $ �   �   	t   H@�  @�y��Oǁ�.`�^���K���w=;��S�X��kb�k4���ά��� ��?���`Uԛ�w�Ƕ=�b�m���?���'�j�Ⱦ��������0��v��<��7�g���h��Ѻ��Gj=�ֽ�'�2Џ>q���(�_�z��<����� �   ��t<�ڵ������Y����mQ9�L4���ѣG���T*�˿�/c>��������`r���x�[��f��g�}�S�(6]qy��;���K��|l}��h�֭���Ψ7�cǎ����5k��WuхQ]��Y�ϝ�'1r�)�L�Ѧ���]�iVﴩz"*㍷!������2�/��ʘ��\� 8�%,���x2--����`�º\�������H������7�8?7�k��_�Zu�����b[�p4`�kk	   ��   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ Й��F�bϽw��VN�8�������j5>�G�Ѿ�{��{r��y��'s�Pc=�ݱ�.�c���������/�������c׮]�<v�TT��ջ,��L�@g:֍���~9�}e����,�_;�?51�����]<Ww�ߑ#G��544����r�=6w�.`�:   $ Й�W���;^ty�T�/^|Ϣ�W����G�h_T��k���Z���w�G�|{���-�(��|O��h�eΏ���m��x�t	tf���Mq��703�=�<��@Kg��X'z�l�4���e�e|l4`&:   $ �   �   	t   H@�  @   �̊�=m���câ�h�Tb��pܿ�D<v`    �̂+Wt��/[V����ml눍�;�[{;��?�  ��ccQ��T���R\4��NM]����8�kW�Ğ�Cq��  smlx(�G����T����c"ԡ�<ʨ���-x�8?��:  s�:6��8��W��>-�{ԡ�:5�vA�Y�Y���m�10<  0WƋ@)e���5��Ԓ@��:Z���:�r �9U���HΚD�	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   ���x�zN˝�b   uK�SS�㱴k�e�6�  �S����i���|��Զ�'c���I�y��P��  ̥���~��JSST����QFMݻ�x\��7�t��Cm�q��#  s�����j������hj����.
����jy,�n}�m�����ų}C  �{�[:[�:^zš��.�N�95�w�ؼ�k�p��J%������ԈC� ȧܛ�M�3+ʳ�o9001   x1�   	t   H@�  @   �   ��@  �:3��kG�x `�6���h�]�6�w���Q,��Xy�mQo��g��t4�o{ot,^�f�}w��D�X���U�ӆO�����:ypW�Ltfd߽0k���y�7����ߣQ���'�2Ї�5�z,����C=v���h�7_'Пg���{.9t   H@�3��v�^�����;���㻣�:t(������T*��g1}�s_�g��L�W]������ݵ;�����ho����Q�������Ol�F�z�����z���/�����X�jU0U�����}���1r���S$Й��M��h�5�z�Mm�Qi>�����E�~�k^���_��@?+�����'�mKcm�,����\���yOl�����;1�͉'��kmm�ŋ�Wu��_;�ۭ{�#�ԉ�S$�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:�3�j5~�#��с�������oē[�F�<5�d�C������  ��O��<S���O��D_��`~��  �J�  @���w'@���a��{fv��.�[�� ���2.���bD�`S6��8N��q�H�v%���)lCGb�@��K"�#�����$J��ؕ����j�����h�
��ٳ���|���׽Ө������   ��ņ�LMME��
Nl```�u�5�v;&'��8�f��֭�^� �!�!�3�<sn��۷�A�V�k۶mq���G�9t�P<؃'�;�-[��K_���E?�p��� ��:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@g)�kMMĞ����OZ|<�����kjj*����x�޽;zM���=�:����~222ccc�k�e�]��Y��C���;���Y�+�,�@g)^2;5O|� V�����`m�#v׮]�ڷw�ޠMNN�,�y��w��x�,�@  �:�r����}Y�b��-x���9z�/���Ϻ0z������X���{�9W_[.�����-?F�7��>ˬ��];�/�y�R	t��W�6N/X��mg�y?����6�y�ױGl��ʹAX��g�%�{��:�"�   �   	t   H@�  @   �   ��@gU4�*.9}C\�u�������g�hL̴   ��*ض~0��3⌍����K��'���  Ȥ�nGT�U#`�t�j�Y�;/;�D���Ն�w~�����'c���  ���Ӛ���Tt:����h4��nX��*:]����q~D��x�E���J� ��To5���8f^�݊N�70�1��:]�7N�0�c�ߺ.����n9 ���=;���p���WM�Dwy��U����*c�P3F&:  'Q����.�U@w	t��>c�BT�v  @��   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ ������>  ���Ntg@�	t�j�3Sq��>���l�M�  N�Fs ڳ3�7�*�^���]FWݺ����<��_{�`  ��V�o�H�~n^�����<[�aet�j��L|��3�8�#��'G���  d�Z7���Ӟ���:ګ��:]��=c�wl&��`K\�u��z{Ʀ���ާ�  2��͹�M��*v�NǍ��   ^�@  �:   $ �   �   	t   H@�  @�e�w��brdw�b���������g՟�����/6�ual����5ӇĞ;����+~"�6o�^3���1�������1���Y����m�X��v,�@gY��,ũ���@?ʡ���~/�Ź?��{2�'�?�W�cm˅���@��7Ů��T�+~�z�~��gF��� �   ��R<2�n��x��W�I���G5�T�v�۷/&''�۴iSl��{[$���b�޽�/֯_��zj��������D��O?=֭[����1::����p�v�i����xFt��xU��o�٩�GI��;���Ǚ��Ī>ic��Q=�֮C�	�ذaC�uV��jZ�����:�����*зm��7o�^3==-���r�W?���sƥ�>wu����_Ձ�3`�:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @���|z�@<��?^�g�/c"X������������h��v������q�}�E/���c�=�F#z���t0�zyܫ�徱�������S������$�Y�M��l����ʛ����m�V+��ǃ�orr2�_>˽�~����'��H   �,�e��Q���	X���T>�i�s���������E�Ͽ��^������,_��ߊ���oF��<g����g�����[����T�ei�?�O	`y���R��c�h��SU�,�4M_v�L   �   ��@  �:   $ �   �   	t   H@�  ��Dkf::�ٹ�e��  P+q>;9^n�ߛ՚�*�ގ��p@�	t  ��=;}L�?7fn+z�ht�@  (�-�ǿ�%��:�  0�N@�	tV��u�hVU<3Պv�B  ��Ϊ���7ŏ^�5���-79ێ;��[y:fZB  @��u?�����o9f��@#�:���`�p��'E:  ��:]ua	�����^|�P��K��v<   �L��UW�x󼏹����Ň���  �L��Ugn��1��yh ���  �~%���F���5�8  �^%�   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@��Z�΂7���  �*�NW����7��1ӭN�N�  ��	t��ݣq��N��o��V�t  ��	t�ꁽ�qϞ�xՙ_�������CO  @��t�'��#�3q��[b�Y�ͫ���_������L;   ��@���׿�ȁ��c���CѬ��[�}l�q�   GtVM}����  ��'�   �   	t   H@�  @   �   ��@  �:   $ �Y��#��  ������j�ޞ�<�ǉ�E�,�葉�ɱ  �^Љ�zU��Ǭ
X$��R<sd�59  ���}��u��$�Y�}G&�  X�:�v��lAo4��3�Ǭ�X$��R�ydb|�c  k]�={���vo_�.�c��Y7�#`�:K��#cO>  ��ufO��~�����E�,Z��y���z��jl������o  �N��v��W������z��3?�H����yQ}��C����^  ��w��96���~���X��R�ǡ�����v� ��T��=;s���fT��'���7�����,�@g�n���7�7�#  `�iOO���j`pA�g�����
X��R}���˨��{k��&��n}  �Zў�:��U#�z���綠��j��K �Y�N�3ZUU}�[���[✫~:  `-�f�5ϱ�����=��h=�%����<����Oe�~=���o�  �	sq>Ϯ��������7n>��,�@g9�W�{�h������p��  Y�g�K�O�������~�ؓ�Ν4��z��D�%�t:SUU}�L��>��ß����_��  �l�u^¼ݚ���͡uQ5�?s{������>�/�:�����,��+c{��_�).z�?����  �B�3�ռ��Z��y�hDc`aǞO�2���s�{�2~5`:�RrUUU_����X���@�௼'  �)!�i�涖��	�Z}�ys���׾s�8�귕������+e|+涢&�}�[�E_  }��R[�`����a�>z��������U��Ǐ<xG<����s{�²t�����]UU}��k���������Ϩ��^ @�(�@�S��|��wk��r��8�Zq���;���ɲN|_�2)(V�ϕ�����];bǧ?���  ���)q�F5��1�nQ�f�'��C�}�ȏ���~!`tVD�����7����̇c�˯�S_�# ��:838��gioG�l.�����7���p��_+��+@��bʂ�%��L��>����v\�/�G��  ���j4��<S��&Gv�=e��c�?_ց?�B:+�2�(�����?���߹!7n	 �^U�{���ټI��%���\��G���;��k1}��#�F�xK�
謨N�3SUՏ�ɻ�}���������i4�wl �ZQo��/��8�\��ث���I��+��Zӓq����C;�sdV�m�k˺�t�
謸����Dz�%��e4��~W������_�w1�~c  ��z����G]fma��f�<�E|n�xy-�ף��l)�z�����������̪_�k�:��+L��e�����*����j������ջ��w �m==  zN}l��`�;��;�w]<��Gf�߼�rY���] �隲��X��e�eT�vm��~�����q��  du�{���{?2��r��e�#]"�骲 ���;��g�jg���w����?�~��  �������}o�g�w�y����u�Ot�@��ʂ�s%ү.�����^�����0��w[\���O;;  �d������{���ѳ����N{{@�	tVEY�}�D�9e�+e�P=�o����mq�[�~\x�/.�Z�  �\황x��|$���њ�:��:��8?�
:��,؞)7��P��r���hԗ�����$�{������wŹ�{�˱ �*�uѝ_�x<������OsWP�_�E�*謺�����(��*��z�����cn�p���o�s�~sl8�  ��6�����o����gF�w���g�:뮀U&�9)��>q�%��Vn����ѧ���`���b��^g��Mq�+^�^|Q  ��t:1��C���[c�7�v��B�z����z�N��IU�7��K���ܾ�����57jC[N�m/�"6�wql<���p�1��3c`x}4� ��ǒ�NN��9���/����ȃw�m:�G��aN�����%��]���k�X��z�Z�Y�竚�� ��5;9�Vk��,�Ke�nY�# 	�N*eyg�y[	�F���2~���mg�Q��)♱g  ��S��2��}���(��d:)^`�txD	�M��2�f��qq[ʨ�o:<Xa�ׯh6�U�����v���aÆ�F��&�;���3A�6m�5�^��˝ �zyS/wbh�Z���	��><��(cGߊg������h@rkbA��_8<X%7�t�窪��X^��7�y{���7�\�/�5��o|��Hyﬕ/�*����~-�k@Y�����^{M � �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @8���������5������l6�j4�ưh������n�g�4&&&>�S��{gvvv2 ���p\ozӛF���k���e��d�"���oo��`��   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	t   H@�  @   �   ��@  �:   $ �   �   	���y����     IEND�B`�PK
     �9s[w�'<�  �  /   images/44e1934a-57d6-434e-9b76-9cc9cf9f98cc.png�PNG

   IHDR   d   �   �=��   	pHYs  �X  �X{�M   tEXtSoftware www.inkscape.org��<  qIDATx��]Y��y�o-]��>�F�iFh$�c��b6��I생�NL�<$���������)ǎ��Ā}&66X�� ��@B�f$�m$�>�ޫ���oUWwuW�t��D��4����֭��˿�V D�2$`0�	B�!C��!CȐ�!dH�2$`04�IQ���6xt���[XO���(Ļ@V"���M�ƎCtI������ĺ��sӾ,Afjߊ�o��T�N�B˲��q�*�C�Cz�4D�{\e�����̉C�<uġM3h�!��N��NÇ�y��W�n�cۥHTk����
��J�H��0d��Ma�����V,��?"�i5
�^�=3����,�Ű�Rw�T�Z.��b+�(@>9)�_V^�/�?��gsȌ�=���/�ա�_4�z��P_��������ۍ��F"����L҆���i�h��-�FZ�o ��x'P�$Cvz&���~��\OOvÒ�; ��S�.+p���@�[��-��g�о~,����G�d27 =v.?��?}��m��x��z��;>_�t�go��W����>�<N��	�􁪤NL���	J��� S��dc �����w׋��,�@R5,��eM\�YF�"-X�id���"#����qǵ��3c����0�z�h��H�����޲���}��>�� j�B8��w`�g����o�'�.�O�M��Dv�#G"��dAF3�+�wt��&0q��3g�s%�ш��K�82�)�q���͜FF��%�!�� �;e����A�w g�m����W�����u_<����z:c*8;c5$57E�ZƵ0��o@*
Y07�Bÿ�8Ά���@$�=�M ��gY��Az�%�AQ粉����R���ڣ!�p	�sn��� �W+`��.����N]��"���4Lku�Ym��n~ߛMK�C��u��a�2$`0�!$��N�Yi�5�{-��zD�t��d��t�l�A`B$WTZ{�[��R ���U�C[W���؛�� !�G`b�V݁~�KZ��R�h�x�ճ����څ���Gv��^�g�%�+���u�8��\���"0��m���0K��S�T޺f��c���O�BE��0����gN��H,a��� �-���\�f��_�S1�b�,K0>6�����-����������4Xt�!`�v<�^�4,]Z��1��v��Ld���u�p�&���AKVC��e��yX���Ca���2-`�Z�R|t���0�i�����"0M��&��x7eTl��6��]���4MLc��EDp�5�h�8܇i���3��CB,�!,�rʻ�3�IP�LԪ%\�Y-���k�	�ū�e�*�$V�|^tݺ�.��+˚5-��5��'I�f�C���/M�^�=�Qt��(Ɯ�7W�N!�j�ǝ����L�$��[Amiw�!Bf&/Z-s����,b������W���
���La��w4r��ҝdi3Q�O�fH�c9d�����Q}��灡8*�~ �t�,iҒ�½����Z%o~^N���ȕ�HR�p� |�uԘ� "C���0~ݶ�U
r�L����`U�x�h�p��(���x��R�����~��_���Z�+���[&w$����;�䇯�������͌1Ϧ�/��f�M�.ĺVp�c���*0z�2�P|��J�~�jg9S����!��G7Gh&E	֭-тĴC� �g�A�s�@���׻6nX�2���x�cId�ϸʐ��\�٢Z+�>1|��"��j*�]}�!����M+_�͐�D�O,L ��`>�a\��ộ5C��h�';K�ax/�d�B�Q��]R�V뭊}*����:����k�*g�̙��_�%+��EQ'��[���dD�I�D���f!I�2AKV���E�UŞQ�hz�O�-cc*Ix�8V��t�s/�>��-�'�#a	��fջU�m��У�ڄZ��!���a�3R7\	;#1���Vp-Y^G��wo���kK`��l�V-R�s�����	P���p��G!�2.���(0|j�r��L�ŠcS �U��t�b��V��vO��
-b��f
��AZ����#�w*����d�.�2�V���!���X���[T���5GÑB�ygIoD̔* ��n��L�ꖺR��\jGۻ`���`�b��Q�ǫ��=�|̝T�M��f�ø����_�$�an���mt�� 1�V��T��Z�l�_O��d�f�\Y\� �}^�0�Xk��w��*��Z�.���m�AY��5!�>�-]i�	�s�X�#�`F!�я2姼߶��ㄯ. �aab�f�=ˆ�d�,�,�3Ė8h$������-��ͧPU��IE�`B����]5m�f��k�l[*n�'�x7��PS!i2��(�_M�Y�k�(yҗ��c�̟L_����S�
�
�	Z�m[�"�%_�*��*�(u�5�ɜE���^��/@'�6�&���,�͹�i����l�;�&�y��i�m�Zkg)�
�4��Cv�U�Si1p3o�~,�zKu~2��O���Iѷ���M�>w
�N��iz0�i叾�юe�!񮕆�X*�$��-�����sҸeM�;��e:y��!�{j�1��M��]�@K��i�x��s^2��!2�����u��N3��ax�im]�IB�U�g ::Tfˢ���[����̈�5`�½#�f�va��]B4�6���6�EH��tJCs��u�,�g���xy+p]�e�]�/2a��C�U� ��W2�@�9-?DX����^�T��g�u<�nZ4`�g��4��{CޚC��]dZ�0�	S#��d�C�����A�\���VQ�fI*�o�!���e����~�X&C���J3�ܾ��d�旟�f�Đ}Hʤ�e��:Z�E"�Ȭ��QA$��2ʄ�Tʓ�tMG���G�);P�z^��Dd�o���a��E�C�5��`t�-��4pϐK� v�>��;�*��F��: �� [g)0I3ǥ�hSN+?�͐����X\Q�6l��;���q���+m�$������b}���k�������Է�`��Ѧ���f8r�2y�wp'�Q��r�"a�w���\����X�*�^�X��zj�ۭ\t��HȐ�#�]%�V�д����w�rz
�&���Q�#H�+|G������t��i�C�5q�u�Ϥ�+ܽ��AH�����̆���ll��*V;ٙ1��~��b_�E��A$ϳ'}<����$����"��*���b:v3*�À���nF�Q'�y]L�&�)�_�)�T�6X�%K��6��V�d���R<*4R��=�t
S��5L줃4�d�(̵x�/��߉h������?�xZ�ӳ�z�
C��-	�Ae9���Z ���j��f�?�Ԉ����i]�-K F����泐=�����vH��\�y�i����G!7~���{��{<~��($'k��ޕ�D�g������u�Cj�m���>{Ί:�9�̴��$?��^A��w�0$Wl@��d`�Cp�*��b��t��=f�Z�tB�6�����lX;�:96|
�H�Ab銒/g�����,F��si�w�$���W2D��_?ꅣ���&h�:�\�0�0]��L�V����c����Cb8x��!Qں���lYZl��1T0��(���Qʠ@�rP������vh��vٲ�Ӟ����-�Vi��K9�(We~�"1$&��c�9g��E󛺓����+�m/�S�g�a�%�u�ruD��t�)Sb5�/&V9��װ�~h�E%�`��rP���^ʟ��D�3��F�a@ F�Aǲ	_��Sn9�����4���(LN�����sC�)mզw�҅yƴu�3+��c�
i��+3��]�]C������#�f4�-�-���o�d�/�ge��e�,U��!���2d	��ֹL�뤞 M���ߌ�?}�4H�T��dR�x�����	���'�.�=�3�6@]_<���7@6����dJ��Ժl�F ���f�����d��"�6d.�Q'6�|�7C:c
־n�t���9��Ql����a���94��z�FW��-��[�Fd\b�YB3Imis�}�4+�g*��H�_z�] ���oPLi�e!{o�����]�H|����%x�M+_�8k��&`z.s�����8�za1"�W�%�[������l!�s�)[#�����9�!ʠ"w���H���];�y���d-G��v�dg�����Q1�%�Ƞ+Z�	`�M�߭��.��{���&�#t=a����i��FY����l�|jֵQ�*tUYN���̤h�L�f�hk�ۯNm�z�WfCQ���dJ!=+,�˲8H�$�8�	��$���E�9w�x�ψZ�,�N�2���=���-�Љ4���[$��_���v��N�!<� ߶۝A55
�o?��KDȑh�s��\X}'ĺʎ��0�}�����SK� %v~��|�#�J������ʠ�Z����?;=&�NlZ���o���V��Xw��u�i�udI*�B�T�(r�n�ru�t��/���d�\D˒���oCU��OA�"��fƚ�^ؼi�˖���Rp`���8��#`��*Q�D�n���`G=�nv����A%�lZ�, ��>]��Tvn�)�t�]�Q���� ��JG`��f���"�%�����d�"�*r�8贬�{�9��n�Gϙ��x��������C��x�Π�����5�ѝ
���{����ǛD�U�a�͊��Ǒ��������t�5�Ɂ��.�Ó��P�/?��s2;�|�y�����-X`��'V�H�b���J#��4��5�I��e����f���=
J�#�L+-�8$���2Xs ����xv���bf�|#�9{�
��T�tR<+=yN�q9���t���Ͳ�\��`U&��z�D@�S��*�b#���eȑ�Bl�e3��3�E�Jۖ��A���D�&_	S�a̳�30Hsz�x.���i��3�.��.$V�����N!��ͻ4(i��XHYLK�M7A��+S�uY=IOL��oVx*-�]$��� Rݞ[?ƍ���9����53���|ٺ��H��;z`��Ae���6�(�vxh�F�w|�Oe?j��bȅ�HӪg��b���H��j�J1�N�(?˱n�6�X@��-��jis�x�L'�T�i ��__|�b|���0�XZ����*ӿtUĂ�,��T���M'��R0�5@&MVb��^?������F��ϊ���u�{,�z�W�,����M�#�����!���I),���C(�T���KCo�O}gN,[rr�rP��y"��l��3T�k!S����`m�6Ȝ]�����[���O]��?�6H�X�ŔUX~�#�=�<�j�g!{�u�v�m�ݲ�v��|S�O������SfP���n�u�:Bh�6����u.�YdH��߈h�B�G_�(���9�ҙl
��^A��3��:��o�P�C�d�,o�6D��A���%}!mҽO�t��%����!r��;(��|�:ln��V��p�-��Y�>�@��w��}�`ц�ڴ?h>�JDZ�0�Q��|�:u^N��qv��A�c;�\��-,+�-a�0��L����m�F]���\���H�-�����w�t2_8�{��[��ʒ����av4��d���'V�tU��e�]^�}��4:�DkE�s�g��!:��Xi1i_ ��|Kn�F-s71%��c�Yc��缃�>e@$�e�����hl�̤Q�}$"�*�a�$ ��@��Ȓ%E�$z����}Z�����s�G2!�Dz�����[R�|�2�ڗz��D���C*�(�����A�\����[w}^0�\�jE��=w��[n���\m��vb��T�?x?�d��/gP�a5n9�fG�*�V��S�M��ٺ�vA:���6<I���#��P�S����\��m�Z���z>B�ʠ2���оvKu۵���]�� �AE�s����'��.MgP�Ƚw]�tbNNe��������H���*N������?��*|VD��o<Z<,L�c��?�὆�!CȐ�aA�����F���|,��l�y��h�!8;�3�&Q	�k��k��ڔǐs�����!i�g��"��Iτ�&�$IM�Ԅ?Ą���7`z����^���Z����:��h�z`� RI�:��G����+�9��_�?ߊ-]�}ō��v�U�G�Agh���+1r:>Yr��zdѕY1��~=��+Fa|�z��2˜CGG����r�g'����>y�W?�~�4Ő�����?�����po���7Kj$RKs���eu�G��%��N�c0�ɝ���KVr������Zұv݊%�Ov0�9pb�{�\!M��^�������5},�,&/>?������$�zon��|����[cڠ��`"�~����We����]-?s��o&������x|i̞;~�C�A���V�ز����ܰW�$�צ�Dܹ<�VF�Q7�s�
ovn�ʑi�t�ev������G�y�޲�s����_y�ɩԙY�dU���`W�C����o�H�?y"��+��K,�K\ө�WEט����~q6�7����^�i��CG�W��35��,h�I+��܋O�O-<���0�;�W�..�=��GW��g�Ϻ��30�5+�o�O�H�>�.�ڽ{w�zT*f�uk_���=��ݻWD���r�L��ܫBn}�Q�E�4�ˮ�Խ/-�����|}��]��$`0�	B�!C��!CȐ�!dH�2$`0�	B�!C��!CȐ�!dH�2$`0�	B�!C��!CȐ��J2��Y���2X�N�i$ܟ�e�U�}�bt����ʃ��_�h��֛���P��lo$ܞʼ��n ���]�P�(���v߯.;C
�D�Q
��1�X�=�'�kZ]��D���<Ӯ7�����y��8ܟ����+ey��D�_Q�ʗ0��^(��=��:���j8_�\�=~Ԏ�7M�����egH����Y��{�[L�RV�2$`0�	B�!C��!CȐ�!dH�2$`0��48�_4O    IEND�B`�PK 
     �9s[���J�O �O                  cirkitFile.jsonPK 
     �9s[                        P jsons/PK 
     �9s[ζ�g{  g{               <P jsons/user_defined.jsonPK 
     �9s[                        �� images/PK 
     �9s[������  ��  /             �� images/27b84e47-6648-4cee-a869-6ff1a6fc12fe.pngPK 
     �9s[�����  �  /             � images/50196d33-890c-4789-8115-a73c306e50dc.pngPK 
     �9s[���HT T /             � images/00941d67-c746-454a-b945-4fddefc776b2.pngPK 
     �9s[�īd}d  }d  /             c
 images/ef87c5cc-d843-475d-a868-97060fb00c54.pngPK 
     �9s[��4k� k� /             -�
 images/fd3ac6b5-800b-45c8-a4ce-2476671127d4.pngPK 
     �9s[F���9  �9  /             �- images/915d9337-ea3e-4fec-8caa-7acd53f715e1.pngPK 
     �9s[z|S�wq wq /             )h images/b949fd05-6e10-4256-9d1b-e11f1f9900de.pngPK 
     �9s[Ìs�    /             �� images/01119c27-1bad-421a-afe4-dfb48490a906.pngPK 
     �9s[�e�e�  �  /             Y� images/3d0a314b-f708-4b2c-819f-35c414b123ec.pngPK 
     �9s[�kZ��  �  /             �� images/6608fa58-7afa-4488-b64c-2b761d69d6bd.pngPK 
     �9s[�����  ��  /             � images/2c98734f-75db-43ce-800c-ea69461525e8.pngPK 
     �9s[���z"  "  /             LQ images/d4c851cf-9fb5-43cd-809f-e1699313b4d2.pngPK 
     �9s[wJ���  ��  /             �e images/f9728bc6-2422-4ead-9082-90351081a874.pngPK 
     �9s[	^�G�  �  /             � images/9ba3df0f-d630-43f7-8169-617793654d93.pngPK 
     �9s[U�p�	�  	�  /             � images/42e39361-2f02-4030-a678-a3271aadd3f6.pngPK 
     �9s[񐼛�  �  /             � images/a4af1710-95e2-4b5e-9600-8e4d90487313.pngPK 
     �9s[t���?  �?  /             � images/e2e2c934-b375-45fc-834c-534243cbf361.pngPK 
     �9s[e���  �  /             � images/6c1978d3-8c4d-4ea9-a1ba-37ab4b096c5d.pngPK 
     �9s[F���Q� Q� /             � images/028dc4b4-5e34-49e4-81aa-ecc68ea503ed.pngPK 
     �9s[���7�  �  /             �� images/06c5fde6-b2c8-47bb-9830-971f0c5559bd.pngPK 
     �9s[�;� � /             p� images/31959ea2-aec5-42cb-a646-ec7cb3b6e41e.pngPK 
     �9s[�Ƚׇ  �  /             �� images/ce527fa2-4558-4370-a5e7-21077342728a.pngPK 
     �9s["1^FHo Ho /             �  images/e2a053a3-24a6-43e1-ac97-395cbc045e87.pngPK 
     �9s[��n  n  /             p images/6b551873-9f16-48c5-b1b9-2fc6ab10f815.pngPK 
     �9s[9&��ސ ސ /             ׈ images/b01488b3-8551-4b4c-b09f-2812c4acc168.pngPK 
     �9s[d��   �   /              images/d3b73945-fe79-451b-b309-b64aab767520.pngPK 
     �9s[��Н�� �� /             �: images/0657d52a-d145-430e-bb7e-5d1be0618b5b.pngPK 
     �9s[T��T$  T$  /             �:# images/8ade0660-1c92-4b58-a3e7-adda420d3982.pngPK 
     �9s[��r�  �  /             Q_# images/022fab5a-d187-48c2-96d7-20ad2a5d1671.pngPK 
     �9s[6ah    /             Ot# images/39d025b2-988a-45cd-b457-87e73cc458ec.pngPK 
     �9s[��9PN  PN  /             �|# images/779eddd4-9cc6-4216-b155-89a4f50be07b.pngPK 
     �9s[w�'<�  �  /             M�# images/44e1934a-57d6-434e-9b76-9cc9cf9f98cc.pngPK    $ $ �  ~�#   